library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_SIGNED.ALL;

entity ConvLayer1_128 is
  generic (
  	       mult_sum      : string := "sum";
           N             : integer := 8; -- input data width
           M             : integer := 8; -- input weight width
           W             : integer := 8; -- output data width      (Note, W+SR <= N+M+4)
           SR            : integer := 2 -- data shift right before output
  	       );
  port    (
           clk     : in std_logic;
           rst     : in std_logic;
  	       d01_in, d65_in    : in std_logic_vector (9*N-1 downto 0);
           d02_in, d66_in    : in std_logic_vector (9*N-1 downto 0);
           d03_in, d67_in    : in std_logic_vector (9*N-1 downto 0);
           d04_in, d68_in    : in std_logic_vector (9*N-1 downto 0);
           d05_in, d69_in    : in std_logic_vector (9*N-1 downto 0);
           d06_in, d70_in    : in std_logic_vector (9*N-1 downto 0);
           d07_in, d71_in    : in std_logic_vector (9*N-1 downto 0);
           d08_in, d72_in    : in std_logic_vector (9*N-1 downto 0);
           d09_in, d73_in    : in std_logic_vector (9*N-1 downto 0);
           d10_in, d74_in    : in std_logic_vector (9*N-1 downto 0);
           d11_in, d75_in    : in std_logic_vector (9*N-1 downto 0);
           d12_in, d76_in    : in std_logic_vector (9*N-1 downto 0);
           d13_in, d77_in    : in std_logic_vector (9*N-1 downto 0);
           d14_in, d78_in    : in std_logic_vector (9*N-1 downto 0);
           d15_in, d79_in    : in std_logic_vector (9*N-1 downto 0);
           d16_in, d80_in    : in std_logic_vector (9*N-1 downto 0);
           d17_in, d81_in    : in std_logic_vector (9*N-1 downto 0);
           d18_in, d82_in    : in std_logic_vector (9*N-1 downto 0);
           d19_in, d83_in    : in std_logic_vector (9*N-1 downto 0);
           d20_in, d84_in    : in std_logic_vector (9*N-1 downto 0);
           d21_in, d85_in    : in std_logic_vector (9*N-1 downto 0);
           d22_in, d86_in    : in std_logic_vector (9*N-1 downto 0);
           d23_in, d87_in    : in std_logic_vector (9*N-1 downto 0);
           d24_in, d88_in    : in std_logic_vector (9*N-1 downto 0);
           d25_in, d89_in    : in std_logic_vector (9*N-1 downto 0);
           d26_in, d90_in    : in std_logic_vector (9*N-1 downto 0);
           d27_in, d91_in    : in std_logic_vector (9*N-1 downto 0);
           d28_in, d92_in    : in std_logic_vector (9*N-1 downto 0);
           d29_in, d93_in    : in std_logic_vector (9*N-1 downto 0);
           d30_in, d94_in    : in std_logic_vector (9*N-1 downto 0);
           d31_in, d95_in    : in std_logic_vector (9*N-1 downto 0);
           d32_in, d96_in    : in std_logic_vector (9*N-1 downto 0);
           d33_in, d97_in    : in std_logic_vector (9*N-1 downto 0);
           d34_in, d98_in    : in std_logic_vector (9*N-1 downto 0);
           d35_in, d99_in    : in std_logic_vector (9*N-1 downto 0);
           d36_in, d100_in   : in std_logic_vector (9*N-1 downto 0);
           d37_in, d101_in   : in std_logic_vector (9*N-1 downto 0);
           d38_in, d102_in   : in std_logic_vector (9*N-1 downto 0);
           d39_in, d103_in   : in std_logic_vector (9*N-1 downto 0);
           d40_in, d104_in   : in std_logic_vector (9*N-1 downto 0);
           d41_in, d105_in   : in std_logic_vector (9*N-1 downto 0);
           d42_in, d106_in   : in std_logic_vector (9*N-1 downto 0);
           d43_in, d107_in   : in std_logic_vector (9*N-1 downto 0);
           d44_in, d108_in   : in std_logic_vector (9*N-1 downto 0);
           d45_in, d109_in   : in std_logic_vector (9*N-1 downto 0);
           d46_in, d110_in   : in std_logic_vector (9*N-1 downto 0);
           d47_in, d111_in   : in std_logic_vector (9*N-1 downto 0);
           d48_in, d112_in   : in std_logic_vector (9*N-1 downto 0);
           d49_in, d113_in   : in std_logic_vector (9*N-1 downto 0);
           d50_in, d114_in   : in std_logic_vector (9*N-1 downto 0);
           d51_in, d115_in   : in std_logic_vector (9*N-1 downto 0);
           d52_in, d116_in   : in std_logic_vector (9*N-1 downto 0);
           d53_in, d117_in   : in std_logic_vector (9*N-1 downto 0);
           d54_in, d118_in   : in std_logic_vector (9*N-1 downto 0);
           d55_in, d119_in   : in std_logic_vector (9*N-1 downto 0);
           d56_in, d120_in   : in std_logic_vector (9*N-1 downto 0);
           d57_in, d121_in   : in std_logic_vector (9*N-1 downto 0);
           d58_in, d122_in   : in std_logic_vector (9*N-1 downto 0);
           d59_in, d123_in   : in std_logic_vector (9*N-1 downto 0);
           d60_in, d124_in   : in std_logic_vector (9*N-1 downto 0);
           d61_in, d125_in   : in std_logic_vector (9*N-1 downto 0);
           d62_in, d126_in   : in std_logic_vector (9*N-1 downto 0);
           d63_in, d127_in   : in std_logic_vector (9*N-1 downto 0);
           d64_in, d128_in   : in std_logic_vector (9*N-1 downto 0);
  	       en_in     : in std_logic;
  	       sof_in    : in std_logic; -- start of frame
  	       --sol     : in std_logic; -- start of line
  	       --eof     : in std_logic; -- end of frame

           w01_in, w65_in    : in std_logic_vector(9*M-1 downto 0);
           w02_in, w66_in    : in std_logic_vector(9*M-1 downto 0);
           w03_in, w67_in    : in std_logic_vector(9*M-1 downto 0);
           w04_in, w68_in    : in std_logic_vector(9*M-1 downto 0);
           w05_in, w69_in    : in std_logic_vector(9*M-1 downto 0);
           w06_in, w70_in    : in std_logic_vector(9*M-1 downto 0);
           w07_in, w71_in    : in std_logic_vector(9*M-1 downto 0);
           w08_in, w72_in    : in std_logic_vector(9*M-1 downto 0);
           w09_in, w73_in    : in std_logic_vector(9*M-1 downto 0);
           w10_in, w74_in    : in std_logic_vector(9*M-1 downto 0);
           w11_in, w75_in    : in std_logic_vector(9*M-1 downto 0);
           w12_in, w76_in    : in std_logic_vector(9*M-1 downto 0);
           w13_in, w77_in    : in std_logic_vector(9*M-1 downto 0);
           w14_in, w78_in    : in std_logic_vector(9*M-1 downto 0);
           w15_in, w79_in    : in std_logic_vector(9*M-1 downto 0);
           w16_in, w80_in    : in std_logic_vector(9*M-1 downto 0);
           w17_in, w81_in    : in std_logic_vector(9*M-1 downto 0);
           w18_in, w82_in    : in std_logic_vector(9*M-1 downto 0);
           w19_in, w83_in    : in std_logic_vector(9*M-1 downto 0);
           w20_in, w84_in    : in std_logic_vector(9*M-1 downto 0);
           w21_in, w85_in    : in std_logic_vector(9*M-1 downto 0);
           w22_in, w86_in    : in std_logic_vector(9*M-1 downto 0);
           w23_in, w87_in    : in std_logic_vector(9*M-1 downto 0);
           w24_in, w88_in    : in std_logic_vector(9*M-1 downto 0);
           w25_in, w89_in    : in std_logic_vector(9*M-1 downto 0);
           w26_in, w90_in    : in std_logic_vector(9*M-1 downto 0);
           w27_in, w91_in    : in std_logic_vector(9*M-1 downto 0);
           w28_in, w92_in    : in std_logic_vector(9*M-1 downto 0);
           w29_in, w93_in    : in std_logic_vector(9*M-1 downto 0);
           w30_in, w94_in    : in std_logic_vector(9*M-1 downto 0);
           w31_in, w95_in    : in std_logic_vector(9*M-1 downto 0);
           w32_in, w96_in    : in std_logic_vector(9*M-1 downto 0);
           w33_in, w97_in    : in std_logic_vector(9*M-1 downto 0);
           w34_in, w98_in    : in std_logic_vector(9*M-1 downto 0);
           w35_in, w99_in    : in std_logic_vector(9*M-1 downto 0);
           w36_in, w100_in   : in std_logic_vector(9*M-1 downto 0);
           w37_in, w101_in   : in std_logic_vector(9*M-1 downto 0);
           w38_in, w102_in   : in std_logic_vector(9*M-1 downto 0);
           w39_in, w103_in   : in std_logic_vector(9*M-1 downto 0);
           w40_in, w104_in   : in std_logic_vector(9*M-1 downto 0);
           w41_in, w105_in   : in std_logic_vector(9*M-1 downto 0);
           w42_in, w106_in   : in std_logic_vector(9*M-1 downto 0);
           w43_in, w107_in   : in std_logic_vector(9*M-1 downto 0);
           w44_in, w108_in   : in std_logic_vector(9*M-1 downto 0);
           w45_in, w109_in   : in std_logic_vector(9*M-1 downto 0);
           w46_in, w110_in   : in std_logic_vector(9*M-1 downto 0);
           w47_in, w111_in   : in std_logic_vector(9*M-1 downto 0);
           w48_in, w112_in   : in std_logic_vector(9*M-1 downto 0);
           w49_in, w113_in   : in std_logic_vector(9*M-1 downto 0);
           w50_in, w114_in   : in std_logic_vector(9*M-1 downto 0);
           w51_in, w115_in   : in std_logic_vector(9*M-1 downto 0);
           w52_in, w116_in   : in std_logic_vector(9*M-1 downto 0);
           w53_in, w117_in   : in std_logic_vector(9*M-1 downto 0);
           w54_in, w118_in   : in std_logic_vector(9*M-1 downto 0);
           w55_in, w119_in   : in std_logic_vector(9*M-1 downto 0);
           w56_in, w120_in   : in std_logic_vector(9*M-1 downto 0);
           w57_in, w121_in   : in std_logic_vector(9*M-1 downto 0);
           w58_in, w122_in   : in std_logic_vector(9*M-1 downto 0);
           w59_in, w123_in   : in std_logic_vector(9*M-1 downto 0);
           w60_in, w124_in   : in std_logic_vector(9*M-1 downto 0);
           w61_in, w125_in   : in std_logic_vector(9*M-1 downto 0);
           w62_in, w126_in   : in std_logic_vector(9*M-1 downto 0);
           w63_in, w127_in   : in std_logic_vector(9*M-1 downto 0);
           w64_in, w128_in   : in std_logic_vector(9*M-1 downto 0);

           d_out   : out std_logic_vector (W-1 downto 0);
           en_out    : out std_logic;
           sof_out   : out std_logic);
end ConvLayer1_128;

architecture a of ConvLayer1_128 is

constant EN_BIT  : integer range 0 to 1 := 0;
constant SOF_BIT : integer range 0 to 1 := 1;

component Binary_adder8 is
  generic (
           N             : integer := 8;                  -- input #1 data width, positive
           M             : integer := 8
           );
  port    (
           clk           : in  std_logic;
           rst           : in  std_logic; 

           en_in         : in  std_logic;                         
           Multiplier    : in  std_logic_vector(N-1 downto 0);    -- positive
           Multiplicand  : in  std_logic_vector(8-1 downto 0);    -- signed

           d_out         : out std_logic_vector (N + M - 1 downto 0);
           en_out        : out std_logic);                        
end component;

component ConvLayer1 is
  generic (
           mult_sum      : string := "sum";
           N             : integer := 8; -- input data width
           M             : integer := 8; -- input weight width
           W             : integer := 8; -- output data width      (Note, W+SR <= N+M+4)
           SR            : integer := 2 -- data shift right before output
           );
  port    (
           clk         : in std_logic;
           rst         : in std_logic;
           data2conv1  : in std_logic_vector (N-1 downto 0);
           data2conv2  : in std_logic_vector (N-1 downto 0);
           data2conv3  : in std_logic_vector (N-1 downto 0);
           data2conv4  : in std_logic_vector (N-1 downto 0);
           data2conv5  : in std_logic_vector (N-1 downto 0);
           data2conv6  : in std_logic_vector (N-1 downto 0);
           data2conv7  : in std_logic_vector (N-1 downto 0);
           data2conv8  : in std_logic_vector (N-1 downto 0);
           data2conv9  : in std_logic_vector (N-1 downto 0);
           en_in       : in std_logic;
           sof_in      : in std_logic; -- start of frame
           --sol     : in std_logic; -- start of line
           --eof     : in std_logic; -- end of frame

          w1           : in std_logic_vector(M-1 downto 0); -- weight matrix
          w2           : in std_logic_vector(M-1 downto 0); -- weight matrix
          w3           : in std_logic_vector(M-1 downto 0); -- weight matrix
          w4           : in std_logic_vector(M-1 downto 0); -- weight matrix
          w5           : in std_logic_vector(M-1 downto 0); -- weight matrix
          w6           : in std_logic_vector(M-1 downto 0); -- weight matrix
          w7           : in std_logic_vector(M-1 downto 0); -- weight matrix
          w8           : in std_logic_vector(M-1 downto 0); -- weight matrix
          w9           : in std_logic_vector(M-1 downto 0); -- weight matrix

           d_out       : out std_logic_vector (W-1 downto 0);
           en_out      : out std_logic;
           sof_out     : out std_logic);
end component;

signal    d01_out, d65_out    : std_logic_vector (W-1 downto 0);
signal    d02_out, d66_out    : std_logic_vector (W-1 downto 0);
signal    d03_out, d67_out    : std_logic_vector (W-1 downto 0);
signal    d04_out, d68_out    : std_logic_vector (W-1 downto 0);
signal    d05_out, d69_out    : std_logic_vector (W-1 downto 0);
signal    d06_out, d70_out    : std_logic_vector (W-1 downto 0);
signal    d07_out, d71_out    : std_logic_vector (W-1 downto 0);
signal    d08_out, d72_out    : std_logic_vector (W-1 downto 0);
signal    d09_out, d73_out    : std_logic_vector (W-1 downto 0);
signal    d10_out, d74_out    : std_logic_vector (W-1 downto 0);
signal    d11_out, d75_out    : std_logic_vector (W-1 downto 0);
signal    d12_out, d76_out    : std_logic_vector (W-1 downto 0);
signal    d13_out, d77_out    : std_logic_vector (W-1 downto 0);
signal    d14_out, d78_out    : std_logic_vector (W-1 downto 0);
signal    d15_out, d79_out    : std_logic_vector (W-1 downto 0);
signal    d16_out, d80_out    : std_logic_vector (W-1 downto 0);
signal    d17_out, d81_out    : std_logic_vector (W-1 downto 0);
signal    d18_out, d82_out    : std_logic_vector (W-1 downto 0);
signal    d19_out, d83_out    : std_logic_vector (W-1 downto 0);
signal    d20_out, d84_out    : std_logic_vector (W-1 downto 0);
signal    d21_out, d85_out    : std_logic_vector (W-1 downto 0);
signal    d22_out, d86_out    : std_logic_vector (W-1 downto 0);
signal    d23_out, d87_out    : std_logic_vector (W-1 downto 0);
signal    d24_out, d88_out    : std_logic_vector (W-1 downto 0);
signal    d25_out, d89_out    : std_logic_vector (W-1 downto 0);
signal    d26_out, d90_out    : std_logic_vector (W-1 downto 0);
signal    d27_out, d91_out    : std_logic_vector (W-1 downto 0);
signal    d28_out, d92_out    : std_logic_vector (W-1 downto 0);
signal    d29_out, d93_out    : std_logic_vector (W-1 downto 0);
signal    d30_out, d94_out    : std_logic_vector (W-1 downto 0);
signal    d31_out, d95_out    : std_logic_vector (W-1 downto 0);
signal    d32_out, d96_out    : std_logic_vector (W-1 downto 0);
signal    d33_out, d97_out    : std_logic_vector (W-1 downto 0);
signal    d34_out, d98_out    : std_logic_vector (W-1 downto 0);
signal    d35_out, d99_out    : std_logic_vector (W-1 downto 0);
signal    d36_out, d100_out   : std_logic_vector (W-1 downto 0);
signal    d37_out, d101_out   : std_logic_vector (W-1 downto 0);
signal    d38_out, d102_out   : std_logic_vector (W-1 downto 0);
signal    d39_out, d103_out   : std_logic_vector (W-1 downto 0);
signal    d40_out, d104_out   : std_logic_vector (W-1 downto 0);
signal    d41_out, d105_out   : std_logic_vector (W-1 downto 0);
signal    d42_out, d106_out   : std_logic_vector (W-1 downto 0);
signal    d43_out, d107_out   : std_logic_vector (W-1 downto 0);
signal    d44_out, d108_out   : std_logic_vector (W-1 downto 0);
signal    d45_out, d109_out   : std_logic_vector (W-1 downto 0);
signal    d46_out, d110_out   : std_logic_vector (W-1 downto 0);
signal    d47_out, d111_out   : std_logic_vector (W-1 downto 0);
signal    d48_out, d112_out   : std_logic_vector (W-1 downto 0);
signal    d49_out, d113_out   : std_logic_vector (W-1 downto 0);
signal    d50_out, d114_out   : std_logic_vector (W-1 downto 0);
signal    d51_out, d115_out   : std_logic_vector (W-1 downto 0);
signal    d52_out, d116_out   : std_logic_vector (W-1 downto 0);
signal    d53_out, d117_out   : std_logic_vector (W-1 downto 0);
signal    d54_out, d118_out   : std_logic_vector (W-1 downto 0);
signal    d55_out, d119_out   : std_logic_vector (W-1 downto 0);
signal    d56_out, d120_out   : std_logic_vector (W-1 downto 0);
signal    d57_out, d121_out   : std_logic_vector (W-1 downto 0);
signal    d58_out, d122_out   : std_logic_vector (W-1 downto 0);
signal    d59_out, d123_out   : std_logic_vector (W-1 downto 0);
signal    d60_out, d124_out   : std_logic_vector (W-1 downto 0);
signal    d61_out, d125_out   : std_logic_vector (W-1 downto 0);
signal    d62_out, d126_out   : std_logic_vector (W-1 downto 0);
signal    d63_out, d127_out   : std_logic_vector (W-1 downto 0);
signal    d64_out, d128_out   : std_logic_vector (W-1 downto 0);

signal    sum1 , sum22     : std_logic_vector (W+1 downto 0); 
signal    sum2 , sum23     : std_logic_vector (W+1 downto 0); 
signal    sum3 , sum24     : std_logic_vector (W+1 downto 0); 
signal    sum4 , sum25     : std_logic_vector (W+1 downto 0); 
signal    sum5 , sum26     : std_logic_vector (W+1 downto 0); 
signal    sum6 , sum27     : std_logic_vector (W+1 downto 0); 
signal    sum7 , sum28     : std_logic_vector (W+1 downto 0); 
signal    sum8 , sum29     : std_logic_vector (W+1 downto 0); 
signal    sum9 , sum30     : std_logic_vector (W+1 downto 0); 
signal    sum10, sum31     : std_logic_vector (W+1 downto 0); 
signal    sum11, sum32     : std_logic_vector (W+1 downto 0); 
signal    sum12, sum33     : std_logic_vector (W+1 downto 0); 
signal    sum13, sum34     : std_logic_vector (W+1 downto 0); 
signal    sum14, sum35     : std_logic_vector (W+1 downto 0); 
signal    sum15, sum36     : std_logic_vector (W+1 downto 0); 
signal    sum16, sum37     : std_logic_vector (W+1 downto 0); 
       
signal    sum17, sum38     : std_logic_vector (W+3 downto 0);   
signal    sum18, sum39     : std_logic_vector (W+3 downto 0);   
signal    sum19, sum40     : std_logic_vector (W+3 downto 0); 
signal    sum20, sum41     : std_logic_vector (W+3 downto 0); 
       
signal    sum21, sum42     : std_logic_vector (W+5 downto 0); 

signal    sum43            : std_logic_vector (W+6 downto 0); 

begin


CL01: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d01_in(9*N-1 downto 8*N),data2conv2 =>d01_in(8*N-1 downto 7*N),data2conv3 =>d01_in(7*N-1 downto 6*N),data2conv4 =>d01_in(6*N-1 downto 5*N),data2conv5 =>d01_in(5*N-1 downto 4*N),data2conv6 =>d01_in(4*N-1 downto 3*N),data2conv7 =>d01_in(3*N-1 downto 2*N),data2conv8 =>d01_in(2*N-1 downto N),data2conv9 =>d01_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d01_in(9*N-1 downto 8*N),w2 => d01_in(8*N-1 downto 7*N),w3 => d01_in(7*N-1 downto 6*N),w4 => d01_in(6*N-1 downto 5*N),w5 => d01_in(5*N-1 downto 4*N),w6 => d01_in(4*N-1 downto 3*N),w7 => d01_in(3*N-1 downto 2*N),w8 => d01_in(2*N-1 downto N),w9 => d01_in(N-1 downto 0 ),d_out => d01_out,en_out =>en_out,sof_out=>sof_out);
CL02: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d02_in(9*N-1 downto 8*N),data2conv2 =>d02_in(8*N-1 downto 7*N),data2conv3 =>d02_in(7*N-1 downto 6*N),data2conv4 =>d02_in(6*N-1 downto 5*N),data2conv5 =>d02_in(5*N-1 downto 4*N),data2conv6 =>d02_in(4*N-1 downto 3*N),data2conv7 =>d02_in(3*N-1 downto 2*N),data2conv8 =>d02_in(2*N-1 downto N),data2conv9 =>d02_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d02_in(9*N-1 downto 8*N),w2 => d02_in(8*N-1 downto 7*N),w3 => d02_in(7*N-1 downto 6*N),w4 => d02_in(6*N-1 downto 5*N),w5 => d02_in(5*N-1 downto 4*N),w6 => d02_in(4*N-1 downto 3*N),w7 => d02_in(3*N-1 downto 2*N),w8 => d02_in(2*N-1 downto N),w9 => d02_in(N-1 downto 0 ),d_out => d02_out,en_out =>open  ,sof_out=>open   );
CL03: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d03_in(9*N-1 downto 8*N),data2conv2 =>d03_in(8*N-1 downto 7*N),data2conv3 =>d03_in(7*N-1 downto 6*N),data2conv4 =>d03_in(6*N-1 downto 5*N),data2conv5 =>d03_in(5*N-1 downto 4*N),data2conv6 =>d03_in(4*N-1 downto 3*N),data2conv7 =>d03_in(3*N-1 downto 2*N),data2conv8 =>d03_in(2*N-1 downto N),data2conv9 =>d03_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d03_in(9*N-1 downto 8*N),w2 => d03_in(8*N-1 downto 7*N),w3 => d03_in(7*N-1 downto 6*N),w4 => d03_in(6*N-1 downto 5*N),w5 => d03_in(5*N-1 downto 4*N),w6 => d03_in(4*N-1 downto 3*N),w7 => d03_in(3*N-1 downto 2*N),w8 => d03_in(2*N-1 downto N),w9 => d03_in(N-1 downto 0 ),d_out => d03_out,en_out =>open  ,sof_out=>open   );
CL04: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d04_in(9*N-1 downto 8*N),data2conv2 =>d04_in(8*N-1 downto 7*N),data2conv3 =>d04_in(7*N-1 downto 6*N),data2conv4 =>d04_in(6*N-1 downto 5*N),data2conv5 =>d04_in(5*N-1 downto 4*N),data2conv6 =>d04_in(4*N-1 downto 3*N),data2conv7 =>d04_in(3*N-1 downto 2*N),data2conv8 =>d04_in(2*N-1 downto N),data2conv9 =>d04_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d04_in(9*N-1 downto 8*N),w2 => d04_in(8*N-1 downto 7*N),w3 => d04_in(7*N-1 downto 6*N),w4 => d04_in(6*N-1 downto 5*N),w5 => d04_in(5*N-1 downto 4*N),w6 => d04_in(4*N-1 downto 3*N),w7 => d04_in(3*N-1 downto 2*N),w8 => d04_in(2*N-1 downto N),w9 => d04_in(N-1 downto 0 ),d_out => d04_out,en_out =>open  ,sof_out=>open   );
CL05: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d05_in(9*N-1 downto 8*N),data2conv2 =>d05_in(8*N-1 downto 7*N),data2conv3 =>d05_in(7*N-1 downto 6*N),data2conv4 =>d05_in(6*N-1 downto 5*N),data2conv5 =>d05_in(5*N-1 downto 4*N),data2conv6 =>d05_in(4*N-1 downto 3*N),data2conv7 =>d05_in(3*N-1 downto 2*N),data2conv8 =>d05_in(2*N-1 downto N),data2conv9 =>d05_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d05_in(9*N-1 downto 8*N),w2 => d05_in(8*N-1 downto 7*N),w3 => d05_in(7*N-1 downto 6*N),w4 => d05_in(6*N-1 downto 5*N),w5 => d05_in(5*N-1 downto 4*N),w6 => d05_in(4*N-1 downto 3*N),w7 => d05_in(3*N-1 downto 2*N),w8 => d05_in(2*N-1 downto N),w9 => d05_in(N-1 downto 0 ),d_out => d05_out,en_out =>open  ,sof_out=>open   );
CL06: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d06_in(9*N-1 downto 8*N),data2conv2 =>d06_in(8*N-1 downto 7*N),data2conv3 =>d06_in(7*N-1 downto 6*N),data2conv4 =>d06_in(6*N-1 downto 5*N),data2conv5 =>d06_in(5*N-1 downto 4*N),data2conv6 =>d06_in(4*N-1 downto 3*N),data2conv7 =>d06_in(3*N-1 downto 2*N),data2conv8 =>d06_in(2*N-1 downto N),data2conv9 =>d06_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d06_in(9*N-1 downto 8*N),w2 => d06_in(8*N-1 downto 7*N),w3 => d06_in(7*N-1 downto 6*N),w4 => d06_in(6*N-1 downto 5*N),w5 => d06_in(5*N-1 downto 4*N),w6 => d06_in(4*N-1 downto 3*N),w7 => d06_in(3*N-1 downto 2*N),w8 => d06_in(2*N-1 downto N),w9 => d06_in(N-1 downto 0 ),d_out => d06_out,en_out =>open  ,sof_out=>open   );
CL07: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d07_in(9*N-1 downto 8*N),data2conv2 =>d07_in(8*N-1 downto 7*N),data2conv3 =>d07_in(7*N-1 downto 6*N),data2conv4 =>d07_in(6*N-1 downto 5*N),data2conv5 =>d07_in(5*N-1 downto 4*N),data2conv6 =>d07_in(4*N-1 downto 3*N),data2conv7 =>d07_in(3*N-1 downto 2*N),data2conv8 =>d07_in(2*N-1 downto N),data2conv9 =>d07_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d07_in(9*N-1 downto 8*N),w2 => d07_in(8*N-1 downto 7*N),w3 => d07_in(7*N-1 downto 6*N),w4 => d07_in(6*N-1 downto 5*N),w5 => d07_in(5*N-1 downto 4*N),w6 => d07_in(4*N-1 downto 3*N),w7 => d07_in(3*N-1 downto 2*N),w8 => d07_in(2*N-1 downto N),w9 => d07_in(N-1 downto 0 ),d_out => d07_out,en_out =>open  ,sof_out=>open   );
CL08: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d08_in(9*N-1 downto 8*N),data2conv2 =>d08_in(8*N-1 downto 7*N),data2conv3 =>d08_in(7*N-1 downto 6*N),data2conv4 =>d08_in(6*N-1 downto 5*N),data2conv5 =>d08_in(5*N-1 downto 4*N),data2conv6 =>d08_in(4*N-1 downto 3*N),data2conv7 =>d08_in(3*N-1 downto 2*N),data2conv8 =>d08_in(2*N-1 downto N),data2conv9 =>d08_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d08_in(9*N-1 downto 8*N),w2 => d08_in(8*N-1 downto 7*N),w3 => d08_in(7*N-1 downto 6*N),w4 => d08_in(6*N-1 downto 5*N),w5 => d08_in(5*N-1 downto 4*N),w6 => d08_in(4*N-1 downto 3*N),w7 => d08_in(3*N-1 downto 2*N),w8 => d08_in(2*N-1 downto N),w9 => d08_in(N-1 downto 0 ),d_out => d08_out,en_out =>open  ,sof_out=>open   );
CL09: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d09_in(9*N-1 downto 8*N),data2conv2 =>d09_in(8*N-1 downto 7*N),data2conv3 =>d09_in(7*N-1 downto 6*N),data2conv4 =>d09_in(6*N-1 downto 5*N),data2conv5 =>d09_in(5*N-1 downto 4*N),data2conv6 =>d09_in(4*N-1 downto 3*N),data2conv7 =>d09_in(3*N-1 downto 2*N),data2conv8 =>d09_in(2*N-1 downto N),data2conv9 =>d09_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d09_in(9*N-1 downto 8*N),w2 => d09_in(8*N-1 downto 7*N),w3 => d09_in(7*N-1 downto 6*N),w4 => d09_in(6*N-1 downto 5*N),w5 => d09_in(5*N-1 downto 4*N),w6 => d09_in(4*N-1 downto 3*N),w7 => d09_in(3*N-1 downto 2*N),w8 => d09_in(2*N-1 downto N),w9 => d09_in(N-1 downto 0 ),d_out => d09_out,en_out =>open  ,sof_out=>open   );
CL10: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d10_in(9*N-1 downto 8*N),data2conv2 =>d10_in(8*N-1 downto 7*N),data2conv3 =>d10_in(7*N-1 downto 6*N),data2conv4 =>d10_in(6*N-1 downto 5*N),data2conv5 =>d10_in(5*N-1 downto 4*N),data2conv6 =>d10_in(4*N-1 downto 3*N),data2conv7 =>d10_in(3*N-1 downto 2*N),data2conv8 =>d10_in(2*N-1 downto N),data2conv9 =>d10_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d10_in(9*N-1 downto 8*N),w2 => d10_in(8*N-1 downto 7*N),w3 => d10_in(7*N-1 downto 6*N),w4 => d10_in(6*N-1 downto 5*N),w5 => d10_in(5*N-1 downto 4*N),w6 => d10_in(4*N-1 downto 3*N),w7 => d10_in(3*N-1 downto 2*N),w8 => d10_in(2*N-1 downto N),w9 => d10_in(N-1 downto 0 ),d_out => d10_out,en_out =>open  ,sof_out=>open   );
CL11: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d11_in(9*N-1 downto 8*N),data2conv2 =>d11_in(8*N-1 downto 7*N),data2conv3 =>d11_in(7*N-1 downto 6*N),data2conv4 =>d11_in(6*N-1 downto 5*N),data2conv5 =>d11_in(5*N-1 downto 4*N),data2conv6 =>d11_in(4*N-1 downto 3*N),data2conv7 =>d11_in(3*N-1 downto 2*N),data2conv8 =>d11_in(2*N-1 downto N),data2conv9 =>d11_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d11_in(9*N-1 downto 8*N),w2 => d11_in(8*N-1 downto 7*N),w3 => d11_in(7*N-1 downto 6*N),w4 => d11_in(6*N-1 downto 5*N),w5 => d11_in(5*N-1 downto 4*N),w6 => d11_in(4*N-1 downto 3*N),w7 => d11_in(3*N-1 downto 2*N),w8 => d11_in(2*N-1 downto N),w9 => d11_in(N-1 downto 0 ),d_out => d11_out,en_out =>open  ,sof_out=>open   );
CL12: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d12_in(9*N-1 downto 8*N),data2conv2 =>d12_in(8*N-1 downto 7*N),data2conv3 =>d12_in(7*N-1 downto 6*N),data2conv4 =>d12_in(6*N-1 downto 5*N),data2conv5 =>d12_in(5*N-1 downto 4*N),data2conv6 =>d12_in(4*N-1 downto 3*N),data2conv7 =>d12_in(3*N-1 downto 2*N),data2conv8 =>d12_in(2*N-1 downto N),data2conv9 =>d12_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d12_in(9*N-1 downto 8*N),w2 => d12_in(8*N-1 downto 7*N),w3 => d12_in(7*N-1 downto 6*N),w4 => d12_in(6*N-1 downto 5*N),w5 => d12_in(5*N-1 downto 4*N),w6 => d12_in(4*N-1 downto 3*N),w7 => d12_in(3*N-1 downto 2*N),w8 => d12_in(2*N-1 downto N),w9 => d12_in(N-1 downto 0 ),d_out => d12_out,en_out =>open  ,sof_out=>open   );
CL13: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d13_in(9*N-1 downto 8*N),data2conv2 =>d13_in(8*N-1 downto 7*N),data2conv3 =>d13_in(7*N-1 downto 6*N),data2conv4 =>d13_in(6*N-1 downto 5*N),data2conv5 =>d13_in(5*N-1 downto 4*N),data2conv6 =>d13_in(4*N-1 downto 3*N),data2conv7 =>d13_in(3*N-1 downto 2*N),data2conv8 =>d13_in(2*N-1 downto N),data2conv9 =>d13_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d13_in(9*N-1 downto 8*N),w2 => d13_in(8*N-1 downto 7*N),w3 => d13_in(7*N-1 downto 6*N),w4 => d13_in(6*N-1 downto 5*N),w5 => d13_in(5*N-1 downto 4*N),w6 => d13_in(4*N-1 downto 3*N),w7 => d13_in(3*N-1 downto 2*N),w8 => d13_in(2*N-1 downto N),w9 => d13_in(N-1 downto 0 ),d_out => d13_out,en_out =>open  ,sof_out=>open   );
CL14: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d14_in(9*N-1 downto 8*N),data2conv2 =>d14_in(8*N-1 downto 7*N),data2conv3 =>d14_in(7*N-1 downto 6*N),data2conv4 =>d14_in(6*N-1 downto 5*N),data2conv5 =>d14_in(5*N-1 downto 4*N),data2conv6 =>d14_in(4*N-1 downto 3*N),data2conv7 =>d14_in(3*N-1 downto 2*N),data2conv8 =>d14_in(2*N-1 downto N),data2conv9 =>d14_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d14_in(9*N-1 downto 8*N),w2 => d14_in(8*N-1 downto 7*N),w3 => d14_in(7*N-1 downto 6*N),w4 => d14_in(6*N-1 downto 5*N),w5 => d14_in(5*N-1 downto 4*N),w6 => d14_in(4*N-1 downto 3*N),w7 => d14_in(3*N-1 downto 2*N),w8 => d14_in(2*N-1 downto N),w9 => d14_in(N-1 downto 0 ),d_out => d14_out,en_out =>open  ,sof_out=>open   );
CL15: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d15_in(9*N-1 downto 8*N),data2conv2 =>d15_in(8*N-1 downto 7*N),data2conv3 =>d15_in(7*N-1 downto 6*N),data2conv4 =>d15_in(6*N-1 downto 5*N),data2conv5 =>d15_in(5*N-1 downto 4*N),data2conv6 =>d15_in(4*N-1 downto 3*N),data2conv7 =>d15_in(3*N-1 downto 2*N),data2conv8 =>d15_in(2*N-1 downto N),data2conv9 =>d15_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d15_in(9*N-1 downto 8*N),w2 => d15_in(8*N-1 downto 7*N),w3 => d15_in(7*N-1 downto 6*N),w4 => d15_in(6*N-1 downto 5*N),w5 => d15_in(5*N-1 downto 4*N),w6 => d15_in(4*N-1 downto 3*N),w7 => d15_in(3*N-1 downto 2*N),w8 => d15_in(2*N-1 downto N),w9 => d15_in(N-1 downto 0 ),d_out => d15_out,en_out =>open  ,sof_out=>open   );
CL16: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d16_in(9*N-1 downto 8*N),data2conv2 =>d16_in(8*N-1 downto 7*N),data2conv3 =>d16_in(7*N-1 downto 6*N),data2conv4 =>d16_in(6*N-1 downto 5*N),data2conv5 =>d16_in(5*N-1 downto 4*N),data2conv6 =>d16_in(4*N-1 downto 3*N),data2conv7 =>d16_in(3*N-1 downto 2*N),data2conv8 =>d16_in(2*N-1 downto N),data2conv9 =>d16_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d16_in(9*N-1 downto 8*N),w2 => d16_in(8*N-1 downto 7*N),w3 => d16_in(7*N-1 downto 6*N),w4 => d16_in(6*N-1 downto 5*N),w5 => d16_in(5*N-1 downto 4*N),w6 => d16_in(4*N-1 downto 3*N),w7 => d16_in(3*N-1 downto 2*N),w8 => d16_in(2*N-1 downto N),w9 => d16_in(N-1 downto 0 ),d_out => d16_out,en_out =>open  ,sof_out=>open   );
CL17: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d17_in(9*N-1 downto 8*N),data2conv2 =>d17_in(8*N-1 downto 7*N),data2conv3 =>d17_in(7*N-1 downto 6*N),data2conv4 =>d17_in(6*N-1 downto 5*N),data2conv5 =>d17_in(5*N-1 downto 4*N),data2conv6 =>d17_in(4*N-1 downto 3*N),data2conv7 =>d17_in(3*N-1 downto 2*N),data2conv8 =>d17_in(2*N-1 downto N),data2conv9 =>d17_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d17_in(9*N-1 downto 8*N),w2 => d17_in(8*N-1 downto 7*N),w3 => d17_in(7*N-1 downto 6*N),w4 => d17_in(6*N-1 downto 5*N),w5 => d17_in(5*N-1 downto 4*N),w6 => d17_in(4*N-1 downto 3*N),w7 => d17_in(3*N-1 downto 2*N),w8 => d17_in(2*N-1 downto N),w9 => d17_in(N-1 downto 0 ),d_out => d17_out,en_out =>open  ,sof_out=>open   );
CL18: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d18_in(9*N-1 downto 8*N),data2conv2 =>d18_in(8*N-1 downto 7*N),data2conv3 =>d18_in(7*N-1 downto 6*N),data2conv4 =>d18_in(6*N-1 downto 5*N),data2conv5 =>d18_in(5*N-1 downto 4*N),data2conv6 =>d18_in(4*N-1 downto 3*N),data2conv7 =>d18_in(3*N-1 downto 2*N),data2conv8 =>d18_in(2*N-1 downto N),data2conv9 =>d18_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d18_in(9*N-1 downto 8*N),w2 => d18_in(8*N-1 downto 7*N),w3 => d18_in(7*N-1 downto 6*N),w4 => d18_in(6*N-1 downto 5*N),w5 => d18_in(5*N-1 downto 4*N),w6 => d18_in(4*N-1 downto 3*N),w7 => d18_in(3*N-1 downto 2*N),w8 => d18_in(2*N-1 downto N),w9 => d18_in(N-1 downto 0 ),d_out => d18_out,en_out =>open  ,sof_out=>open   );
CL19: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d19_in(9*N-1 downto 8*N),data2conv2 =>d19_in(8*N-1 downto 7*N),data2conv3 =>d19_in(7*N-1 downto 6*N),data2conv4 =>d19_in(6*N-1 downto 5*N),data2conv5 =>d19_in(5*N-1 downto 4*N),data2conv6 =>d19_in(4*N-1 downto 3*N),data2conv7 =>d19_in(3*N-1 downto 2*N),data2conv8 =>d19_in(2*N-1 downto N),data2conv9 =>d19_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d19_in(9*N-1 downto 8*N),w2 => d19_in(8*N-1 downto 7*N),w3 => d19_in(7*N-1 downto 6*N),w4 => d19_in(6*N-1 downto 5*N),w5 => d19_in(5*N-1 downto 4*N),w6 => d19_in(4*N-1 downto 3*N),w7 => d19_in(3*N-1 downto 2*N),w8 => d19_in(2*N-1 downto N),w9 => d19_in(N-1 downto 0 ),d_out => d19_out,en_out =>open  ,sof_out=>open   );
CL20: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d20_in(9*N-1 downto 8*N),data2conv2 =>d20_in(8*N-1 downto 7*N),data2conv3 =>d20_in(7*N-1 downto 6*N),data2conv4 =>d20_in(6*N-1 downto 5*N),data2conv5 =>d20_in(5*N-1 downto 4*N),data2conv6 =>d20_in(4*N-1 downto 3*N),data2conv7 =>d20_in(3*N-1 downto 2*N),data2conv8 =>d20_in(2*N-1 downto N),data2conv9 =>d20_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d20_in(9*N-1 downto 8*N),w2 => d20_in(8*N-1 downto 7*N),w3 => d20_in(7*N-1 downto 6*N),w4 => d20_in(6*N-1 downto 5*N),w5 => d20_in(5*N-1 downto 4*N),w6 => d20_in(4*N-1 downto 3*N),w7 => d20_in(3*N-1 downto 2*N),w8 => d20_in(2*N-1 downto N),w9 => d20_in(N-1 downto 0 ),d_out => d20_out,en_out =>open  ,sof_out=>open   );
CL21: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d21_in(9*N-1 downto 8*N),data2conv2 =>d21_in(8*N-1 downto 7*N),data2conv3 =>d21_in(7*N-1 downto 6*N),data2conv4 =>d21_in(6*N-1 downto 5*N),data2conv5 =>d21_in(5*N-1 downto 4*N),data2conv6 =>d21_in(4*N-1 downto 3*N),data2conv7 =>d21_in(3*N-1 downto 2*N),data2conv8 =>d21_in(2*N-1 downto N),data2conv9 =>d21_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d21_in(9*N-1 downto 8*N),w2 => d21_in(8*N-1 downto 7*N),w3 => d21_in(7*N-1 downto 6*N),w4 => d21_in(6*N-1 downto 5*N),w5 => d21_in(5*N-1 downto 4*N),w6 => d21_in(4*N-1 downto 3*N),w7 => d21_in(3*N-1 downto 2*N),w8 => d21_in(2*N-1 downto N),w9 => d21_in(N-1 downto 0 ),d_out => d21_out,en_out =>open  ,sof_out=>open   );
CL22: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d22_in(9*N-1 downto 8*N),data2conv2 =>d22_in(8*N-1 downto 7*N),data2conv3 =>d22_in(7*N-1 downto 6*N),data2conv4 =>d22_in(6*N-1 downto 5*N),data2conv5 =>d22_in(5*N-1 downto 4*N),data2conv6 =>d22_in(4*N-1 downto 3*N),data2conv7 =>d22_in(3*N-1 downto 2*N),data2conv8 =>d22_in(2*N-1 downto N),data2conv9 =>d22_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d22_in(9*N-1 downto 8*N),w2 => d22_in(8*N-1 downto 7*N),w3 => d22_in(7*N-1 downto 6*N),w4 => d22_in(6*N-1 downto 5*N),w5 => d22_in(5*N-1 downto 4*N),w6 => d22_in(4*N-1 downto 3*N),w7 => d22_in(3*N-1 downto 2*N),w8 => d22_in(2*N-1 downto N),w9 => d22_in(N-1 downto 0 ),d_out => d22_out,en_out =>open  ,sof_out=>open   );
CL23: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d23_in(9*N-1 downto 8*N),data2conv2 =>d23_in(8*N-1 downto 7*N),data2conv3 =>d23_in(7*N-1 downto 6*N),data2conv4 =>d23_in(6*N-1 downto 5*N),data2conv5 =>d23_in(5*N-1 downto 4*N),data2conv6 =>d23_in(4*N-1 downto 3*N),data2conv7 =>d23_in(3*N-1 downto 2*N),data2conv8 =>d23_in(2*N-1 downto N),data2conv9 =>d23_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d23_in(9*N-1 downto 8*N),w2 => d23_in(8*N-1 downto 7*N),w3 => d23_in(7*N-1 downto 6*N),w4 => d23_in(6*N-1 downto 5*N),w5 => d23_in(5*N-1 downto 4*N),w6 => d23_in(4*N-1 downto 3*N),w7 => d23_in(3*N-1 downto 2*N),w8 => d23_in(2*N-1 downto N),w9 => d23_in(N-1 downto 0 ),d_out => d23_out,en_out =>open  ,sof_out=>open   );
CL24: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d24_in(9*N-1 downto 8*N),data2conv2 =>d24_in(8*N-1 downto 7*N),data2conv3 =>d24_in(7*N-1 downto 6*N),data2conv4 =>d24_in(6*N-1 downto 5*N),data2conv5 =>d24_in(5*N-1 downto 4*N),data2conv6 =>d24_in(4*N-1 downto 3*N),data2conv7 =>d24_in(3*N-1 downto 2*N),data2conv8 =>d24_in(2*N-1 downto N),data2conv9 =>d24_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d24_in(9*N-1 downto 8*N),w2 => d24_in(8*N-1 downto 7*N),w3 => d24_in(7*N-1 downto 6*N),w4 => d24_in(6*N-1 downto 5*N),w5 => d24_in(5*N-1 downto 4*N),w6 => d24_in(4*N-1 downto 3*N),w7 => d24_in(3*N-1 downto 2*N),w8 => d24_in(2*N-1 downto N),w9 => d24_in(N-1 downto 0 ),d_out => d24_out,en_out =>open  ,sof_out=>open   );
CL25: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d25_in(9*N-1 downto 8*N),data2conv2 =>d25_in(8*N-1 downto 7*N),data2conv3 =>d25_in(7*N-1 downto 6*N),data2conv4 =>d25_in(6*N-1 downto 5*N),data2conv5 =>d25_in(5*N-1 downto 4*N),data2conv6 =>d25_in(4*N-1 downto 3*N),data2conv7 =>d25_in(3*N-1 downto 2*N),data2conv8 =>d25_in(2*N-1 downto N),data2conv9 =>d25_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d25_in(9*N-1 downto 8*N),w2 => d25_in(8*N-1 downto 7*N),w3 => d25_in(7*N-1 downto 6*N),w4 => d25_in(6*N-1 downto 5*N),w5 => d25_in(5*N-1 downto 4*N),w6 => d25_in(4*N-1 downto 3*N),w7 => d25_in(3*N-1 downto 2*N),w8 => d25_in(2*N-1 downto N),w9 => d25_in(N-1 downto 0 ),d_out => d25_out,en_out =>open  ,sof_out=>open   );
CL26: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d26_in(9*N-1 downto 8*N),data2conv2 =>d26_in(8*N-1 downto 7*N),data2conv3 =>d26_in(7*N-1 downto 6*N),data2conv4 =>d26_in(6*N-1 downto 5*N),data2conv5 =>d26_in(5*N-1 downto 4*N),data2conv6 =>d26_in(4*N-1 downto 3*N),data2conv7 =>d26_in(3*N-1 downto 2*N),data2conv8 =>d26_in(2*N-1 downto N),data2conv9 =>d26_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d26_in(9*N-1 downto 8*N),w2 => d26_in(8*N-1 downto 7*N),w3 => d26_in(7*N-1 downto 6*N),w4 => d26_in(6*N-1 downto 5*N),w5 => d26_in(5*N-1 downto 4*N),w6 => d26_in(4*N-1 downto 3*N),w7 => d26_in(3*N-1 downto 2*N),w8 => d26_in(2*N-1 downto N),w9 => d26_in(N-1 downto 0 ),d_out => d26_out,en_out =>open  ,sof_out=>open   );
CL27: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d27_in(9*N-1 downto 8*N),data2conv2 =>d27_in(8*N-1 downto 7*N),data2conv3 =>d27_in(7*N-1 downto 6*N),data2conv4 =>d27_in(6*N-1 downto 5*N),data2conv5 =>d27_in(5*N-1 downto 4*N),data2conv6 =>d27_in(4*N-1 downto 3*N),data2conv7 =>d27_in(3*N-1 downto 2*N),data2conv8 =>d27_in(2*N-1 downto N),data2conv9 =>d27_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d27_in(9*N-1 downto 8*N),w2 => d27_in(8*N-1 downto 7*N),w3 => d27_in(7*N-1 downto 6*N),w4 => d27_in(6*N-1 downto 5*N),w5 => d27_in(5*N-1 downto 4*N),w6 => d27_in(4*N-1 downto 3*N),w7 => d27_in(3*N-1 downto 2*N),w8 => d27_in(2*N-1 downto N),w9 => d27_in(N-1 downto 0 ),d_out => d27_out,en_out =>open  ,sof_out=>open   );
CL28: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d28_in(9*N-1 downto 8*N),data2conv2 =>d28_in(8*N-1 downto 7*N),data2conv3 =>d28_in(7*N-1 downto 6*N),data2conv4 =>d28_in(6*N-1 downto 5*N),data2conv5 =>d28_in(5*N-1 downto 4*N),data2conv6 =>d28_in(4*N-1 downto 3*N),data2conv7 =>d28_in(3*N-1 downto 2*N),data2conv8 =>d28_in(2*N-1 downto N),data2conv9 =>d28_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d28_in(9*N-1 downto 8*N),w2 => d28_in(8*N-1 downto 7*N),w3 => d28_in(7*N-1 downto 6*N),w4 => d28_in(6*N-1 downto 5*N),w5 => d28_in(5*N-1 downto 4*N),w6 => d28_in(4*N-1 downto 3*N),w7 => d28_in(3*N-1 downto 2*N),w8 => d28_in(2*N-1 downto N),w9 => d28_in(N-1 downto 0 ),d_out => d28_out,en_out =>open  ,sof_out=>open   );
CL29: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d29_in(9*N-1 downto 8*N),data2conv2 =>d29_in(8*N-1 downto 7*N),data2conv3 =>d29_in(7*N-1 downto 6*N),data2conv4 =>d29_in(6*N-1 downto 5*N),data2conv5 =>d29_in(5*N-1 downto 4*N),data2conv6 =>d29_in(4*N-1 downto 3*N),data2conv7 =>d29_in(3*N-1 downto 2*N),data2conv8 =>d29_in(2*N-1 downto N),data2conv9 =>d29_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d29_in(9*N-1 downto 8*N),w2 => d29_in(8*N-1 downto 7*N),w3 => d29_in(7*N-1 downto 6*N),w4 => d29_in(6*N-1 downto 5*N),w5 => d29_in(5*N-1 downto 4*N),w6 => d29_in(4*N-1 downto 3*N),w7 => d29_in(3*N-1 downto 2*N),w8 => d29_in(2*N-1 downto N),w9 => d29_in(N-1 downto 0 ),d_out => d29_out,en_out =>open  ,sof_out=>open   );
CL30: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d30_in(9*N-1 downto 8*N),data2conv2 =>d30_in(8*N-1 downto 7*N),data2conv3 =>d30_in(7*N-1 downto 6*N),data2conv4 =>d30_in(6*N-1 downto 5*N),data2conv5 =>d30_in(5*N-1 downto 4*N),data2conv6 =>d30_in(4*N-1 downto 3*N),data2conv7 =>d30_in(3*N-1 downto 2*N),data2conv8 =>d30_in(2*N-1 downto N),data2conv9 =>d30_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d30_in(9*N-1 downto 8*N),w2 => d30_in(8*N-1 downto 7*N),w3 => d30_in(7*N-1 downto 6*N),w4 => d30_in(6*N-1 downto 5*N),w5 => d30_in(5*N-1 downto 4*N),w6 => d30_in(4*N-1 downto 3*N),w7 => d30_in(3*N-1 downto 2*N),w8 => d30_in(2*N-1 downto N),w9 => d30_in(N-1 downto 0 ),d_out => d30_out,en_out =>open  ,sof_out=>open   );
CL31: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d31_in(9*N-1 downto 8*N),data2conv2 =>d31_in(8*N-1 downto 7*N),data2conv3 =>d31_in(7*N-1 downto 6*N),data2conv4 =>d31_in(6*N-1 downto 5*N),data2conv5 =>d31_in(5*N-1 downto 4*N),data2conv6 =>d31_in(4*N-1 downto 3*N),data2conv7 =>d31_in(3*N-1 downto 2*N),data2conv8 =>d31_in(2*N-1 downto N),data2conv9 =>d31_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d31_in(9*N-1 downto 8*N),w2 => d31_in(8*N-1 downto 7*N),w3 => d31_in(7*N-1 downto 6*N),w4 => d31_in(6*N-1 downto 5*N),w5 => d31_in(5*N-1 downto 4*N),w6 => d31_in(4*N-1 downto 3*N),w7 => d31_in(3*N-1 downto 2*N),w8 => d31_in(2*N-1 downto N),w9 => d31_in(N-1 downto 0 ),d_out => d31_out,en_out =>open  ,sof_out=>open   );
CL32: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d32_in(9*N-1 downto 8*N),data2conv2 =>d32_in(8*N-1 downto 7*N),data2conv3 =>d32_in(7*N-1 downto 6*N),data2conv4 =>d32_in(6*N-1 downto 5*N),data2conv5 =>d32_in(5*N-1 downto 4*N),data2conv6 =>d32_in(4*N-1 downto 3*N),data2conv7 =>d32_in(3*N-1 downto 2*N),data2conv8 =>d32_in(2*N-1 downto N),data2conv9 =>d32_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d32_in(9*N-1 downto 8*N),w2 => d32_in(8*N-1 downto 7*N),w3 => d32_in(7*N-1 downto 6*N),w4 => d32_in(6*N-1 downto 5*N),w5 => d32_in(5*N-1 downto 4*N),w6 => d32_in(4*N-1 downto 3*N),w7 => d32_in(3*N-1 downto 2*N),w8 => d32_in(2*N-1 downto N),w9 => d32_in(N-1 downto 0 ),d_out => d32_out,en_out =>open  ,sof_out=>open   );
CL33: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d33_in(9*N-1 downto 8*N),data2conv2 =>d33_in(8*N-1 downto 7*N),data2conv3 =>d33_in(7*N-1 downto 6*N),data2conv4 =>d33_in(6*N-1 downto 5*N),data2conv5 =>d33_in(5*N-1 downto 4*N),data2conv6 =>d33_in(4*N-1 downto 3*N),data2conv7 =>d33_in(3*N-1 downto 2*N),data2conv8 =>d33_in(2*N-1 downto N),data2conv9 =>d33_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d33_in(9*N-1 downto 8*N),w2 => d33_in(8*N-1 downto 7*N),w3 => d33_in(7*N-1 downto 6*N),w4 => d33_in(6*N-1 downto 5*N),w5 => d33_in(5*N-1 downto 4*N),w6 => d33_in(4*N-1 downto 3*N),w7 => d33_in(3*N-1 downto 2*N),w8 => d33_in(2*N-1 downto N),w9 => d33_in(N-1 downto 0 ),d_out => d33_out,en_out =>open  ,sof_out=>open   );
CL34: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d34_in(9*N-1 downto 8*N),data2conv2 =>d34_in(8*N-1 downto 7*N),data2conv3 =>d34_in(7*N-1 downto 6*N),data2conv4 =>d34_in(6*N-1 downto 5*N),data2conv5 =>d34_in(5*N-1 downto 4*N),data2conv6 =>d34_in(4*N-1 downto 3*N),data2conv7 =>d34_in(3*N-1 downto 2*N),data2conv8 =>d34_in(2*N-1 downto N),data2conv9 =>d34_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d34_in(9*N-1 downto 8*N),w2 => d34_in(8*N-1 downto 7*N),w3 => d34_in(7*N-1 downto 6*N),w4 => d34_in(6*N-1 downto 5*N),w5 => d34_in(5*N-1 downto 4*N),w6 => d34_in(4*N-1 downto 3*N),w7 => d34_in(3*N-1 downto 2*N),w8 => d34_in(2*N-1 downto N),w9 => d34_in(N-1 downto 0 ),d_out => d34_out,en_out =>open  ,sof_out=>open   );
CL35: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d35_in(9*N-1 downto 8*N),data2conv2 =>d35_in(8*N-1 downto 7*N),data2conv3 =>d35_in(7*N-1 downto 6*N),data2conv4 =>d35_in(6*N-1 downto 5*N),data2conv5 =>d35_in(5*N-1 downto 4*N),data2conv6 =>d35_in(4*N-1 downto 3*N),data2conv7 =>d35_in(3*N-1 downto 2*N),data2conv8 =>d35_in(2*N-1 downto N),data2conv9 =>d35_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d35_in(9*N-1 downto 8*N),w2 => d35_in(8*N-1 downto 7*N),w3 => d35_in(7*N-1 downto 6*N),w4 => d35_in(6*N-1 downto 5*N),w5 => d35_in(5*N-1 downto 4*N),w6 => d35_in(4*N-1 downto 3*N),w7 => d35_in(3*N-1 downto 2*N),w8 => d35_in(2*N-1 downto N),w9 => d35_in(N-1 downto 0 ),d_out => d35_out,en_out =>open  ,sof_out=>open   );
CL36: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d36_in(9*N-1 downto 8*N),data2conv2 =>d36_in(8*N-1 downto 7*N),data2conv3 =>d36_in(7*N-1 downto 6*N),data2conv4 =>d36_in(6*N-1 downto 5*N),data2conv5 =>d36_in(5*N-1 downto 4*N),data2conv6 =>d36_in(4*N-1 downto 3*N),data2conv7 =>d36_in(3*N-1 downto 2*N),data2conv8 =>d36_in(2*N-1 downto N),data2conv9 =>d36_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d36_in(9*N-1 downto 8*N),w2 => d36_in(8*N-1 downto 7*N),w3 => d36_in(7*N-1 downto 6*N),w4 => d36_in(6*N-1 downto 5*N),w5 => d36_in(5*N-1 downto 4*N),w6 => d36_in(4*N-1 downto 3*N),w7 => d36_in(3*N-1 downto 2*N),w8 => d36_in(2*N-1 downto N),w9 => d36_in(N-1 downto 0 ),d_out => d36_out,en_out =>open  ,sof_out=>open   );
CL37: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d37_in(9*N-1 downto 8*N),data2conv2 =>d37_in(8*N-1 downto 7*N),data2conv3 =>d37_in(7*N-1 downto 6*N),data2conv4 =>d37_in(6*N-1 downto 5*N),data2conv5 =>d37_in(5*N-1 downto 4*N),data2conv6 =>d37_in(4*N-1 downto 3*N),data2conv7 =>d37_in(3*N-1 downto 2*N),data2conv8 =>d37_in(2*N-1 downto N),data2conv9 =>d37_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d37_in(9*N-1 downto 8*N),w2 => d37_in(8*N-1 downto 7*N),w3 => d37_in(7*N-1 downto 6*N),w4 => d37_in(6*N-1 downto 5*N),w5 => d37_in(5*N-1 downto 4*N),w6 => d37_in(4*N-1 downto 3*N),w7 => d37_in(3*N-1 downto 2*N),w8 => d37_in(2*N-1 downto N),w9 => d37_in(N-1 downto 0 ),d_out => d37_out,en_out =>open  ,sof_out=>open   );
CL38: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d38_in(9*N-1 downto 8*N),data2conv2 =>d38_in(8*N-1 downto 7*N),data2conv3 =>d38_in(7*N-1 downto 6*N),data2conv4 =>d38_in(6*N-1 downto 5*N),data2conv5 =>d38_in(5*N-1 downto 4*N),data2conv6 =>d38_in(4*N-1 downto 3*N),data2conv7 =>d38_in(3*N-1 downto 2*N),data2conv8 =>d38_in(2*N-1 downto N),data2conv9 =>d38_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d38_in(9*N-1 downto 8*N),w2 => d38_in(8*N-1 downto 7*N),w3 => d38_in(7*N-1 downto 6*N),w4 => d38_in(6*N-1 downto 5*N),w5 => d38_in(5*N-1 downto 4*N),w6 => d38_in(4*N-1 downto 3*N),w7 => d38_in(3*N-1 downto 2*N),w8 => d38_in(2*N-1 downto N),w9 => d38_in(N-1 downto 0 ),d_out => d38_out,en_out =>open  ,sof_out=>open   );
CL39: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d39_in(9*N-1 downto 8*N),data2conv2 =>d39_in(8*N-1 downto 7*N),data2conv3 =>d39_in(7*N-1 downto 6*N),data2conv4 =>d39_in(6*N-1 downto 5*N),data2conv5 =>d39_in(5*N-1 downto 4*N),data2conv6 =>d39_in(4*N-1 downto 3*N),data2conv7 =>d39_in(3*N-1 downto 2*N),data2conv8 =>d39_in(2*N-1 downto N),data2conv9 =>d39_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d39_in(9*N-1 downto 8*N),w2 => d39_in(8*N-1 downto 7*N),w3 => d39_in(7*N-1 downto 6*N),w4 => d39_in(6*N-1 downto 5*N),w5 => d39_in(5*N-1 downto 4*N),w6 => d39_in(4*N-1 downto 3*N),w7 => d39_in(3*N-1 downto 2*N),w8 => d39_in(2*N-1 downto N),w9 => d39_in(N-1 downto 0 ),d_out => d39_out,en_out =>open  ,sof_out=>open   );
CL40: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d40_in(9*N-1 downto 8*N),data2conv2 =>d40_in(8*N-1 downto 7*N),data2conv3 =>d40_in(7*N-1 downto 6*N),data2conv4 =>d40_in(6*N-1 downto 5*N),data2conv5 =>d40_in(5*N-1 downto 4*N),data2conv6 =>d40_in(4*N-1 downto 3*N),data2conv7 =>d40_in(3*N-1 downto 2*N),data2conv8 =>d40_in(2*N-1 downto N),data2conv9 =>d40_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d40_in(9*N-1 downto 8*N),w2 => d40_in(8*N-1 downto 7*N),w3 => d40_in(7*N-1 downto 6*N),w4 => d40_in(6*N-1 downto 5*N),w5 => d40_in(5*N-1 downto 4*N),w6 => d40_in(4*N-1 downto 3*N),w7 => d40_in(3*N-1 downto 2*N),w8 => d40_in(2*N-1 downto N),w9 => d40_in(N-1 downto 0 ),d_out => d40_out,en_out =>open  ,sof_out=>open   );
CL41: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d41_in(9*N-1 downto 8*N),data2conv2 =>d41_in(8*N-1 downto 7*N),data2conv3 =>d41_in(7*N-1 downto 6*N),data2conv4 =>d41_in(6*N-1 downto 5*N),data2conv5 =>d41_in(5*N-1 downto 4*N),data2conv6 =>d41_in(4*N-1 downto 3*N),data2conv7 =>d41_in(3*N-1 downto 2*N),data2conv8 =>d41_in(2*N-1 downto N),data2conv9 =>d41_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d41_in(9*N-1 downto 8*N),w2 => d41_in(8*N-1 downto 7*N),w3 => d41_in(7*N-1 downto 6*N),w4 => d41_in(6*N-1 downto 5*N),w5 => d41_in(5*N-1 downto 4*N),w6 => d41_in(4*N-1 downto 3*N),w7 => d41_in(3*N-1 downto 2*N),w8 => d41_in(2*N-1 downto N),w9 => d41_in(N-1 downto 0 ),d_out => d41_out,en_out =>open  ,sof_out=>open   );
CL42: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d42_in(9*N-1 downto 8*N),data2conv2 =>d42_in(8*N-1 downto 7*N),data2conv3 =>d42_in(7*N-1 downto 6*N),data2conv4 =>d42_in(6*N-1 downto 5*N),data2conv5 =>d42_in(5*N-1 downto 4*N),data2conv6 =>d42_in(4*N-1 downto 3*N),data2conv7 =>d42_in(3*N-1 downto 2*N),data2conv8 =>d42_in(2*N-1 downto N),data2conv9 =>d42_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d42_in(9*N-1 downto 8*N),w2 => d42_in(8*N-1 downto 7*N),w3 => d42_in(7*N-1 downto 6*N),w4 => d42_in(6*N-1 downto 5*N),w5 => d42_in(5*N-1 downto 4*N),w6 => d42_in(4*N-1 downto 3*N),w7 => d42_in(3*N-1 downto 2*N),w8 => d42_in(2*N-1 downto N),w9 => d42_in(N-1 downto 0 ),d_out => d42_out,en_out =>open  ,sof_out=>open   );
CL43: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d43_in(9*N-1 downto 8*N),data2conv2 =>d43_in(8*N-1 downto 7*N),data2conv3 =>d43_in(7*N-1 downto 6*N),data2conv4 =>d43_in(6*N-1 downto 5*N),data2conv5 =>d43_in(5*N-1 downto 4*N),data2conv6 =>d43_in(4*N-1 downto 3*N),data2conv7 =>d43_in(3*N-1 downto 2*N),data2conv8 =>d43_in(2*N-1 downto N),data2conv9 =>d43_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d43_in(9*N-1 downto 8*N),w2 => d43_in(8*N-1 downto 7*N),w3 => d43_in(7*N-1 downto 6*N),w4 => d43_in(6*N-1 downto 5*N),w5 => d43_in(5*N-1 downto 4*N),w6 => d43_in(4*N-1 downto 3*N),w7 => d43_in(3*N-1 downto 2*N),w8 => d43_in(2*N-1 downto N),w9 => d43_in(N-1 downto 0 ),d_out => d43_out,en_out =>open  ,sof_out=>open   );
CL44: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d44_in(9*N-1 downto 8*N),data2conv2 =>d44_in(8*N-1 downto 7*N),data2conv3 =>d44_in(7*N-1 downto 6*N),data2conv4 =>d44_in(6*N-1 downto 5*N),data2conv5 =>d44_in(5*N-1 downto 4*N),data2conv6 =>d44_in(4*N-1 downto 3*N),data2conv7 =>d44_in(3*N-1 downto 2*N),data2conv8 =>d44_in(2*N-1 downto N),data2conv9 =>d44_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d44_in(9*N-1 downto 8*N),w2 => d44_in(8*N-1 downto 7*N),w3 => d44_in(7*N-1 downto 6*N),w4 => d44_in(6*N-1 downto 5*N),w5 => d44_in(5*N-1 downto 4*N),w6 => d44_in(4*N-1 downto 3*N),w7 => d44_in(3*N-1 downto 2*N),w8 => d44_in(2*N-1 downto N),w9 => d44_in(N-1 downto 0 ),d_out => d44_out,en_out =>open  ,sof_out=>open   );
CL45: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d45_in(9*N-1 downto 8*N),data2conv2 =>d45_in(8*N-1 downto 7*N),data2conv3 =>d45_in(7*N-1 downto 6*N),data2conv4 =>d45_in(6*N-1 downto 5*N),data2conv5 =>d45_in(5*N-1 downto 4*N),data2conv6 =>d45_in(4*N-1 downto 3*N),data2conv7 =>d45_in(3*N-1 downto 2*N),data2conv8 =>d45_in(2*N-1 downto N),data2conv9 =>d45_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d45_in(9*N-1 downto 8*N),w2 => d45_in(8*N-1 downto 7*N),w3 => d45_in(7*N-1 downto 6*N),w4 => d45_in(6*N-1 downto 5*N),w5 => d45_in(5*N-1 downto 4*N),w6 => d45_in(4*N-1 downto 3*N),w7 => d45_in(3*N-1 downto 2*N),w8 => d45_in(2*N-1 downto N),w9 => d45_in(N-1 downto 0 ),d_out => d45_out,en_out =>open  ,sof_out=>open   );
CL46: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d46_in(9*N-1 downto 8*N),data2conv2 =>d46_in(8*N-1 downto 7*N),data2conv3 =>d46_in(7*N-1 downto 6*N),data2conv4 =>d46_in(6*N-1 downto 5*N),data2conv5 =>d46_in(5*N-1 downto 4*N),data2conv6 =>d46_in(4*N-1 downto 3*N),data2conv7 =>d46_in(3*N-1 downto 2*N),data2conv8 =>d46_in(2*N-1 downto N),data2conv9 =>d46_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d46_in(9*N-1 downto 8*N),w2 => d46_in(8*N-1 downto 7*N),w3 => d46_in(7*N-1 downto 6*N),w4 => d46_in(6*N-1 downto 5*N),w5 => d46_in(5*N-1 downto 4*N),w6 => d46_in(4*N-1 downto 3*N),w7 => d46_in(3*N-1 downto 2*N),w8 => d46_in(2*N-1 downto N),w9 => d46_in(N-1 downto 0 ),d_out => d46_out,en_out =>open  ,sof_out=>open   );
CL47: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d47_in(9*N-1 downto 8*N),data2conv2 =>d47_in(8*N-1 downto 7*N),data2conv3 =>d47_in(7*N-1 downto 6*N),data2conv4 =>d47_in(6*N-1 downto 5*N),data2conv5 =>d47_in(5*N-1 downto 4*N),data2conv6 =>d47_in(4*N-1 downto 3*N),data2conv7 =>d47_in(3*N-1 downto 2*N),data2conv8 =>d47_in(2*N-1 downto N),data2conv9 =>d47_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d47_in(9*N-1 downto 8*N),w2 => d47_in(8*N-1 downto 7*N),w3 => d47_in(7*N-1 downto 6*N),w4 => d47_in(6*N-1 downto 5*N),w5 => d47_in(5*N-1 downto 4*N),w6 => d47_in(4*N-1 downto 3*N),w7 => d47_in(3*N-1 downto 2*N),w8 => d47_in(2*N-1 downto N),w9 => d47_in(N-1 downto 0 ),d_out => d47_out,en_out =>open  ,sof_out=>open   );
CL48: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d48_in(9*N-1 downto 8*N),data2conv2 =>d48_in(8*N-1 downto 7*N),data2conv3 =>d48_in(7*N-1 downto 6*N),data2conv4 =>d48_in(6*N-1 downto 5*N),data2conv5 =>d48_in(5*N-1 downto 4*N),data2conv6 =>d48_in(4*N-1 downto 3*N),data2conv7 =>d48_in(3*N-1 downto 2*N),data2conv8 =>d48_in(2*N-1 downto N),data2conv9 =>d48_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d48_in(9*N-1 downto 8*N),w2 => d48_in(8*N-1 downto 7*N),w3 => d48_in(7*N-1 downto 6*N),w4 => d48_in(6*N-1 downto 5*N),w5 => d48_in(5*N-1 downto 4*N),w6 => d48_in(4*N-1 downto 3*N),w7 => d48_in(3*N-1 downto 2*N),w8 => d48_in(2*N-1 downto N),w9 => d48_in(N-1 downto 0 ),d_out => d48_out,en_out =>open  ,sof_out=>open   );
CL49: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d49_in(9*N-1 downto 8*N),data2conv2 =>d49_in(8*N-1 downto 7*N),data2conv3 =>d49_in(7*N-1 downto 6*N),data2conv4 =>d49_in(6*N-1 downto 5*N),data2conv5 =>d49_in(5*N-1 downto 4*N),data2conv6 =>d49_in(4*N-1 downto 3*N),data2conv7 =>d49_in(3*N-1 downto 2*N),data2conv8 =>d49_in(2*N-1 downto N),data2conv9 =>d49_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d49_in(9*N-1 downto 8*N),w2 => d49_in(8*N-1 downto 7*N),w3 => d49_in(7*N-1 downto 6*N),w4 => d49_in(6*N-1 downto 5*N),w5 => d49_in(5*N-1 downto 4*N),w6 => d49_in(4*N-1 downto 3*N),w7 => d49_in(3*N-1 downto 2*N),w8 => d49_in(2*N-1 downto N),w9 => d49_in(N-1 downto 0 ),d_out => d49_out,en_out =>open  ,sof_out=>open   );
CL50: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d50_in(9*N-1 downto 8*N),data2conv2 =>d50_in(8*N-1 downto 7*N),data2conv3 =>d50_in(7*N-1 downto 6*N),data2conv4 =>d50_in(6*N-1 downto 5*N),data2conv5 =>d50_in(5*N-1 downto 4*N),data2conv6 =>d50_in(4*N-1 downto 3*N),data2conv7 =>d50_in(3*N-1 downto 2*N),data2conv8 =>d50_in(2*N-1 downto N),data2conv9 =>d50_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d50_in(9*N-1 downto 8*N),w2 => d50_in(8*N-1 downto 7*N),w3 => d50_in(7*N-1 downto 6*N),w4 => d50_in(6*N-1 downto 5*N),w5 => d50_in(5*N-1 downto 4*N),w6 => d50_in(4*N-1 downto 3*N),w7 => d50_in(3*N-1 downto 2*N),w8 => d50_in(2*N-1 downto N),w9 => d50_in(N-1 downto 0 ),d_out => d50_out,en_out =>open  ,sof_out=>open   );
CL51: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d51_in(9*N-1 downto 8*N),data2conv2 =>d51_in(8*N-1 downto 7*N),data2conv3 =>d51_in(7*N-1 downto 6*N),data2conv4 =>d51_in(6*N-1 downto 5*N),data2conv5 =>d51_in(5*N-1 downto 4*N),data2conv6 =>d51_in(4*N-1 downto 3*N),data2conv7 =>d51_in(3*N-1 downto 2*N),data2conv8 =>d51_in(2*N-1 downto N),data2conv9 =>d51_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d51_in(9*N-1 downto 8*N),w2 => d51_in(8*N-1 downto 7*N),w3 => d51_in(7*N-1 downto 6*N),w4 => d51_in(6*N-1 downto 5*N),w5 => d51_in(5*N-1 downto 4*N),w6 => d51_in(4*N-1 downto 3*N),w7 => d51_in(3*N-1 downto 2*N),w8 => d51_in(2*N-1 downto N),w9 => d51_in(N-1 downto 0 ),d_out => d51_out,en_out =>open  ,sof_out=>open   );
CL52: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d52_in(9*N-1 downto 8*N),data2conv2 =>d52_in(8*N-1 downto 7*N),data2conv3 =>d52_in(7*N-1 downto 6*N),data2conv4 =>d52_in(6*N-1 downto 5*N),data2conv5 =>d52_in(5*N-1 downto 4*N),data2conv6 =>d52_in(4*N-1 downto 3*N),data2conv7 =>d52_in(3*N-1 downto 2*N),data2conv8 =>d52_in(2*N-1 downto N),data2conv9 =>d52_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d52_in(9*N-1 downto 8*N),w2 => d52_in(8*N-1 downto 7*N),w3 => d52_in(7*N-1 downto 6*N),w4 => d52_in(6*N-1 downto 5*N),w5 => d52_in(5*N-1 downto 4*N),w6 => d52_in(4*N-1 downto 3*N),w7 => d52_in(3*N-1 downto 2*N),w8 => d52_in(2*N-1 downto N),w9 => d52_in(N-1 downto 0 ),d_out => d52_out,en_out =>open  ,sof_out=>open   );
CL53: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d53_in(9*N-1 downto 8*N),data2conv2 =>d53_in(8*N-1 downto 7*N),data2conv3 =>d53_in(7*N-1 downto 6*N),data2conv4 =>d53_in(6*N-1 downto 5*N),data2conv5 =>d53_in(5*N-1 downto 4*N),data2conv6 =>d53_in(4*N-1 downto 3*N),data2conv7 =>d53_in(3*N-1 downto 2*N),data2conv8 =>d53_in(2*N-1 downto N),data2conv9 =>d53_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d53_in(9*N-1 downto 8*N),w2 => d53_in(8*N-1 downto 7*N),w3 => d53_in(7*N-1 downto 6*N),w4 => d53_in(6*N-1 downto 5*N),w5 => d53_in(5*N-1 downto 4*N),w6 => d53_in(4*N-1 downto 3*N),w7 => d53_in(3*N-1 downto 2*N),w8 => d53_in(2*N-1 downto N),w9 => d53_in(N-1 downto 0 ),d_out => d53_out,en_out =>open  ,sof_out=>open   );
CL54: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d54_in(9*N-1 downto 8*N),data2conv2 =>d54_in(8*N-1 downto 7*N),data2conv3 =>d54_in(7*N-1 downto 6*N),data2conv4 =>d54_in(6*N-1 downto 5*N),data2conv5 =>d54_in(5*N-1 downto 4*N),data2conv6 =>d54_in(4*N-1 downto 3*N),data2conv7 =>d54_in(3*N-1 downto 2*N),data2conv8 =>d54_in(2*N-1 downto N),data2conv9 =>d54_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d54_in(9*N-1 downto 8*N),w2 => d54_in(8*N-1 downto 7*N),w3 => d54_in(7*N-1 downto 6*N),w4 => d54_in(6*N-1 downto 5*N),w5 => d54_in(5*N-1 downto 4*N),w6 => d54_in(4*N-1 downto 3*N),w7 => d54_in(3*N-1 downto 2*N),w8 => d54_in(2*N-1 downto N),w9 => d54_in(N-1 downto 0 ),d_out => d54_out,en_out =>open  ,sof_out=>open   );
CL55: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d55_in(9*N-1 downto 8*N),data2conv2 =>d55_in(8*N-1 downto 7*N),data2conv3 =>d55_in(7*N-1 downto 6*N),data2conv4 =>d55_in(6*N-1 downto 5*N),data2conv5 =>d55_in(5*N-1 downto 4*N),data2conv6 =>d55_in(4*N-1 downto 3*N),data2conv7 =>d55_in(3*N-1 downto 2*N),data2conv8 =>d55_in(2*N-1 downto N),data2conv9 =>d55_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d55_in(9*N-1 downto 8*N),w2 => d55_in(8*N-1 downto 7*N),w3 => d55_in(7*N-1 downto 6*N),w4 => d55_in(6*N-1 downto 5*N),w5 => d55_in(5*N-1 downto 4*N),w6 => d55_in(4*N-1 downto 3*N),w7 => d55_in(3*N-1 downto 2*N),w8 => d55_in(2*N-1 downto N),w9 => d55_in(N-1 downto 0 ),d_out => d55_out,en_out =>open  ,sof_out=>open   );
CL56: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d56_in(9*N-1 downto 8*N),data2conv2 =>d56_in(8*N-1 downto 7*N),data2conv3 =>d56_in(7*N-1 downto 6*N),data2conv4 =>d56_in(6*N-1 downto 5*N),data2conv5 =>d56_in(5*N-1 downto 4*N),data2conv6 =>d56_in(4*N-1 downto 3*N),data2conv7 =>d56_in(3*N-1 downto 2*N),data2conv8 =>d56_in(2*N-1 downto N),data2conv9 =>d56_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d56_in(9*N-1 downto 8*N),w2 => d56_in(8*N-1 downto 7*N),w3 => d56_in(7*N-1 downto 6*N),w4 => d56_in(6*N-1 downto 5*N),w5 => d56_in(5*N-1 downto 4*N),w6 => d56_in(4*N-1 downto 3*N),w7 => d56_in(3*N-1 downto 2*N),w8 => d56_in(2*N-1 downto N),w9 => d56_in(N-1 downto 0 ),d_out => d56_out,en_out =>open  ,sof_out=>open   );
CL57: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d57_in(9*N-1 downto 8*N),data2conv2 =>d57_in(8*N-1 downto 7*N),data2conv3 =>d57_in(7*N-1 downto 6*N),data2conv4 =>d57_in(6*N-1 downto 5*N),data2conv5 =>d57_in(5*N-1 downto 4*N),data2conv6 =>d57_in(4*N-1 downto 3*N),data2conv7 =>d57_in(3*N-1 downto 2*N),data2conv8 =>d57_in(2*N-1 downto N),data2conv9 =>d57_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d57_in(9*N-1 downto 8*N),w2 => d57_in(8*N-1 downto 7*N),w3 => d57_in(7*N-1 downto 6*N),w4 => d57_in(6*N-1 downto 5*N),w5 => d57_in(5*N-1 downto 4*N),w6 => d57_in(4*N-1 downto 3*N),w7 => d57_in(3*N-1 downto 2*N),w8 => d57_in(2*N-1 downto N),w9 => d57_in(N-1 downto 0 ),d_out => d57_out,en_out =>open  ,sof_out=>open   );
CL58: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d58_in(9*N-1 downto 8*N),data2conv2 =>d58_in(8*N-1 downto 7*N),data2conv3 =>d58_in(7*N-1 downto 6*N),data2conv4 =>d58_in(6*N-1 downto 5*N),data2conv5 =>d58_in(5*N-1 downto 4*N),data2conv6 =>d58_in(4*N-1 downto 3*N),data2conv7 =>d58_in(3*N-1 downto 2*N),data2conv8 =>d58_in(2*N-1 downto N),data2conv9 =>d58_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d58_in(9*N-1 downto 8*N),w2 => d58_in(8*N-1 downto 7*N),w3 => d58_in(7*N-1 downto 6*N),w4 => d58_in(6*N-1 downto 5*N),w5 => d58_in(5*N-1 downto 4*N),w6 => d58_in(4*N-1 downto 3*N),w7 => d58_in(3*N-1 downto 2*N),w8 => d58_in(2*N-1 downto N),w9 => d58_in(N-1 downto 0 ),d_out => d58_out,en_out =>open  ,sof_out=>open   );
CL59: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d59_in(9*N-1 downto 8*N),data2conv2 =>d59_in(8*N-1 downto 7*N),data2conv3 =>d59_in(7*N-1 downto 6*N),data2conv4 =>d59_in(6*N-1 downto 5*N),data2conv5 =>d59_in(5*N-1 downto 4*N),data2conv6 =>d59_in(4*N-1 downto 3*N),data2conv7 =>d59_in(3*N-1 downto 2*N),data2conv8 =>d59_in(2*N-1 downto N),data2conv9 =>d59_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d59_in(9*N-1 downto 8*N),w2 => d59_in(8*N-1 downto 7*N),w3 => d59_in(7*N-1 downto 6*N),w4 => d59_in(6*N-1 downto 5*N),w5 => d59_in(5*N-1 downto 4*N),w6 => d59_in(4*N-1 downto 3*N),w7 => d59_in(3*N-1 downto 2*N),w8 => d59_in(2*N-1 downto N),w9 => d59_in(N-1 downto 0 ),d_out => d59_out,en_out =>open  ,sof_out=>open   );
CL60: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d60_in(9*N-1 downto 8*N),data2conv2 =>d60_in(8*N-1 downto 7*N),data2conv3 =>d60_in(7*N-1 downto 6*N),data2conv4 =>d60_in(6*N-1 downto 5*N),data2conv5 =>d60_in(5*N-1 downto 4*N),data2conv6 =>d60_in(4*N-1 downto 3*N),data2conv7 =>d60_in(3*N-1 downto 2*N),data2conv8 =>d60_in(2*N-1 downto N),data2conv9 =>d60_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d60_in(9*N-1 downto 8*N),w2 => d60_in(8*N-1 downto 7*N),w3 => d60_in(7*N-1 downto 6*N),w4 => d60_in(6*N-1 downto 5*N),w5 => d60_in(5*N-1 downto 4*N),w6 => d60_in(4*N-1 downto 3*N),w7 => d60_in(3*N-1 downto 2*N),w8 => d60_in(2*N-1 downto N),w9 => d60_in(N-1 downto 0 ),d_out => d60_out,en_out =>open  ,sof_out=>open   );
CL61: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d61_in(9*N-1 downto 8*N),data2conv2 =>d61_in(8*N-1 downto 7*N),data2conv3 =>d61_in(7*N-1 downto 6*N),data2conv4 =>d61_in(6*N-1 downto 5*N),data2conv5 =>d61_in(5*N-1 downto 4*N),data2conv6 =>d61_in(4*N-1 downto 3*N),data2conv7 =>d61_in(3*N-1 downto 2*N),data2conv8 =>d61_in(2*N-1 downto N),data2conv9 =>d61_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d61_in(9*N-1 downto 8*N),w2 => d61_in(8*N-1 downto 7*N),w3 => d61_in(7*N-1 downto 6*N),w4 => d61_in(6*N-1 downto 5*N),w5 => d61_in(5*N-1 downto 4*N),w6 => d61_in(4*N-1 downto 3*N),w7 => d61_in(3*N-1 downto 2*N),w8 => d61_in(2*N-1 downto N),w9 => d61_in(N-1 downto 0 ),d_out => d61_out,en_out =>open  ,sof_out=>open   );
CL62: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d62_in(9*N-1 downto 8*N),data2conv2 =>d62_in(8*N-1 downto 7*N),data2conv3 =>d62_in(7*N-1 downto 6*N),data2conv4 =>d62_in(6*N-1 downto 5*N),data2conv5 =>d62_in(5*N-1 downto 4*N),data2conv6 =>d62_in(4*N-1 downto 3*N),data2conv7 =>d62_in(3*N-1 downto 2*N),data2conv8 =>d62_in(2*N-1 downto N),data2conv9 =>d62_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d62_in(9*N-1 downto 8*N),w2 => d62_in(8*N-1 downto 7*N),w3 => d62_in(7*N-1 downto 6*N),w4 => d62_in(6*N-1 downto 5*N),w5 => d62_in(5*N-1 downto 4*N),w6 => d62_in(4*N-1 downto 3*N),w7 => d62_in(3*N-1 downto 2*N),w8 => d62_in(2*N-1 downto N),w9 => d62_in(N-1 downto 0 ),d_out => d62_out,en_out =>open  ,sof_out=>open   );
CL63: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d63_in(9*N-1 downto 8*N),data2conv2 =>d63_in(8*N-1 downto 7*N),data2conv3 =>d63_in(7*N-1 downto 6*N),data2conv4 =>d63_in(6*N-1 downto 5*N),data2conv5 =>d63_in(5*N-1 downto 4*N),data2conv6 =>d63_in(4*N-1 downto 3*N),data2conv7 =>d63_in(3*N-1 downto 2*N),data2conv8 =>d63_in(2*N-1 downto N),data2conv9 =>d63_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d63_in(9*N-1 downto 8*N),w2 => d63_in(8*N-1 downto 7*N),w3 => d63_in(7*N-1 downto 6*N),w4 => d63_in(6*N-1 downto 5*N),w5 => d63_in(5*N-1 downto 4*N),w6 => d63_in(4*N-1 downto 3*N),w7 => d63_in(3*N-1 downto 2*N),w8 => d63_in(2*N-1 downto N),w9 => d63_in(N-1 downto 0 ),d_out => d63_out,en_out =>open  ,sof_out=>open   );
CL64: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d64_in(9*N-1 downto 8*N),data2conv2 =>d64_in(8*N-1 downto 7*N),data2conv3 =>d64_in(7*N-1 downto 6*N),data2conv4 =>d64_in(6*N-1 downto 5*N),data2conv5 =>d64_in(5*N-1 downto 4*N),data2conv6 =>d64_in(4*N-1 downto 3*N),data2conv7 =>d64_in(3*N-1 downto 2*N),data2conv8 =>d64_in(2*N-1 downto N),data2conv9 =>d64_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d64_in(9*N-1 downto 8*N),w2 => d64_in(8*N-1 downto 7*N),w3 => d64_in(7*N-1 downto 6*N),w4 => d64_in(6*N-1 downto 5*N),w5 => d64_in(5*N-1 downto 4*N),w6 => d64_in(4*N-1 downto 3*N),w7 => d64_in(3*N-1 downto 2*N),w8 => d64_in(2*N-1 downto N),w9 => d64_in(N-1 downto 0 ),d_out => d64_out,en_out =>open  ,sof_out=>open   );

CL65 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d65_in (9*N-1 downto 8*N),data2conv2 =>d65_in (8*N-1 downto 7*N),data2conv3 =>d65_in (7*N-1 downto 6*N),data2conv4 =>d65_in (6*N-1 downto 5*N),data2conv5 =>d65_in (5*N-1 downto 4*N),data2conv6 =>d65_in (4*N-1 downto 3*N),data2conv7 =>d65_in (3*N-1 downto 2*N),data2conv8 =>d65_in (2*N-1 downto N),data2conv9 =>d65_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d65_in (9*N-1 downto 8*N),w2 => d65_in (8*N-1 downto 7*N),w3 => d65_in (7*N-1 downto 6*N),w4 => d65_in (6*N-1 downto 5*N),w5 => d65_in (5*N-1 downto 4*N),w6 => d65_in (4*N-1 downto 3*N),w7 => d65_in (3*N-1 downto 2*N),w8 => d65_in (2*N-1 downto N),w9 => d65_in (N-1 downto 0 ),d_out => d65_out ,en_out =>open  ,sof_out=>open   );
CL66 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d66_in (9*N-1 downto 8*N),data2conv2 =>d66_in (8*N-1 downto 7*N),data2conv3 =>d66_in (7*N-1 downto 6*N),data2conv4 =>d66_in (6*N-1 downto 5*N),data2conv5 =>d66_in (5*N-1 downto 4*N),data2conv6 =>d66_in (4*N-1 downto 3*N),data2conv7 =>d66_in (3*N-1 downto 2*N),data2conv8 =>d66_in (2*N-1 downto N),data2conv9 =>d66_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d66_in (9*N-1 downto 8*N),w2 => d66_in (8*N-1 downto 7*N),w3 => d66_in (7*N-1 downto 6*N),w4 => d66_in (6*N-1 downto 5*N),w5 => d66_in (5*N-1 downto 4*N),w6 => d66_in (4*N-1 downto 3*N),w7 => d66_in (3*N-1 downto 2*N),w8 => d66_in (2*N-1 downto N),w9 => d66_in (N-1 downto 0 ),d_out => d66_out ,en_out =>open  ,sof_out=>open   );
CL67 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d67_in (9*N-1 downto 8*N),data2conv2 =>d67_in (8*N-1 downto 7*N),data2conv3 =>d67_in (7*N-1 downto 6*N),data2conv4 =>d67_in (6*N-1 downto 5*N),data2conv5 =>d67_in (5*N-1 downto 4*N),data2conv6 =>d67_in (4*N-1 downto 3*N),data2conv7 =>d67_in (3*N-1 downto 2*N),data2conv8 =>d67_in (2*N-1 downto N),data2conv9 =>d67_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d67_in (9*N-1 downto 8*N),w2 => d67_in (8*N-1 downto 7*N),w3 => d67_in (7*N-1 downto 6*N),w4 => d67_in (6*N-1 downto 5*N),w5 => d67_in (5*N-1 downto 4*N),w6 => d67_in (4*N-1 downto 3*N),w7 => d67_in (3*N-1 downto 2*N),w8 => d67_in (2*N-1 downto N),w9 => d67_in (N-1 downto 0 ),d_out => d67_out ,en_out =>open  ,sof_out=>open   );
CL68 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d68_in (9*N-1 downto 8*N),data2conv2 =>d68_in (8*N-1 downto 7*N),data2conv3 =>d68_in (7*N-1 downto 6*N),data2conv4 =>d68_in (6*N-1 downto 5*N),data2conv5 =>d68_in (5*N-1 downto 4*N),data2conv6 =>d68_in (4*N-1 downto 3*N),data2conv7 =>d68_in (3*N-1 downto 2*N),data2conv8 =>d68_in (2*N-1 downto N),data2conv9 =>d68_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d68_in (9*N-1 downto 8*N),w2 => d68_in (8*N-1 downto 7*N),w3 => d68_in (7*N-1 downto 6*N),w4 => d68_in (6*N-1 downto 5*N),w5 => d68_in (5*N-1 downto 4*N),w6 => d68_in (4*N-1 downto 3*N),w7 => d68_in (3*N-1 downto 2*N),w8 => d68_in (2*N-1 downto N),w9 => d68_in (N-1 downto 0 ),d_out => d68_out ,en_out =>open  ,sof_out=>open   );
CL69 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d69_in (9*N-1 downto 8*N),data2conv2 =>d69_in (8*N-1 downto 7*N),data2conv3 =>d69_in (7*N-1 downto 6*N),data2conv4 =>d69_in (6*N-1 downto 5*N),data2conv5 =>d69_in (5*N-1 downto 4*N),data2conv6 =>d69_in (4*N-1 downto 3*N),data2conv7 =>d69_in (3*N-1 downto 2*N),data2conv8 =>d69_in (2*N-1 downto N),data2conv9 =>d69_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d69_in (9*N-1 downto 8*N),w2 => d69_in (8*N-1 downto 7*N),w3 => d69_in (7*N-1 downto 6*N),w4 => d69_in (6*N-1 downto 5*N),w5 => d69_in (5*N-1 downto 4*N),w6 => d69_in (4*N-1 downto 3*N),w7 => d69_in (3*N-1 downto 2*N),w8 => d69_in (2*N-1 downto N),w9 => d69_in (N-1 downto 0 ),d_out => d69_out ,en_out =>open  ,sof_out=>open   );
CL70 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d70_in (9*N-1 downto 8*N),data2conv2 =>d70_in (8*N-1 downto 7*N),data2conv3 =>d70_in (7*N-1 downto 6*N),data2conv4 =>d70_in (6*N-1 downto 5*N),data2conv5 =>d70_in (5*N-1 downto 4*N),data2conv6 =>d70_in (4*N-1 downto 3*N),data2conv7 =>d70_in (3*N-1 downto 2*N),data2conv8 =>d70_in (2*N-1 downto N),data2conv9 =>d70_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d70_in (9*N-1 downto 8*N),w2 => d70_in (8*N-1 downto 7*N),w3 => d70_in (7*N-1 downto 6*N),w4 => d70_in (6*N-1 downto 5*N),w5 => d70_in (5*N-1 downto 4*N),w6 => d70_in (4*N-1 downto 3*N),w7 => d70_in (3*N-1 downto 2*N),w8 => d70_in (2*N-1 downto N),w9 => d70_in (N-1 downto 0 ),d_out => d70_out ,en_out =>open  ,sof_out=>open   );
CL71 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d71_in (9*N-1 downto 8*N),data2conv2 =>d71_in (8*N-1 downto 7*N),data2conv3 =>d71_in (7*N-1 downto 6*N),data2conv4 =>d71_in (6*N-1 downto 5*N),data2conv5 =>d71_in (5*N-1 downto 4*N),data2conv6 =>d71_in (4*N-1 downto 3*N),data2conv7 =>d71_in (3*N-1 downto 2*N),data2conv8 =>d71_in (2*N-1 downto N),data2conv9 =>d71_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d71_in (9*N-1 downto 8*N),w2 => d71_in (8*N-1 downto 7*N),w3 => d71_in (7*N-1 downto 6*N),w4 => d71_in (6*N-1 downto 5*N),w5 => d71_in (5*N-1 downto 4*N),w6 => d71_in (4*N-1 downto 3*N),w7 => d71_in (3*N-1 downto 2*N),w8 => d71_in (2*N-1 downto N),w9 => d71_in (N-1 downto 0 ),d_out => d71_out ,en_out =>open  ,sof_out=>open   );
CL72 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d72_in (9*N-1 downto 8*N),data2conv2 =>d72_in (8*N-1 downto 7*N),data2conv3 =>d72_in (7*N-1 downto 6*N),data2conv4 =>d72_in (6*N-1 downto 5*N),data2conv5 =>d72_in (5*N-1 downto 4*N),data2conv6 =>d72_in (4*N-1 downto 3*N),data2conv7 =>d72_in (3*N-1 downto 2*N),data2conv8 =>d72_in (2*N-1 downto N),data2conv9 =>d72_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d72_in (9*N-1 downto 8*N),w2 => d72_in (8*N-1 downto 7*N),w3 => d72_in (7*N-1 downto 6*N),w4 => d72_in (6*N-1 downto 5*N),w5 => d72_in (5*N-1 downto 4*N),w6 => d72_in (4*N-1 downto 3*N),w7 => d72_in (3*N-1 downto 2*N),w8 => d72_in (2*N-1 downto N),w9 => d72_in (N-1 downto 0 ),d_out => d72_out ,en_out =>open  ,sof_out=>open   );
CL73 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d73_in (9*N-1 downto 8*N),data2conv2 =>d73_in (8*N-1 downto 7*N),data2conv3 =>d73_in (7*N-1 downto 6*N),data2conv4 =>d73_in (6*N-1 downto 5*N),data2conv5 =>d73_in (5*N-1 downto 4*N),data2conv6 =>d73_in (4*N-1 downto 3*N),data2conv7 =>d73_in (3*N-1 downto 2*N),data2conv8 =>d73_in (2*N-1 downto N),data2conv9 =>d73_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d73_in (9*N-1 downto 8*N),w2 => d73_in (8*N-1 downto 7*N),w3 => d73_in (7*N-1 downto 6*N),w4 => d73_in (6*N-1 downto 5*N),w5 => d73_in (5*N-1 downto 4*N),w6 => d73_in (4*N-1 downto 3*N),w7 => d73_in (3*N-1 downto 2*N),w8 => d73_in (2*N-1 downto N),w9 => d73_in (N-1 downto 0 ),d_out => d73_out ,en_out =>open  ,sof_out=>open   );
CL74 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d74_in (9*N-1 downto 8*N),data2conv2 =>d74_in (8*N-1 downto 7*N),data2conv3 =>d74_in (7*N-1 downto 6*N),data2conv4 =>d74_in (6*N-1 downto 5*N),data2conv5 =>d74_in (5*N-1 downto 4*N),data2conv6 =>d74_in (4*N-1 downto 3*N),data2conv7 =>d74_in (3*N-1 downto 2*N),data2conv8 =>d74_in (2*N-1 downto N),data2conv9 =>d74_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d74_in (9*N-1 downto 8*N),w2 => d74_in (8*N-1 downto 7*N),w3 => d74_in (7*N-1 downto 6*N),w4 => d74_in (6*N-1 downto 5*N),w5 => d74_in (5*N-1 downto 4*N),w6 => d74_in (4*N-1 downto 3*N),w7 => d74_in (3*N-1 downto 2*N),w8 => d74_in (2*N-1 downto N),w9 => d74_in (N-1 downto 0 ),d_out => d74_out ,en_out =>open  ,sof_out=>open   );
CL75 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d75_in (9*N-1 downto 8*N),data2conv2 =>d75_in (8*N-1 downto 7*N),data2conv3 =>d75_in (7*N-1 downto 6*N),data2conv4 =>d75_in (6*N-1 downto 5*N),data2conv5 =>d75_in (5*N-1 downto 4*N),data2conv6 =>d75_in (4*N-1 downto 3*N),data2conv7 =>d75_in (3*N-1 downto 2*N),data2conv8 =>d75_in (2*N-1 downto N),data2conv9 =>d75_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d75_in (9*N-1 downto 8*N),w2 => d75_in (8*N-1 downto 7*N),w3 => d75_in (7*N-1 downto 6*N),w4 => d75_in (6*N-1 downto 5*N),w5 => d75_in (5*N-1 downto 4*N),w6 => d75_in (4*N-1 downto 3*N),w7 => d75_in (3*N-1 downto 2*N),w8 => d75_in (2*N-1 downto N),w9 => d75_in (N-1 downto 0 ),d_out => d75_out ,en_out =>open  ,sof_out=>open   );
CL76 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d76_in (9*N-1 downto 8*N),data2conv2 =>d76_in (8*N-1 downto 7*N),data2conv3 =>d76_in (7*N-1 downto 6*N),data2conv4 =>d76_in (6*N-1 downto 5*N),data2conv5 =>d76_in (5*N-1 downto 4*N),data2conv6 =>d76_in (4*N-1 downto 3*N),data2conv7 =>d76_in (3*N-1 downto 2*N),data2conv8 =>d76_in (2*N-1 downto N),data2conv9 =>d76_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d76_in (9*N-1 downto 8*N),w2 => d76_in (8*N-1 downto 7*N),w3 => d76_in (7*N-1 downto 6*N),w4 => d76_in (6*N-1 downto 5*N),w5 => d76_in (5*N-1 downto 4*N),w6 => d76_in (4*N-1 downto 3*N),w7 => d76_in (3*N-1 downto 2*N),w8 => d76_in (2*N-1 downto N),w9 => d76_in (N-1 downto 0 ),d_out => d76_out ,en_out =>open  ,sof_out=>open   );
CL77 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d77_in (9*N-1 downto 8*N),data2conv2 =>d77_in (8*N-1 downto 7*N),data2conv3 =>d77_in (7*N-1 downto 6*N),data2conv4 =>d77_in (6*N-1 downto 5*N),data2conv5 =>d77_in (5*N-1 downto 4*N),data2conv6 =>d77_in (4*N-1 downto 3*N),data2conv7 =>d77_in (3*N-1 downto 2*N),data2conv8 =>d77_in (2*N-1 downto N),data2conv9 =>d77_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d77_in (9*N-1 downto 8*N),w2 => d77_in (8*N-1 downto 7*N),w3 => d77_in (7*N-1 downto 6*N),w4 => d77_in (6*N-1 downto 5*N),w5 => d77_in (5*N-1 downto 4*N),w6 => d77_in (4*N-1 downto 3*N),w7 => d77_in (3*N-1 downto 2*N),w8 => d77_in (2*N-1 downto N),w9 => d77_in (N-1 downto 0 ),d_out => d77_out ,en_out =>open  ,sof_out=>open   );
CL78 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d78_in (9*N-1 downto 8*N),data2conv2 =>d78_in (8*N-1 downto 7*N),data2conv3 =>d78_in (7*N-1 downto 6*N),data2conv4 =>d78_in (6*N-1 downto 5*N),data2conv5 =>d78_in (5*N-1 downto 4*N),data2conv6 =>d78_in (4*N-1 downto 3*N),data2conv7 =>d78_in (3*N-1 downto 2*N),data2conv8 =>d78_in (2*N-1 downto N),data2conv9 =>d78_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d78_in (9*N-1 downto 8*N),w2 => d78_in (8*N-1 downto 7*N),w3 => d78_in (7*N-1 downto 6*N),w4 => d78_in (6*N-1 downto 5*N),w5 => d78_in (5*N-1 downto 4*N),w6 => d78_in (4*N-1 downto 3*N),w7 => d78_in (3*N-1 downto 2*N),w8 => d78_in (2*N-1 downto N),w9 => d78_in (N-1 downto 0 ),d_out => d78_out ,en_out =>open  ,sof_out=>open   );
CL79 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d79_in (9*N-1 downto 8*N),data2conv2 =>d79_in (8*N-1 downto 7*N),data2conv3 =>d79_in (7*N-1 downto 6*N),data2conv4 =>d79_in (6*N-1 downto 5*N),data2conv5 =>d79_in (5*N-1 downto 4*N),data2conv6 =>d79_in (4*N-1 downto 3*N),data2conv7 =>d79_in (3*N-1 downto 2*N),data2conv8 =>d79_in (2*N-1 downto N),data2conv9 =>d79_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d79_in (9*N-1 downto 8*N),w2 => d79_in (8*N-1 downto 7*N),w3 => d79_in (7*N-1 downto 6*N),w4 => d79_in (6*N-1 downto 5*N),w5 => d79_in (5*N-1 downto 4*N),w6 => d79_in (4*N-1 downto 3*N),w7 => d79_in (3*N-1 downto 2*N),w8 => d79_in (2*N-1 downto N),w9 => d79_in (N-1 downto 0 ),d_out => d79_out ,en_out =>open  ,sof_out=>open   );
CL80 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d80_in (9*N-1 downto 8*N),data2conv2 =>d80_in (8*N-1 downto 7*N),data2conv3 =>d80_in (7*N-1 downto 6*N),data2conv4 =>d80_in (6*N-1 downto 5*N),data2conv5 =>d80_in (5*N-1 downto 4*N),data2conv6 =>d80_in (4*N-1 downto 3*N),data2conv7 =>d80_in (3*N-1 downto 2*N),data2conv8 =>d80_in (2*N-1 downto N),data2conv9 =>d80_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d80_in (9*N-1 downto 8*N),w2 => d80_in (8*N-1 downto 7*N),w3 => d80_in (7*N-1 downto 6*N),w4 => d80_in (6*N-1 downto 5*N),w5 => d80_in (5*N-1 downto 4*N),w6 => d80_in (4*N-1 downto 3*N),w7 => d80_in (3*N-1 downto 2*N),w8 => d80_in (2*N-1 downto N),w9 => d80_in (N-1 downto 0 ),d_out => d80_out ,en_out =>open  ,sof_out=>open   );
CL81 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d81_in (9*N-1 downto 8*N),data2conv2 =>d81_in (8*N-1 downto 7*N),data2conv3 =>d81_in (7*N-1 downto 6*N),data2conv4 =>d81_in (6*N-1 downto 5*N),data2conv5 =>d81_in (5*N-1 downto 4*N),data2conv6 =>d81_in (4*N-1 downto 3*N),data2conv7 =>d81_in (3*N-1 downto 2*N),data2conv8 =>d81_in (2*N-1 downto N),data2conv9 =>d81_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d81_in (9*N-1 downto 8*N),w2 => d81_in (8*N-1 downto 7*N),w3 => d81_in (7*N-1 downto 6*N),w4 => d81_in (6*N-1 downto 5*N),w5 => d81_in (5*N-1 downto 4*N),w6 => d81_in (4*N-1 downto 3*N),w7 => d81_in (3*N-1 downto 2*N),w8 => d81_in (2*N-1 downto N),w9 => d81_in (N-1 downto 0 ),d_out => d81_out ,en_out =>open  ,sof_out=>open   );
CL82 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d82_in (9*N-1 downto 8*N),data2conv2 =>d82_in (8*N-1 downto 7*N),data2conv3 =>d82_in (7*N-1 downto 6*N),data2conv4 =>d82_in (6*N-1 downto 5*N),data2conv5 =>d82_in (5*N-1 downto 4*N),data2conv6 =>d82_in (4*N-1 downto 3*N),data2conv7 =>d82_in (3*N-1 downto 2*N),data2conv8 =>d82_in (2*N-1 downto N),data2conv9 =>d82_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d82_in (9*N-1 downto 8*N),w2 => d82_in (8*N-1 downto 7*N),w3 => d82_in (7*N-1 downto 6*N),w4 => d82_in (6*N-1 downto 5*N),w5 => d82_in (5*N-1 downto 4*N),w6 => d82_in (4*N-1 downto 3*N),w7 => d82_in (3*N-1 downto 2*N),w8 => d82_in (2*N-1 downto N),w9 => d82_in (N-1 downto 0 ),d_out => d82_out ,en_out =>open  ,sof_out=>open   );
CL83 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d83_in (9*N-1 downto 8*N),data2conv2 =>d83_in (8*N-1 downto 7*N),data2conv3 =>d83_in (7*N-1 downto 6*N),data2conv4 =>d83_in (6*N-1 downto 5*N),data2conv5 =>d83_in (5*N-1 downto 4*N),data2conv6 =>d83_in (4*N-1 downto 3*N),data2conv7 =>d83_in (3*N-1 downto 2*N),data2conv8 =>d83_in (2*N-1 downto N),data2conv9 =>d83_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d83_in (9*N-1 downto 8*N),w2 => d83_in (8*N-1 downto 7*N),w3 => d83_in (7*N-1 downto 6*N),w4 => d83_in (6*N-1 downto 5*N),w5 => d83_in (5*N-1 downto 4*N),w6 => d83_in (4*N-1 downto 3*N),w7 => d83_in (3*N-1 downto 2*N),w8 => d83_in (2*N-1 downto N),w9 => d83_in (N-1 downto 0 ),d_out => d83_out ,en_out =>open  ,sof_out=>open   );
CL84 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d84_in (9*N-1 downto 8*N),data2conv2 =>d84_in (8*N-1 downto 7*N),data2conv3 =>d84_in (7*N-1 downto 6*N),data2conv4 =>d84_in (6*N-1 downto 5*N),data2conv5 =>d84_in (5*N-1 downto 4*N),data2conv6 =>d84_in (4*N-1 downto 3*N),data2conv7 =>d84_in (3*N-1 downto 2*N),data2conv8 =>d84_in (2*N-1 downto N),data2conv9 =>d84_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d84_in (9*N-1 downto 8*N),w2 => d84_in (8*N-1 downto 7*N),w3 => d84_in (7*N-1 downto 6*N),w4 => d84_in (6*N-1 downto 5*N),w5 => d84_in (5*N-1 downto 4*N),w6 => d84_in (4*N-1 downto 3*N),w7 => d84_in (3*N-1 downto 2*N),w8 => d84_in (2*N-1 downto N),w9 => d84_in (N-1 downto 0 ),d_out => d84_out ,en_out =>open  ,sof_out=>open   );
CL85 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d85_in (9*N-1 downto 8*N),data2conv2 =>d85_in (8*N-1 downto 7*N),data2conv3 =>d85_in (7*N-1 downto 6*N),data2conv4 =>d85_in (6*N-1 downto 5*N),data2conv5 =>d85_in (5*N-1 downto 4*N),data2conv6 =>d85_in (4*N-1 downto 3*N),data2conv7 =>d85_in (3*N-1 downto 2*N),data2conv8 =>d85_in (2*N-1 downto N),data2conv9 =>d85_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d85_in (9*N-1 downto 8*N),w2 => d85_in (8*N-1 downto 7*N),w3 => d85_in (7*N-1 downto 6*N),w4 => d85_in (6*N-1 downto 5*N),w5 => d85_in (5*N-1 downto 4*N),w6 => d85_in (4*N-1 downto 3*N),w7 => d85_in (3*N-1 downto 2*N),w8 => d85_in (2*N-1 downto N),w9 => d85_in (N-1 downto 0 ),d_out => d85_out ,en_out =>open  ,sof_out=>open   );
CL86 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d86_in (9*N-1 downto 8*N),data2conv2 =>d86_in (8*N-1 downto 7*N),data2conv3 =>d86_in (7*N-1 downto 6*N),data2conv4 =>d86_in (6*N-1 downto 5*N),data2conv5 =>d86_in (5*N-1 downto 4*N),data2conv6 =>d86_in (4*N-1 downto 3*N),data2conv7 =>d86_in (3*N-1 downto 2*N),data2conv8 =>d86_in (2*N-1 downto N),data2conv9 =>d86_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d86_in (9*N-1 downto 8*N),w2 => d86_in (8*N-1 downto 7*N),w3 => d86_in (7*N-1 downto 6*N),w4 => d86_in (6*N-1 downto 5*N),w5 => d86_in (5*N-1 downto 4*N),w6 => d86_in (4*N-1 downto 3*N),w7 => d86_in (3*N-1 downto 2*N),w8 => d86_in (2*N-1 downto N),w9 => d86_in (N-1 downto 0 ),d_out => d86_out ,en_out =>open  ,sof_out=>open   );
CL87 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d87_in (9*N-1 downto 8*N),data2conv2 =>d87_in (8*N-1 downto 7*N),data2conv3 =>d87_in (7*N-1 downto 6*N),data2conv4 =>d87_in (6*N-1 downto 5*N),data2conv5 =>d87_in (5*N-1 downto 4*N),data2conv6 =>d87_in (4*N-1 downto 3*N),data2conv7 =>d87_in (3*N-1 downto 2*N),data2conv8 =>d87_in (2*N-1 downto N),data2conv9 =>d87_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d87_in (9*N-1 downto 8*N),w2 => d87_in (8*N-1 downto 7*N),w3 => d87_in (7*N-1 downto 6*N),w4 => d87_in (6*N-1 downto 5*N),w5 => d87_in (5*N-1 downto 4*N),w6 => d87_in (4*N-1 downto 3*N),w7 => d87_in (3*N-1 downto 2*N),w8 => d87_in (2*N-1 downto N),w9 => d87_in (N-1 downto 0 ),d_out => d87_out ,en_out =>open  ,sof_out=>open   );
CL88 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d88_in (9*N-1 downto 8*N),data2conv2 =>d88_in (8*N-1 downto 7*N),data2conv3 =>d88_in (7*N-1 downto 6*N),data2conv4 =>d88_in (6*N-1 downto 5*N),data2conv5 =>d88_in (5*N-1 downto 4*N),data2conv6 =>d88_in (4*N-1 downto 3*N),data2conv7 =>d88_in (3*N-1 downto 2*N),data2conv8 =>d88_in (2*N-1 downto N),data2conv9 =>d88_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d88_in (9*N-1 downto 8*N),w2 => d88_in (8*N-1 downto 7*N),w3 => d88_in (7*N-1 downto 6*N),w4 => d88_in (6*N-1 downto 5*N),w5 => d88_in (5*N-1 downto 4*N),w6 => d88_in (4*N-1 downto 3*N),w7 => d88_in (3*N-1 downto 2*N),w8 => d88_in (2*N-1 downto N),w9 => d88_in (N-1 downto 0 ),d_out => d88_out ,en_out =>open  ,sof_out=>open   );
CL89 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d89_in (9*N-1 downto 8*N),data2conv2 =>d89_in (8*N-1 downto 7*N),data2conv3 =>d89_in (7*N-1 downto 6*N),data2conv4 =>d89_in (6*N-1 downto 5*N),data2conv5 =>d89_in (5*N-1 downto 4*N),data2conv6 =>d89_in (4*N-1 downto 3*N),data2conv7 =>d89_in (3*N-1 downto 2*N),data2conv8 =>d89_in (2*N-1 downto N),data2conv9 =>d89_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d89_in (9*N-1 downto 8*N),w2 => d89_in (8*N-1 downto 7*N),w3 => d89_in (7*N-1 downto 6*N),w4 => d89_in (6*N-1 downto 5*N),w5 => d89_in (5*N-1 downto 4*N),w6 => d89_in (4*N-1 downto 3*N),w7 => d89_in (3*N-1 downto 2*N),w8 => d89_in (2*N-1 downto N),w9 => d89_in (N-1 downto 0 ),d_out => d89_out ,en_out =>open  ,sof_out=>open   );
CL90 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d90_in (9*N-1 downto 8*N),data2conv2 =>d90_in (8*N-1 downto 7*N),data2conv3 =>d90_in (7*N-1 downto 6*N),data2conv4 =>d90_in (6*N-1 downto 5*N),data2conv5 =>d90_in (5*N-1 downto 4*N),data2conv6 =>d90_in (4*N-1 downto 3*N),data2conv7 =>d90_in (3*N-1 downto 2*N),data2conv8 =>d90_in (2*N-1 downto N),data2conv9 =>d90_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d90_in (9*N-1 downto 8*N),w2 => d90_in (8*N-1 downto 7*N),w3 => d90_in (7*N-1 downto 6*N),w4 => d90_in (6*N-1 downto 5*N),w5 => d90_in (5*N-1 downto 4*N),w6 => d90_in (4*N-1 downto 3*N),w7 => d90_in (3*N-1 downto 2*N),w8 => d90_in (2*N-1 downto N),w9 => d90_in (N-1 downto 0 ),d_out => d90_out ,en_out =>open  ,sof_out=>open   );
CL91 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d91_in (9*N-1 downto 8*N),data2conv2 =>d91_in (8*N-1 downto 7*N),data2conv3 =>d91_in (7*N-1 downto 6*N),data2conv4 =>d91_in (6*N-1 downto 5*N),data2conv5 =>d91_in (5*N-1 downto 4*N),data2conv6 =>d91_in (4*N-1 downto 3*N),data2conv7 =>d91_in (3*N-1 downto 2*N),data2conv8 =>d91_in (2*N-1 downto N),data2conv9 =>d91_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d91_in (9*N-1 downto 8*N),w2 => d91_in (8*N-1 downto 7*N),w3 => d91_in (7*N-1 downto 6*N),w4 => d91_in (6*N-1 downto 5*N),w5 => d91_in (5*N-1 downto 4*N),w6 => d91_in (4*N-1 downto 3*N),w7 => d91_in (3*N-1 downto 2*N),w8 => d91_in (2*N-1 downto N),w9 => d91_in (N-1 downto 0 ),d_out => d91_out ,en_out =>open  ,sof_out=>open   );
CL92 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d92_in (9*N-1 downto 8*N),data2conv2 =>d92_in (8*N-1 downto 7*N),data2conv3 =>d92_in (7*N-1 downto 6*N),data2conv4 =>d92_in (6*N-1 downto 5*N),data2conv5 =>d92_in (5*N-1 downto 4*N),data2conv6 =>d92_in (4*N-1 downto 3*N),data2conv7 =>d92_in (3*N-1 downto 2*N),data2conv8 =>d92_in (2*N-1 downto N),data2conv9 =>d92_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d92_in (9*N-1 downto 8*N),w2 => d92_in (8*N-1 downto 7*N),w3 => d92_in (7*N-1 downto 6*N),w4 => d92_in (6*N-1 downto 5*N),w5 => d92_in (5*N-1 downto 4*N),w6 => d92_in (4*N-1 downto 3*N),w7 => d92_in (3*N-1 downto 2*N),w8 => d92_in (2*N-1 downto N),w9 => d92_in (N-1 downto 0 ),d_out => d92_out ,en_out =>open  ,sof_out=>open   );
CL93 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d93_in (9*N-1 downto 8*N),data2conv2 =>d93_in (8*N-1 downto 7*N),data2conv3 =>d93_in (7*N-1 downto 6*N),data2conv4 =>d93_in (6*N-1 downto 5*N),data2conv5 =>d93_in (5*N-1 downto 4*N),data2conv6 =>d93_in (4*N-1 downto 3*N),data2conv7 =>d93_in (3*N-1 downto 2*N),data2conv8 =>d93_in (2*N-1 downto N),data2conv9 =>d93_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d93_in (9*N-1 downto 8*N),w2 => d93_in (8*N-1 downto 7*N),w3 => d93_in (7*N-1 downto 6*N),w4 => d93_in (6*N-1 downto 5*N),w5 => d93_in (5*N-1 downto 4*N),w6 => d93_in (4*N-1 downto 3*N),w7 => d93_in (3*N-1 downto 2*N),w8 => d93_in (2*N-1 downto N),w9 => d93_in (N-1 downto 0 ),d_out => d93_out ,en_out =>open  ,sof_out=>open   );
CL94 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d94_in (9*N-1 downto 8*N),data2conv2 =>d94_in (8*N-1 downto 7*N),data2conv3 =>d94_in (7*N-1 downto 6*N),data2conv4 =>d94_in (6*N-1 downto 5*N),data2conv5 =>d94_in (5*N-1 downto 4*N),data2conv6 =>d94_in (4*N-1 downto 3*N),data2conv7 =>d94_in (3*N-1 downto 2*N),data2conv8 =>d94_in (2*N-1 downto N),data2conv9 =>d94_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d94_in (9*N-1 downto 8*N),w2 => d94_in (8*N-1 downto 7*N),w3 => d94_in (7*N-1 downto 6*N),w4 => d94_in (6*N-1 downto 5*N),w5 => d94_in (5*N-1 downto 4*N),w6 => d94_in (4*N-1 downto 3*N),w7 => d94_in (3*N-1 downto 2*N),w8 => d94_in (2*N-1 downto N),w9 => d94_in (N-1 downto 0 ),d_out => d94_out ,en_out =>open  ,sof_out=>open   );
CL95 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d95_in (9*N-1 downto 8*N),data2conv2 =>d95_in (8*N-1 downto 7*N),data2conv3 =>d95_in (7*N-1 downto 6*N),data2conv4 =>d95_in (6*N-1 downto 5*N),data2conv5 =>d95_in (5*N-1 downto 4*N),data2conv6 =>d95_in (4*N-1 downto 3*N),data2conv7 =>d95_in (3*N-1 downto 2*N),data2conv8 =>d95_in (2*N-1 downto N),data2conv9 =>d95_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d95_in (9*N-1 downto 8*N),w2 => d95_in (8*N-1 downto 7*N),w3 => d95_in (7*N-1 downto 6*N),w4 => d95_in (6*N-1 downto 5*N),w5 => d95_in (5*N-1 downto 4*N),w6 => d95_in (4*N-1 downto 3*N),w7 => d95_in (3*N-1 downto 2*N),w8 => d95_in (2*N-1 downto N),w9 => d95_in (N-1 downto 0 ),d_out => d95_out ,en_out =>open  ,sof_out=>open   );
CL96 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d96_in (9*N-1 downto 8*N),data2conv2 =>d96_in (8*N-1 downto 7*N),data2conv3 =>d96_in (7*N-1 downto 6*N),data2conv4 =>d96_in (6*N-1 downto 5*N),data2conv5 =>d96_in (5*N-1 downto 4*N),data2conv6 =>d96_in (4*N-1 downto 3*N),data2conv7 =>d96_in (3*N-1 downto 2*N),data2conv8 =>d96_in (2*N-1 downto N),data2conv9 =>d96_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d96_in (9*N-1 downto 8*N),w2 => d96_in (8*N-1 downto 7*N),w3 => d96_in (7*N-1 downto 6*N),w4 => d96_in (6*N-1 downto 5*N),w5 => d96_in (5*N-1 downto 4*N),w6 => d96_in (4*N-1 downto 3*N),w7 => d96_in (3*N-1 downto 2*N),w8 => d96_in (2*N-1 downto N),w9 => d96_in (N-1 downto 0 ),d_out => d96_out ,en_out =>open  ,sof_out=>open   );
CL97 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d97_in (9*N-1 downto 8*N),data2conv2 =>d97_in (8*N-1 downto 7*N),data2conv3 =>d97_in (7*N-1 downto 6*N),data2conv4 =>d97_in (6*N-1 downto 5*N),data2conv5 =>d97_in (5*N-1 downto 4*N),data2conv6 =>d97_in (4*N-1 downto 3*N),data2conv7 =>d97_in (3*N-1 downto 2*N),data2conv8 =>d97_in (2*N-1 downto N),data2conv9 =>d97_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d97_in (9*N-1 downto 8*N),w2 => d97_in (8*N-1 downto 7*N),w3 => d97_in (7*N-1 downto 6*N),w4 => d97_in (6*N-1 downto 5*N),w5 => d97_in (5*N-1 downto 4*N),w6 => d97_in (4*N-1 downto 3*N),w7 => d97_in (3*N-1 downto 2*N),w8 => d97_in (2*N-1 downto N),w9 => d97_in (N-1 downto 0 ),d_out => d97_out ,en_out =>open  ,sof_out=>open   );
CL98 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d98_in (9*N-1 downto 8*N),data2conv2 =>d98_in (8*N-1 downto 7*N),data2conv3 =>d98_in (7*N-1 downto 6*N),data2conv4 =>d98_in (6*N-1 downto 5*N),data2conv5 =>d98_in (5*N-1 downto 4*N),data2conv6 =>d98_in (4*N-1 downto 3*N),data2conv7 =>d98_in (3*N-1 downto 2*N),data2conv8 =>d98_in (2*N-1 downto N),data2conv9 =>d98_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d98_in (9*N-1 downto 8*N),w2 => d98_in (8*N-1 downto 7*N),w3 => d98_in (7*N-1 downto 6*N),w4 => d98_in (6*N-1 downto 5*N),w5 => d98_in (5*N-1 downto 4*N),w6 => d98_in (4*N-1 downto 3*N),w7 => d98_in (3*N-1 downto 2*N),w8 => d98_in (2*N-1 downto N),w9 => d98_in (N-1 downto 0 ),d_out => d98_out ,en_out =>open  ,sof_out=>open   );
CL99 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d99_in (9*N-1 downto 8*N),data2conv2 =>d99_in (8*N-1 downto 7*N),data2conv3 =>d99_in (7*N-1 downto 6*N),data2conv4 =>d99_in (6*N-1 downto 5*N),data2conv5 =>d99_in (5*N-1 downto 4*N),data2conv6 =>d99_in (4*N-1 downto 3*N),data2conv7 =>d99_in (3*N-1 downto 2*N),data2conv8 =>d99_in (2*N-1 downto N),data2conv9 =>d99_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d99_in (9*N-1 downto 8*N),w2 => d99_in (8*N-1 downto 7*N),w3 => d99_in (7*N-1 downto 6*N),w4 => d99_in (6*N-1 downto 5*N),w5 => d99_in (5*N-1 downto 4*N),w6 => d99_in (4*N-1 downto 3*N),w7 => d99_in (3*N-1 downto 2*N),w8 => d99_in (2*N-1 downto N),w9 => d99_in (N-1 downto 0 ),d_out => d99_out ,en_out =>open  ,sof_out=>open   );
CL100: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d100_in(9*N-1 downto 8*N),data2conv2 =>d100_in(8*N-1 downto 7*N),data2conv3 =>d100_in(7*N-1 downto 6*N),data2conv4 =>d100_in(6*N-1 downto 5*N),data2conv5 =>d100_in(5*N-1 downto 4*N),data2conv6 =>d100_in(4*N-1 downto 3*N),data2conv7 =>d100_in(3*N-1 downto 2*N),data2conv8 =>d100_in(2*N-1 downto N),data2conv9 =>d100_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d100_in(9*N-1 downto 8*N),w2 => d100_in(8*N-1 downto 7*N),w3 => d100_in(7*N-1 downto 6*N),w4 => d100_in(6*N-1 downto 5*N),w5 => d100_in(5*N-1 downto 4*N),w6 => d100_in(4*N-1 downto 3*N),w7 => d100_in(3*N-1 downto 2*N),w8 => d100_in(2*N-1 downto N),w9 => d100_in(N-1 downto 0 ),d_out => d100_out,en_out =>open  ,sof_out=>open   );
CL101: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d101_in(9*N-1 downto 8*N),data2conv2 =>d101_in(8*N-1 downto 7*N),data2conv3 =>d101_in(7*N-1 downto 6*N),data2conv4 =>d101_in(6*N-1 downto 5*N),data2conv5 =>d101_in(5*N-1 downto 4*N),data2conv6 =>d101_in(4*N-1 downto 3*N),data2conv7 =>d101_in(3*N-1 downto 2*N),data2conv8 =>d101_in(2*N-1 downto N),data2conv9 =>d101_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d101_in(9*N-1 downto 8*N),w2 => d101_in(8*N-1 downto 7*N),w3 => d101_in(7*N-1 downto 6*N),w4 => d101_in(6*N-1 downto 5*N),w5 => d101_in(5*N-1 downto 4*N),w6 => d101_in(4*N-1 downto 3*N),w7 => d101_in(3*N-1 downto 2*N),w8 => d101_in(2*N-1 downto N),w9 => d101_in(N-1 downto 0 ),d_out => d101_out,en_out =>open  ,sof_out=>open   );
CL102: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d102_in(9*N-1 downto 8*N),data2conv2 =>d102_in(8*N-1 downto 7*N),data2conv3 =>d102_in(7*N-1 downto 6*N),data2conv4 =>d102_in(6*N-1 downto 5*N),data2conv5 =>d102_in(5*N-1 downto 4*N),data2conv6 =>d102_in(4*N-1 downto 3*N),data2conv7 =>d102_in(3*N-1 downto 2*N),data2conv8 =>d102_in(2*N-1 downto N),data2conv9 =>d102_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d102_in(9*N-1 downto 8*N),w2 => d102_in(8*N-1 downto 7*N),w3 => d102_in(7*N-1 downto 6*N),w4 => d102_in(6*N-1 downto 5*N),w5 => d102_in(5*N-1 downto 4*N),w6 => d102_in(4*N-1 downto 3*N),w7 => d102_in(3*N-1 downto 2*N),w8 => d102_in(2*N-1 downto N),w9 => d102_in(N-1 downto 0 ),d_out => d102_out,en_out =>open  ,sof_out=>open   );
CL103: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d103_in(9*N-1 downto 8*N),data2conv2 =>d103_in(8*N-1 downto 7*N),data2conv3 =>d103_in(7*N-1 downto 6*N),data2conv4 =>d103_in(6*N-1 downto 5*N),data2conv5 =>d103_in(5*N-1 downto 4*N),data2conv6 =>d103_in(4*N-1 downto 3*N),data2conv7 =>d103_in(3*N-1 downto 2*N),data2conv8 =>d103_in(2*N-1 downto N),data2conv9 =>d103_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d103_in(9*N-1 downto 8*N),w2 => d103_in(8*N-1 downto 7*N),w3 => d103_in(7*N-1 downto 6*N),w4 => d103_in(6*N-1 downto 5*N),w5 => d103_in(5*N-1 downto 4*N),w6 => d103_in(4*N-1 downto 3*N),w7 => d103_in(3*N-1 downto 2*N),w8 => d103_in(2*N-1 downto N),w9 => d103_in(N-1 downto 0 ),d_out => d103_out,en_out =>open  ,sof_out=>open   );
CL104: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d104_in(9*N-1 downto 8*N),data2conv2 =>d104_in(8*N-1 downto 7*N),data2conv3 =>d104_in(7*N-1 downto 6*N),data2conv4 =>d104_in(6*N-1 downto 5*N),data2conv5 =>d104_in(5*N-1 downto 4*N),data2conv6 =>d104_in(4*N-1 downto 3*N),data2conv7 =>d104_in(3*N-1 downto 2*N),data2conv8 =>d104_in(2*N-1 downto N),data2conv9 =>d104_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d104_in(9*N-1 downto 8*N),w2 => d104_in(8*N-1 downto 7*N),w3 => d104_in(7*N-1 downto 6*N),w4 => d104_in(6*N-1 downto 5*N),w5 => d104_in(5*N-1 downto 4*N),w6 => d104_in(4*N-1 downto 3*N),w7 => d104_in(3*N-1 downto 2*N),w8 => d104_in(2*N-1 downto N),w9 => d104_in(N-1 downto 0 ),d_out => d104_out,en_out =>open  ,sof_out=>open   );
CL105: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d105_in(9*N-1 downto 8*N),data2conv2 =>d105_in(8*N-1 downto 7*N),data2conv3 =>d105_in(7*N-1 downto 6*N),data2conv4 =>d105_in(6*N-1 downto 5*N),data2conv5 =>d105_in(5*N-1 downto 4*N),data2conv6 =>d105_in(4*N-1 downto 3*N),data2conv7 =>d105_in(3*N-1 downto 2*N),data2conv8 =>d105_in(2*N-1 downto N),data2conv9 =>d105_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d105_in(9*N-1 downto 8*N),w2 => d105_in(8*N-1 downto 7*N),w3 => d105_in(7*N-1 downto 6*N),w4 => d105_in(6*N-1 downto 5*N),w5 => d105_in(5*N-1 downto 4*N),w6 => d105_in(4*N-1 downto 3*N),w7 => d105_in(3*N-1 downto 2*N),w8 => d105_in(2*N-1 downto N),w9 => d105_in(N-1 downto 0 ),d_out => d105_out,en_out =>open  ,sof_out=>open   );
CL106: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d106_in(9*N-1 downto 8*N),data2conv2 =>d106_in(8*N-1 downto 7*N),data2conv3 =>d106_in(7*N-1 downto 6*N),data2conv4 =>d106_in(6*N-1 downto 5*N),data2conv5 =>d106_in(5*N-1 downto 4*N),data2conv6 =>d106_in(4*N-1 downto 3*N),data2conv7 =>d106_in(3*N-1 downto 2*N),data2conv8 =>d106_in(2*N-1 downto N),data2conv9 =>d106_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d106_in(9*N-1 downto 8*N),w2 => d106_in(8*N-1 downto 7*N),w3 => d106_in(7*N-1 downto 6*N),w4 => d106_in(6*N-1 downto 5*N),w5 => d106_in(5*N-1 downto 4*N),w6 => d106_in(4*N-1 downto 3*N),w7 => d106_in(3*N-1 downto 2*N),w8 => d106_in(2*N-1 downto N),w9 => d106_in(N-1 downto 0 ),d_out => d106_out,en_out =>open  ,sof_out=>open   );
CL107: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d107_in(9*N-1 downto 8*N),data2conv2 =>d107_in(8*N-1 downto 7*N),data2conv3 =>d107_in(7*N-1 downto 6*N),data2conv4 =>d107_in(6*N-1 downto 5*N),data2conv5 =>d107_in(5*N-1 downto 4*N),data2conv6 =>d107_in(4*N-1 downto 3*N),data2conv7 =>d107_in(3*N-1 downto 2*N),data2conv8 =>d107_in(2*N-1 downto N),data2conv9 =>d107_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d107_in(9*N-1 downto 8*N),w2 => d107_in(8*N-1 downto 7*N),w3 => d107_in(7*N-1 downto 6*N),w4 => d107_in(6*N-1 downto 5*N),w5 => d107_in(5*N-1 downto 4*N),w6 => d107_in(4*N-1 downto 3*N),w7 => d107_in(3*N-1 downto 2*N),w8 => d107_in(2*N-1 downto N),w9 => d107_in(N-1 downto 0 ),d_out => d107_out,en_out =>open  ,sof_out=>open   );
CL108: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d108_in(9*N-1 downto 8*N),data2conv2 =>d108_in(8*N-1 downto 7*N),data2conv3 =>d108_in(7*N-1 downto 6*N),data2conv4 =>d108_in(6*N-1 downto 5*N),data2conv5 =>d108_in(5*N-1 downto 4*N),data2conv6 =>d108_in(4*N-1 downto 3*N),data2conv7 =>d108_in(3*N-1 downto 2*N),data2conv8 =>d108_in(2*N-1 downto N),data2conv9 =>d108_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d108_in(9*N-1 downto 8*N),w2 => d108_in(8*N-1 downto 7*N),w3 => d108_in(7*N-1 downto 6*N),w4 => d108_in(6*N-1 downto 5*N),w5 => d108_in(5*N-1 downto 4*N),w6 => d108_in(4*N-1 downto 3*N),w7 => d108_in(3*N-1 downto 2*N),w8 => d108_in(2*N-1 downto N),w9 => d108_in(N-1 downto 0 ),d_out => d108_out,en_out =>open  ,sof_out=>open   );
CL109: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d109_in(9*N-1 downto 8*N),data2conv2 =>d109_in(8*N-1 downto 7*N),data2conv3 =>d109_in(7*N-1 downto 6*N),data2conv4 =>d109_in(6*N-1 downto 5*N),data2conv5 =>d109_in(5*N-1 downto 4*N),data2conv6 =>d109_in(4*N-1 downto 3*N),data2conv7 =>d109_in(3*N-1 downto 2*N),data2conv8 =>d109_in(2*N-1 downto N),data2conv9 =>d109_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d109_in(9*N-1 downto 8*N),w2 => d109_in(8*N-1 downto 7*N),w3 => d109_in(7*N-1 downto 6*N),w4 => d109_in(6*N-1 downto 5*N),w5 => d109_in(5*N-1 downto 4*N),w6 => d109_in(4*N-1 downto 3*N),w7 => d109_in(3*N-1 downto 2*N),w8 => d109_in(2*N-1 downto N),w9 => d109_in(N-1 downto 0 ),d_out => d109_out,en_out =>open  ,sof_out=>open   );
CL110: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d110_in(9*N-1 downto 8*N),data2conv2 =>d110_in(8*N-1 downto 7*N),data2conv3 =>d110_in(7*N-1 downto 6*N),data2conv4 =>d110_in(6*N-1 downto 5*N),data2conv5 =>d110_in(5*N-1 downto 4*N),data2conv6 =>d110_in(4*N-1 downto 3*N),data2conv7 =>d110_in(3*N-1 downto 2*N),data2conv8 =>d110_in(2*N-1 downto N),data2conv9 =>d110_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d110_in(9*N-1 downto 8*N),w2 => d110_in(8*N-1 downto 7*N),w3 => d110_in(7*N-1 downto 6*N),w4 => d110_in(6*N-1 downto 5*N),w5 => d110_in(5*N-1 downto 4*N),w6 => d110_in(4*N-1 downto 3*N),w7 => d110_in(3*N-1 downto 2*N),w8 => d110_in(2*N-1 downto N),w9 => d110_in(N-1 downto 0 ),d_out => d110_out,en_out =>open  ,sof_out=>open   );
CL111: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d111_in(9*N-1 downto 8*N),data2conv2 =>d111_in(8*N-1 downto 7*N),data2conv3 =>d111_in(7*N-1 downto 6*N),data2conv4 =>d111_in(6*N-1 downto 5*N),data2conv5 =>d111_in(5*N-1 downto 4*N),data2conv6 =>d111_in(4*N-1 downto 3*N),data2conv7 =>d111_in(3*N-1 downto 2*N),data2conv8 =>d111_in(2*N-1 downto N),data2conv9 =>d111_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d111_in(9*N-1 downto 8*N),w2 => d111_in(8*N-1 downto 7*N),w3 => d111_in(7*N-1 downto 6*N),w4 => d111_in(6*N-1 downto 5*N),w5 => d111_in(5*N-1 downto 4*N),w6 => d111_in(4*N-1 downto 3*N),w7 => d111_in(3*N-1 downto 2*N),w8 => d111_in(2*N-1 downto N),w9 => d111_in(N-1 downto 0 ),d_out => d111_out,en_out =>open  ,sof_out=>open   );
CL112: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d112_in(9*N-1 downto 8*N),data2conv2 =>d112_in(8*N-1 downto 7*N),data2conv3 =>d112_in(7*N-1 downto 6*N),data2conv4 =>d112_in(6*N-1 downto 5*N),data2conv5 =>d112_in(5*N-1 downto 4*N),data2conv6 =>d112_in(4*N-1 downto 3*N),data2conv7 =>d112_in(3*N-1 downto 2*N),data2conv8 =>d112_in(2*N-1 downto N),data2conv9 =>d112_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d112_in(9*N-1 downto 8*N),w2 => d112_in(8*N-1 downto 7*N),w3 => d112_in(7*N-1 downto 6*N),w4 => d112_in(6*N-1 downto 5*N),w5 => d112_in(5*N-1 downto 4*N),w6 => d112_in(4*N-1 downto 3*N),w7 => d112_in(3*N-1 downto 2*N),w8 => d112_in(2*N-1 downto N),w9 => d112_in(N-1 downto 0 ),d_out => d112_out,en_out =>open  ,sof_out=>open   );
CL113: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d113_in(9*N-1 downto 8*N),data2conv2 =>d113_in(8*N-1 downto 7*N),data2conv3 =>d113_in(7*N-1 downto 6*N),data2conv4 =>d113_in(6*N-1 downto 5*N),data2conv5 =>d113_in(5*N-1 downto 4*N),data2conv6 =>d113_in(4*N-1 downto 3*N),data2conv7 =>d113_in(3*N-1 downto 2*N),data2conv8 =>d113_in(2*N-1 downto N),data2conv9 =>d113_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d113_in(9*N-1 downto 8*N),w2 => d113_in(8*N-1 downto 7*N),w3 => d113_in(7*N-1 downto 6*N),w4 => d113_in(6*N-1 downto 5*N),w5 => d113_in(5*N-1 downto 4*N),w6 => d113_in(4*N-1 downto 3*N),w7 => d113_in(3*N-1 downto 2*N),w8 => d113_in(2*N-1 downto N),w9 => d113_in(N-1 downto 0 ),d_out => d113_out,en_out =>open  ,sof_out=>open   );
CL114: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d114_in(9*N-1 downto 8*N),data2conv2 =>d114_in(8*N-1 downto 7*N),data2conv3 =>d114_in(7*N-1 downto 6*N),data2conv4 =>d114_in(6*N-1 downto 5*N),data2conv5 =>d114_in(5*N-1 downto 4*N),data2conv6 =>d114_in(4*N-1 downto 3*N),data2conv7 =>d114_in(3*N-1 downto 2*N),data2conv8 =>d114_in(2*N-1 downto N),data2conv9 =>d114_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d114_in(9*N-1 downto 8*N),w2 => d114_in(8*N-1 downto 7*N),w3 => d114_in(7*N-1 downto 6*N),w4 => d114_in(6*N-1 downto 5*N),w5 => d114_in(5*N-1 downto 4*N),w6 => d114_in(4*N-1 downto 3*N),w7 => d114_in(3*N-1 downto 2*N),w8 => d114_in(2*N-1 downto N),w9 => d114_in(N-1 downto 0 ),d_out => d114_out,en_out =>open  ,sof_out=>open   );
CL115: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d115_in(9*N-1 downto 8*N),data2conv2 =>d115_in(8*N-1 downto 7*N),data2conv3 =>d115_in(7*N-1 downto 6*N),data2conv4 =>d115_in(6*N-1 downto 5*N),data2conv5 =>d115_in(5*N-1 downto 4*N),data2conv6 =>d115_in(4*N-1 downto 3*N),data2conv7 =>d115_in(3*N-1 downto 2*N),data2conv8 =>d115_in(2*N-1 downto N),data2conv9 =>d115_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d115_in(9*N-1 downto 8*N),w2 => d115_in(8*N-1 downto 7*N),w3 => d115_in(7*N-1 downto 6*N),w4 => d115_in(6*N-1 downto 5*N),w5 => d115_in(5*N-1 downto 4*N),w6 => d115_in(4*N-1 downto 3*N),w7 => d115_in(3*N-1 downto 2*N),w8 => d115_in(2*N-1 downto N),w9 => d115_in(N-1 downto 0 ),d_out => d115_out,en_out =>open  ,sof_out=>open   );
CL116: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d116_in(9*N-1 downto 8*N),data2conv2 =>d116_in(8*N-1 downto 7*N),data2conv3 =>d116_in(7*N-1 downto 6*N),data2conv4 =>d116_in(6*N-1 downto 5*N),data2conv5 =>d116_in(5*N-1 downto 4*N),data2conv6 =>d116_in(4*N-1 downto 3*N),data2conv7 =>d116_in(3*N-1 downto 2*N),data2conv8 =>d116_in(2*N-1 downto N),data2conv9 =>d116_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d116_in(9*N-1 downto 8*N),w2 => d116_in(8*N-1 downto 7*N),w3 => d116_in(7*N-1 downto 6*N),w4 => d116_in(6*N-1 downto 5*N),w5 => d116_in(5*N-1 downto 4*N),w6 => d116_in(4*N-1 downto 3*N),w7 => d116_in(3*N-1 downto 2*N),w8 => d116_in(2*N-1 downto N),w9 => d116_in(N-1 downto 0 ),d_out => d116_out,en_out =>open  ,sof_out=>open   );
CL117: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d117_in(9*N-1 downto 8*N),data2conv2 =>d117_in(8*N-1 downto 7*N),data2conv3 =>d117_in(7*N-1 downto 6*N),data2conv4 =>d117_in(6*N-1 downto 5*N),data2conv5 =>d117_in(5*N-1 downto 4*N),data2conv6 =>d117_in(4*N-1 downto 3*N),data2conv7 =>d117_in(3*N-1 downto 2*N),data2conv8 =>d117_in(2*N-1 downto N),data2conv9 =>d117_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d117_in(9*N-1 downto 8*N),w2 => d117_in(8*N-1 downto 7*N),w3 => d117_in(7*N-1 downto 6*N),w4 => d117_in(6*N-1 downto 5*N),w5 => d117_in(5*N-1 downto 4*N),w6 => d117_in(4*N-1 downto 3*N),w7 => d117_in(3*N-1 downto 2*N),w8 => d117_in(2*N-1 downto N),w9 => d117_in(N-1 downto 0 ),d_out => d117_out,en_out =>open  ,sof_out=>open   );
CL118: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d118_in(9*N-1 downto 8*N),data2conv2 =>d118_in(8*N-1 downto 7*N),data2conv3 =>d118_in(7*N-1 downto 6*N),data2conv4 =>d118_in(6*N-1 downto 5*N),data2conv5 =>d118_in(5*N-1 downto 4*N),data2conv6 =>d118_in(4*N-1 downto 3*N),data2conv7 =>d118_in(3*N-1 downto 2*N),data2conv8 =>d118_in(2*N-1 downto N),data2conv9 =>d118_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d118_in(9*N-1 downto 8*N),w2 => d118_in(8*N-1 downto 7*N),w3 => d118_in(7*N-1 downto 6*N),w4 => d118_in(6*N-1 downto 5*N),w5 => d118_in(5*N-1 downto 4*N),w6 => d118_in(4*N-1 downto 3*N),w7 => d118_in(3*N-1 downto 2*N),w8 => d118_in(2*N-1 downto N),w9 => d118_in(N-1 downto 0 ),d_out => d118_out,en_out =>open  ,sof_out=>open   );
CL119: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d119_in(9*N-1 downto 8*N),data2conv2 =>d119_in(8*N-1 downto 7*N),data2conv3 =>d119_in(7*N-1 downto 6*N),data2conv4 =>d119_in(6*N-1 downto 5*N),data2conv5 =>d119_in(5*N-1 downto 4*N),data2conv6 =>d119_in(4*N-1 downto 3*N),data2conv7 =>d119_in(3*N-1 downto 2*N),data2conv8 =>d119_in(2*N-1 downto N),data2conv9 =>d119_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d119_in(9*N-1 downto 8*N),w2 => d119_in(8*N-1 downto 7*N),w3 => d119_in(7*N-1 downto 6*N),w4 => d119_in(6*N-1 downto 5*N),w5 => d119_in(5*N-1 downto 4*N),w6 => d119_in(4*N-1 downto 3*N),w7 => d119_in(3*N-1 downto 2*N),w8 => d119_in(2*N-1 downto N),w9 => d119_in(N-1 downto 0 ),d_out => d119_out,en_out =>open  ,sof_out=>open   );
CL120: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d120_in(9*N-1 downto 8*N),data2conv2 =>d120_in(8*N-1 downto 7*N),data2conv3 =>d120_in(7*N-1 downto 6*N),data2conv4 =>d120_in(6*N-1 downto 5*N),data2conv5 =>d120_in(5*N-1 downto 4*N),data2conv6 =>d120_in(4*N-1 downto 3*N),data2conv7 =>d120_in(3*N-1 downto 2*N),data2conv8 =>d120_in(2*N-1 downto N),data2conv9 =>d120_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d120_in(9*N-1 downto 8*N),w2 => d120_in(8*N-1 downto 7*N),w3 => d120_in(7*N-1 downto 6*N),w4 => d120_in(6*N-1 downto 5*N),w5 => d120_in(5*N-1 downto 4*N),w6 => d120_in(4*N-1 downto 3*N),w7 => d120_in(3*N-1 downto 2*N),w8 => d120_in(2*N-1 downto N),w9 => d120_in(N-1 downto 0 ),d_out => d120_out,en_out =>open  ,sof_out=>open   );
CL121: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d121_in(9*N-1 downto 8*N),data2conv2 =>d121_in(8*N-1 downto 7*N),data2conv3 =>d121_in(7*N-1 downto 6*N),data2conv4 =>d121_in(6*N-1 downto 5*N),data2conv5 =>d121_in(5*N-1 downto 4*N),data2conv6 =>d121_in(4*N-1 downto 3*N),data2conv7 =>d121_in(3*N-1 downto 2*N),data2conv8 =>d121_in(2*N-1 downto N),data2conv9 =>d121_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d121_in(9*N-1 downto 8*N),w2 => d121_in(8*N-1 downto 7*N),w3 => d121_in(7*N-1 downto 6*N),w4 => d121_in(6*N-1 downto 5*N),w5 => d121_in(5*N-1 downto 4*N),w6 => d121_in(4*N-1 downto 3*N),w7 => d121_in(3*N-1 downto 2*N),w8 => d121_in(2*N-1 downto N),w9 => d121_in(N-1 downto 0 ),d_out => d121_out,en_out =>open  ,sof_out=>open   );
CL122: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d122_in(9*N-1 downto 8*N),data2conv2 =>d122_in(8*N-1 downto 7*N),data2conv3 =>d122_in(7*N-1 downto 6*N),data2conv4 =>d122_in(6*N-1 downto 5*N),data2conv5 =>d122_in(5*N-1 downto 4*N),data2conv6 =>d122_in(4*N-1 downto 3*N),data2conv7 =>d122_in(3*N-1 downto 2*N),data2conv8 =>d122_in(2*N-1 downto N),data2conv9 =>d122_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d122_in(9*N-1 downto 8*N),w2 => d122_in(8*N-1 downto 7*N),w3 => d122_in(7*N-1 downto 6*N),w4 => d122_in(6*N-1 downto 5*N),w5 => d122_in(5*N-1 downto 4*N),w6 => d122_in(4*N-1 downto 3*N),w7 => d122_in(3*N-1 downto 2*N),w8 => d122_in(2*N-1 downto N),w9 => d122_in(N-1 downto 0 ),d_out => d122_out,en_out =>open  ,sof_out=>open   );
CL123: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d123_in(9*N-1 downto 8*N),data2conv2 =>d123_in(8*N-1 downto 7*N),data2conv3 =>d123_in(7*N-1 downto 6*N),data2conv4 =>d123_in(6*N-1 downto 5*N),data2conv5 =>d123_in(5*N-1 downto 4*N),data2conv6 =>d123_in(4*N-1 downto 3*N),data2conv7 =>d123_in(3*N-1 downto 2*N),data2conv8 =>d123_in(2*N-1 downto N),data2conv9 =>d123_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d123_in(9*N-1 downto 8*N),w2 => d123_in(8*N-1 downto 7*N),w3 => d123_in(7*N-1 downto 6*N),w4 => d123_in(6*N-1 downto 5*N),w5 => d123_in(5*N-1 downto 4*N),w6 => d123_in(4*N-1 downto 3*N),w7 => d123_in(3*N-1 downto 2*N),w8 => d123_in(2*N-1 downto N),w9 => d123_in(N-1 downto 0 ),d_out => d123_out,en_out =>open  ,sof_out=>open   );
CL124: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d124_in(9*N-1 downto 8*N),data2conv2 =>d124_in(8*N-1 downto 7*N),data2conv3 =>d124_in(7*N-1 downto 6*N),data2conv4 =>d124_in(6*N-1 downto 5*N),data2conv5 =>d124_in(5*N-1 downto 4*N),data2conv6 =>d124_in(4*N-1 downto 3*N),data2conv7 =>d124_in(3*N-1 downto 2*N),data2conv8 =>d124_in(2*N-1 downto N),data2conv9 =>d124_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d124_in(9*N-1 downto 8*N),w2 => d124_in(8*N-1 downto 7*N),w3 => d124_in(7*N-1 downto 6*N),w4 => d124_in(6*N-1 downto 5*N),w5 => d124_in(5*N-1 downto 4*N),w6 => d124_in(4*N-1 downto 3*N),w7 => d124_in(3*N-1 downto 2*N),w8 => d124_in(2*N-1 downto N),w9 => d124_in(N-1 downto 0 ),d_out => d124_out,en_out =>open  ,sof_out=>open   );
CL125: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d125_in(9*N-1 downto 8*N),data2conv2 =>d125_in(8*N-1 downto 7*N),data2conv3 =>d125_in(7*N-1 downto 6*N),data2conv4 =>d125_in(6*N-1 downto 5*N),data2conv5 =>d125_in(5*N-1 downto 4*N),data2conv6 =>d125_in(4*N-1 downto 3*N),data2conv7 =>d125_in(3*N-1 downto 2*N),data2conv8 =>d125_in(2*N-1 downto N),data2conv9 =>d125_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d125_in(9*N-1 downto 8*N),w2 => d125_in(8*N-1 downto 7*N),w3 => d125_in(7*N-1 downto 6*N),w4 => d125_in(6*N-1 downto 5*N),w5 => d125_in(5*N-1 downto 4*N),w6 => d125_in(4*N-1 downto 3*N),w7 => d125_in(3*N-1 downto 2*N),w8 => d125_in(2*N-1 downto N),w9 => d125_in(N-1 downto 0 ),d_out => d125_out,en_out =>open  ,sof_out=>open   );
CL126: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d126_in(9*N-1 downto 8*N),data2conv2 =>d126_in(8*N-1 downto 7*N),data2conv3 =>d126_in(7*N-1 downto 6*N),data2conv4 =>d126_in(6*N-1 downto 5*N),data2conv5 =>d126_in(5*N-1 downto 4*N),data2conv6 =>d126_in(4*N-1 downto 3*N),data2conv7 =>d126_in(3*N-1 downto 2*N),data2conv8 =>d126_in(2*N-1 downto N),data2conv9 =>d126_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d126_in(9*N-1 downto 8*N),w2 => d126_in(8*N-1 downto 7*N),w3 => d126_in(7*N-1 downto 6*N),w4 => d126_in(6*N-1 downto 5*N),w5 => d126_in(5*N-1 downto 4*N),w6 => d126_in(4*N-1 downto 3*N),w7 => d126_in(3*N-1 downto 2*N),w8 => d126_in(2*N-1 downto N),w9 => d126_in(N-1 downto 0 ),d_out => d126_out,en_out =>open  ,sof_out=>open   );
CL127: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d127_in(9*N-1 downto 8*N),data2conv2 =>d127_in(8*N-1 downto 7*N),data2conv3 =>d127_in(7*N-1 downto 6*N),data2conv4 =>d127_in(6*N-1 downto 5*N),data2conv5 =>d127_in(5*N-1 downto 4*N),data2conv6 =>d127_in(4*N-1 downto 3*N),data2conv7 =>d127_in(3*N-1 downto 2*N),data2conv8 =>d127_in(2*N-1 downto N),data2conv9 =>d127_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d127_in(9*N-1 downto 8*N),w2 => d127_in(8*N-1 downto 7*N),w3 => d127_in(7*N-1 downto 6*N),w4 => d127_in(6*N-1 downto 5*N),w5 => d127_in(5*N-1 downto 4*N),w6 => d127_in(4*N-1 downto 3*N),w7 => d127_in(3*N-1 downto 2*N),w8 => d127_in(2*N-1 downto N),w9 => d127_in(N-1 downto 0 ),d_out => d127_out,en_out =>open  ,sof_out=>open   );
CL128: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d128_in(9*N-1 downto 8*N),data2conv2 =>d128_in(8*N-1 downto 7*N),data2conv3 =>d128_in(7*N-1 downto 6*N),data2conv4 =>d128_in(6*N-1 downto 5*N),data2conv5 =>d128_in(5*N-1 downto 4*N),data2conv6 =>d128_in(4*N-1 downto 3*N),data2conv7 =>d128_in(3*N-1 downto 2*N),data2conv8 =>d128_in(2*N-1 downto N),data2conv9 =>d128_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d128_in(9*N-1 downto 8*N),w2 => d128_in(8*N-1 downto 7*N),w3 => d128_in(7*N-1 downto 6*N),w4 => d128_in(6*N-1 downto 5*N),w5 => d128_in(5*N-1 downto 4*N),w6 => d128_in(4*N-1 downto 3*N),w7 => d128_in(3*N-1 downto 2*N),w8 => d128_in(2*N-1 downto N),w9 => d128_in(N-1 downto 0 ),d_out => d128_out,en_out =>open  ,sof_out=>open   );

  p_sums: process (clk)
  begin
    if rising_edge(clk) then
       sum1  <= (d01_out(d01_out'left) & d01_out(d01_out'left) & d01_out) +  (d02_out(d02_out'left) & d02_out(d02_out'left) & d02_out) + (d03_out(d03_out'left) & d03_out(d03_out'left) & d03_out) +  (d03_out(d03_out'left) & d03_out(d03_out'left) & d03_out);  
       sum2  <= (d05_out(d05_out'left) & d05_out(d05_out'left) & d05_out) +  (d06_out(d06_out'left) & d06_out(d06_out'left) & d06_out) + (d07_out(d07_out'left) & d07_out(d07_out'left) & d07_out) +  (d07_out(d07_out'left) & d07_out(d07_out'left) & d07_out);  
       sum3  <= (d09_out(d09_out'left) & d09_out(d09_out'left) & d09_out) +  (d10_out(d10_out'left) & d10_out(d10_out'left) & d10_out) + (d11_out(d11_out'left) & d11_out(d11_out'left) & d11_out) +  (d11_out(d11_out'left) & d11_out(d11_out'left) & d11_out);  
       sum4  <= (d13_out(d13_out'left) & d13_out(d13_out'left) & d13_out) +  (d14_out(d14_out'left) & d14_out(d14_out'left) & d14_out) + (d15_out(d15_out'left) & d15_out(d15_out'left) & d15_out) +  (d15_out(d15_out'left) & d15_out(d15_out'left) & d15_out);  
       sum5  <= (d17_out(d17_out'left) & d17_out(d17_out'left) & d17_out) +  (d18_out(d18_out'left) & d18_out(d18_out'left) & d18_out) + (d19_out(d19_out'left) & d19_out(d19_out'left) & d19_out) +  (d19_out(d19_out'left) & d19_out(d19_out'left) & d19_out);  
       sum6  <= (d21_out(d21_out'left) & d21_out(d21_out'left) & d21_out) +  (d22_out(d22_out'left) & d22_out(d22_out'left) & d22_out) + (d23_out(d23_out'left) & d23_out(d23_out'left) & d23_out) +  (d23_out(d23_out'left) & d23_out(d23_out'left) & d23_out);  
       sum7  <= (d25_out(d25_out'left) & d25_out(d25_out'left) & d25_out) +  (d26_out(d26_out'left) & d26_out(d26_out'left) & d26_out) + (d27_out(d27_out'left) & d27_out(d27_out'left) & d27_out) +  (d27_out(d27_out'left) & d27_out(d27_out'left) & d27_out);  
       sum8  <= (d29_out(d29_out'left) & d29_out(d29_out'left) & d29_out) +  (d30_out(d30_out'left) & d30_out(d30_out'left) & d30_out) + (d31_out(d31_out'left) & d31_out(d31_out'left) & d31_out) +  (d31_out(d31_out'left) & d31_out(d31_out'left) & d31_out);  
       sum9  <= (d33_out(d33_out'left) & d33_out(d33_out'left) & d33_out) +  (d34_out(d34_out'left) & d34_out(d34_out'left) & d34_out) + (d35_out(d35_out'left) & d35_out(d35_out'left) & d35_out) +  (d35_out(d35_out'left) & d35_out(d35_out'left) & d35_out);  
       sum10 <= (d37_out(d37_out'left) & d37_out(d37_out'left) & d37_out) +  (d38_out(d38_out'left) & d38_out(d38_out'left) & d38_out) + (d39_out(d39_out'left) & d39_out(d39_out'left) & d39_out) +  (d39_out(d39_out'left) & d39_out(d39_out'left) & d39_out);  
       sum11 <= (d41_out(d41_out'left) & d41_out(d41_out'left) & d41_out) +  (d42_out(d42_out'left) & d42_out(d42_out'left) & d42_out) + (d43_out(d43_out'left) & d43_out(d43_out'left) & d43_out) +  (d43_out(d43_out'left) & d43_out(d43_out'left) & d43_out);  
       sum12 <= (d45_out(d45_out'left) & d45_out(d45_out'left) & d45_out) +  (d46_out(d46_out'left) & d46_out(d46_out'left) & d46_out) + (d47_out(d47_out'left) & d47_out(d47_out'left) & d47_out) +  (d47_out(d47_out'left) & d47_out(d47_out'left) & d47_out);  
       sum13 <= (d49_out(d49_out'left) & d49_out(d49_out'left) & d49_out) +  (d50_out(d50_out'left) & d50_out(d50_out'left) & d50_out) + (d51_out(d51_out'left) & d51_out(d51_out'left) & d51_out) +  (d51_out(d51_out'left) & d51_out(d51_out'left) & d51_out);  
       sum14 <= (d53_out(d53_out'left) & d53_out(d53_out'left) & d53_out) +  (d54_out(d54_out'left) & d54_out(d54_out'left) & d54_out) + (d55_out(d55_out'left) & d55_out(d55_out'left) & d55_out) +  (d55_out(d55_out'left) & d55_out(d55_out'left) & d55_out);  
       sum15 <= (d57_out(d57_out'left) & d57_out(d57_out'left) & d57_out) +  (d58_out(d58_out'left) & d58_out(d58_out'left) & d58_out) + (d59_out(d59_out'left) & d59_out(d59_out'left) & d59_out) +  (d59_out(d59_out'left) & d59_out(d59_out'left) & d59_out);  
       sum16 <= (d61_out(d61_out'left) & d61_out(d61_out'left) & d61_out) +  (d62_out(d62_out'left) & d62_out(d62_out'left) & d62_out) + (d63_out(d63_out'left) & d63_out(d63_out'left) & d63_out) +  (d63_out(d63_out'left) & d63_out(d63_out'left) & d63_out);  
       sum22 <= (d65_out (d65_out 'left) & d65_out (d65_out 'left) & d65_out ) + (d66_out (d66_out 'left) & d66_out (d66_out 'left) & d66_out ) + (d67_out (d67_out 'left) & d67_out (d67_out 'left) & d67_out ) + (d68_out (d68_out 'left) & d68_out (d68_out 'left) & d68_out );
       sum23 <= (d69_out (d69_out 'left) & d69_out (d69_out 'left) & d69_out ) + (d70_out (d70_out 'left) & d70_out (d70_out 'left) & d70_out ) + (d71_out (d71_out 'left) & d71_out (d71_out 'left) & d71_out ) + (d72_out (d72_out 'left) & d72_out (d72_out 'left) & d72_out );
       sum24 <= (d73_out (d73_out 'left) & d73_out (d73_out 'left) & d73_out ) + (d74_out (d74_out 'left) & d74_out (d74_out 'left) & d74_out ) + (d75_out (d75_out 'left) & d75_out (d75_out 'left) & d75_out ) + (d76_out (d76_out 'left) & d76_out (d76_out 'left) & d76_out );
       sum25 <= (d77_out (d77_out 'left) & d77_out (d77_out 'left) & d77_out ) + (d78_out (d78_out 'left) & d78_out (d78_out 'left) & d78_out ) + (d79_out (d79_out 'left) & d79_out (d79_out 'left) & d79_out ) + (d80_out (d80_out 'left) & d80_out (d80_out 'left) & d80_out );
       sum26 <= (d81_out (d81_out 'left) & d81_out (d81_out 'left) & d81_out ) + (d82_out (d82_out 'left) & d82_out (d82_out 'left) & d82_out ) + (d83_out (d83_out 'left) & d83_out (d83_out 'left) & d83_out ) + (d84_out (d84_out 'left) & d84_out (d84_out 'left) & d84_out );
       sum27 <= (d85_out (d85_out 'left) & d85_out (d85_out 'left) & d85_out ) + (d86_out (d86_out 'left) & d86_out (d86_out 'left) & d86_out ) + (d87_out (d87_out 'left) & d87_out (d87_out 'left) & d87_out ) + (d88_out (d88_out 'left) & d88_out (d88_out 'left) & d88_out );
       sum28 <= (d89_out (d89_out 'left) & d89_out (d89_out 'left) & d89_out ) + (d90_out (d90_out 'left) & d90_out (d90_out 'left) & d90_out ) + (d91_out (d91_out 'left) & d91_out (d91_out 'left) & d91_out ) + (d92_out (d92_out 'left) & d92_out (d92_out 'left) & d92_out );
       sum29 <= (d93_out (d93_out 'left) & d93_out (d93_out 'left) & d93_out ) + (d94_out (d94_out 'left) & d94_out (d94_out 'left) & d94_out ) + (d95_out (d95_out 'left) & d95_out (d95_out 'left) & d95_out ) + (d96_out (d96_out 'left) & d96_out (d96_out 'left) & d96_out );
       sum30 <= (d97_out (d97_out 'left) & d97_out (d97_out 'left) & d97_out ) + (d98_out (d98_out 'left) & d98_out (d98_out 'left) & d98_out ) + (d99_out (d99_out 'left) & d99_out (d99_out 'left) & d99_out ) + (d100_out(d100_out'left) & d100_out(d100_out'left) & d100_out);
       sum31 <= (d101_out(d101_out'left) & d101_out(d101_out'left) & d101_out) + (d102_out(d102_out'left) & d102_out(d102_out'left) & d102_out) + (d103_out(d103_out'left) & d103_out(d103_out'left) & d103_out) + (d104_out(d104_out'left) & d104_out(d104_out'left) & d104_out);
       sum32 <= (d105_out(d105_out'left) & d105_out(d105_out'left) & d105_out) + (d106_out(d106_out'left) & d106_out(d106_out'left) & d106_out) + (d107_out(d107_out'left) & d107_out(d107_out'left) & d107_out) + (d108_out(d108_out'left) & d108_out(d108_out'left) & d108_out);
       sum33 <= (d109_out(d109_out'left) & d109_out(d109_out'left) & d109_out) + (d110_out(d110_out'left) & d110_out(d110_out'left) & d110_out) + (d111_out(d111_out'left) & d111_out(d111_out'left) & d111_out) + (d112_out(d112_out'left) & d112_out(d112_out'left) & d112_out);
       sum34 <= (d113_out(d113_out'left) & d113_out(d113_out'left) & d113_out) + (d114_out(d114_out'left) & d114_out(d114_out'left) & d114_out) + (d115_out(d115_out'left) & d115_out(d115_out'left) & d115_out) + (d116_out(d116_out'left) & d116_out(d116_out'left) & d116_out);
       sum35 <= (d117_out(d117_out'left) & d117_out(d117_out'left) & d117_out) + (d118_out(d118_out'left) & d118_out(d118_out'left) & d118_out) + (d119_out(d119_out'left) & d119_out(d119_out'left) & d119_out) + (d120_out(d120_out'left) & d120_out(d120_out'left) & d120_out);
       sum36 <= (d121_out(d121_out'left) & d121_out(d121_out'left) & d121_out) + (d122_out(d122_out'left) & d122_out(d122_out'left) & d122_out) + (d123_out(d123_out'left) & d123_out(d123_out'left) & d123_out) + (d124_out(d124_out'left) & d124_out(d124_out'left) & d124_out);
       sum37 <= (d125_out(d125_out'left) & d125_out(d125_out'left) & d125_out) + (d126_out(d126_out'left) & d126_out(d126_out'left) & d126_out) + (d127_out(d127_out'left) & d127_out(d127_out'left) & d127_out) + (d128_out(d128_out'left) & d128_out(d128_out'left) & d128_out);


       sum17 <= (sum1(sum1  'left) & sum1(sum1  'left) & sum1 ) + (sum2(sum2  'left) & sum2(sum2  'left) & sum2 ) + (sum3(sum3  'left) & sum3(sum3  'left) & sum3 ) + (sum4(sum4  'left) & sum4(sum4  'left) & sum4 );  
       sum18 <= (sum5(sum5  'left) & sum5(sum5  'left) & sum5 ) + (sum6(sum6  'left) & sum6(sum6  'left) & sum6 ) + (sum7(sum7  'left) & sum7(sum7  'left) & sum7 ) + (sum8(sum8  'left) & sum8(sum8  'left) & sum8 );  
       sum19 <= (sum9(sum9  'left) & sum9(sum9  'left) & sum9 ) + (sum10(sum10'left) & sum10(sum10'left) & sum10) + (sum11(sum11'left) & sum11(sum11'left) & sum11) + (sum12(sum12'left) & sum12(sum12'left) & sum12);
       sum20 <= (sum13(sum13'left) & sum13(sum13'left) & sum13) + (sum14(sum14'left) & sum14(sum14'left) & sum14) + (sum15(sum15'left) & sum15(sum15'left) & sum15) + (sum16(sum16'left) & sum16(sum16'left) & sum16);
       sum38 <= (sum22(sum22'left) & sum22(sum22'left) & sum22) + (sum23(sum23'left) & sum23(sum23'left) & sum23) + (sum24(sum24'left) & sum24(sum24'left) & sum24) + (sum25(sum25'left) & sum25(sum25'left) & sum25);
       sum39 <= (sum26(sum26'left) & sum26(sum26'left) & sum26) + (sum27(sum27'left) & sum27(sum27'left) & sum27) + (sum28(sum28'left) & sum28(sum28'left) & sum28) + (sum29(sum29'left) & sum29(sum29'left) & sum29);
       sum40 <= (sum30(sum30'left) & sum30(sum30'left) & sum30) + (sum31(sum31'left) & sum31(sum31'left) & sum31) + (sum32(sum32'left) & sum32(sum32'left) & sum32) + (sum33(sum33'left) & sum33(sum33'left) & sum33);
       sum41 <= (sum34(sum34'left) & sum34(sum34'left) & sum34) + (sum35(sum35'left) & sum35(sum35'left) & sum35) + (sum36(sum36'left) & sum36(sum36'left) & sum36) + (sum37(sum37'left) & sum37(sum37'left) & sum37);

       
       sum21 <= (sum17(sum17'left) & sum17(sum17'left) & sum17) + (sum18(sum18'left) & sum18(sum18'left) & sum18) + (sum19(sum19'left) & sum19(sum19'left) & sum19) + (sum20(sum20'left) & sum20(sum20'left) & sum20); 
       sum42 <= (sum38(sum38'left) & sum38(sum38'left) & sum38) + (sum39(sum39'left) & sum39(sum39'left) & sum39) + (sum40(sum40'left) & sum40(sum40'left) & sum40) + (sum41(sum41'left) & sum41(sum41'left) & sum41);

       sum43 <= (sum21(sum21'left) & sum21) + (sum42(sum42'left) & sum42);
    end if;
  end process p_sums;

d_out <= sum43(sum43'left downto sum43'left -W +1);

end a;