library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_SIGNED.ALL;

entity Huffman128 is
  generic (
           N             : integer := 4;  -- input data width
           M             : integer := 8;  -- max code width
           Wh            : integer := 16;  -- Huffman unit output data width (Note W>=M)
           Wb            : integer := 512; -- output buffer data width
           Huff_enc_en   : boolean := TRUE; -- Huffman encoder Enable/Bypass
           depth         : integer := 500; -- buffer depth
           burst         : integer := 10   -- buffer read burst
  	       );
  port    (
           clk           : in  std_logic;
           rst           : in  std_logic; 

           init_en       : in  std_logic;                         -- initialising convert table
           alpha_data    : in  std_logic_vector(N-1 downto 0);    
           alpha_code    : in  std_logic_vector(M-1 downto 0);    
           alpha_width   : in  std_logic_vector(  3 downto 0);

  	       d01_in          : in std_logic_vector (N-1 downto 0);
           d02_in          : in std_logic_vector (N-1 downto 0);
           d03_in          : in std_logic_vector (N-1 downto 0);
           d04_in          : in std_logic_vector (N-1 downto 0);
           d05_in          : in std_logic_vector (N-1 downto 0);
           d06_in          : in std_logic_vector (N-1 downto 0);
           d07_in          : in std_logic_vector (N-1 downto 0);
           d08_in          : in std_logic_vector (N-1 downto 0);
           d09_in          : in std_logic_vector (N-1 downto 0);
           d10_in          : in std_logic_vector (N-1 downto 0);
           d11_in          : in std_logic_vector (N-1 downto 0);
           d12_in          : in std_logic_vector (N-1 downto 0);
           d13_in          : in std_logic_vector (N-1 downto 0);
           d14_in          : in std_logic_vector (N-1 downto 0);
           d15_in          : in std_logic_vector (N-1 downto 0);
           d16_in          : in std_logic_vector (N-1 downto 0);
           d17_in          : in std_logic_vector (N-1 downto 0);
           d18_in          : in std_logic_vector (N-1 downto 0);
           d19_in          : in std_logic_vector (N-1 downto 0);
           d20_in          : in std_logic_vector (N-1 downto 0);
           d21_in          : in std_logic_vector (N-1 downto 0);
           d22_in          : in std_logic_vector (N-1 downto 0);
           d23_in          : in std_logic_vector (N-1 downto 0);
           d24_in          : in std_logic_vector (N-1 downto 0);
           d25_in          : in std_logic_vector (N-1 downto 0);
           d26_in          : in std_logic_vector (N-1 downto 0);
           d27_in          : in std_logic_vector (N-1 downto 0);
           d28_in          : in std_logic_vector (N-1 downto 0);
           d29_in          : in std_logic_vector (N-1 downto 0);
           d30_in          : in std_logic_vector (N-1 downto 0);
           d31_in          : in std_logic_vector (N-1 downto 0);
           d32_in          : in std_logic_vector (N-1 downto 0);
           d33_in          : in std_logic_vector (N-1 downto 0);
           d34_in          : in std_logic_vector (N-1 downto 0);
           d35_in          : in std_logic_vector (N-1 downto 0);
           d36_in          : in std_logic_vector (N-1 downto 0);
           d37_in          : in std_logic_vector (N-1 downto 0);
           d38_in          : in std_logic_vector (N-1 downto 0);
           d39_in          : in std_logic_vector (N-1 downto 0);
           d40_in          : in std_logic_vector (N-1 downto 0);
           d41_in          : in std_logic_vector (N-1 downto 0);
           d42_in          : in std_logic_vector (N-1 downto 0);
           d43_in          : in std_logic_vector (N-1 downto 0);
           d44_in          : in std_logic_vector (N-1 downto 0);
           d45_in          : in std_logic_vector (N-1 downto 0);
           d46_in          : in std_logic_vector (N-1 downto 0);
           d47_in          : in std_logic_vector (N-1 downto 0);
           d48_in          : in std_logic_vector (N-1 downto 0);
           d49_in          : in std_logic_vector (N-1 downto 0);
           d50_in          : in std_logic_vector (N-1 downto 0);
           d51_in          : in std_logic_vector (N-1 downto 0);
           d52_in          : in std_logic_vector (N-1 downto 0);
           d53_in          : in std_logic_vector (N-1 downto 0);
           d54_in          : in std_logic_vector (N-1 downto 0);
           d55_in          : in std_logic_vector (N-1 downto 0);
           d56_in          : in std_logic_vector (N-1 downto 0);
           d57_in          : in std_logic_vector (N-1 downto 0);
           d58_in          : in std_logic_vector (N-1 downto 0);
           d59_in          : in std_logic_vector (N-1 downto 0);
           d60_in          : in std_logic_vector (N-1 downto 0);
           d61_in          : in std_logic_vector (N-1 downto 0);
           d62_in          : in std_logic_vector (N-1 downto 0);
           d63_in          : in std_logic_vector (N-1 downto 0);
           d64_in          : in std_logic_vector (N-1 downto 0);

           d65_in          : in std_logic_vector (N-1 downto 0);
           d66_in          : in std_logic_vector (N-1 downto 0);
           d67_in          : in std_logic_vector (N-1 downto 0);
           d68_in          : in std_logic_vector (N-1 downto 0);
           d69_in          : in std_logic_vector (N-1 downto 0);
           d70_in          : in std_logic_vector (N-1 downto 0);
           d71_in          : in std_logic_vector (N-1 downto 0);
           d72_in          : in std_logic_vector (N-1 downto 0);
           d73_in          : in std_logic_vector (N-1 downto 0);
           d74_in          : in std_logic_vector (N-1 downto 0);
           d75_in          : in std_logic_vector (N-1 downto 0);
           d76_in          : in std_logic_vector (N-1 downto 0);
           d77_in          : in std_logic_vector (N-1 downto 0);
           d78_in          : in std_logic_vector (N-1 downto 0);
           d79_in          : in std_logic_vector (N-1 downto 0);
           d80_in          : in std_logic_vector (N-1 downto 0);
           d81_in          : in std_logic_vector (N-1 downto 0);
           d82_in          : in std_logic_vector (N-1 downto 0);
           d83_in          : in std_logic_vector (N-1 downto 0);
           d84_in          : in std_logic_vector (N-1 downto 0);
           d85_in          : in std_logic_vector (N-1 downto 0);
           d86_in          : in std_logic_vector (N-1 downto 0);
           d87_in          : in std_logic_vector (N-1 downto 0);
           d88_in          : in std_logic_vector (N-1 downto 0);
           d89_in          : in std_logic_vector (N-1 downto 0);
           d90_in          : in std_logic_vector (N-1 downto 0);
           d91_in          : in std_logic_vector (N-1 downto 0);
           d92_in          : in std_logic_vector (N-1 downto 0);
           d93_in          : in std_logic_vector (N-1 downto 0);
           d94_in          : in std_logic_vector (N-1 downto 0);
           d95_in          : in std_logic_vector (N-1 downto 0);
           d96_in          : in std_logic_vector (N-1 downto 0);
           d97_in          : in std_logic_vector (N-1 downto 0);
           d98_in          : in std_logic_vector (N-1 downto 0);
           d99_in          : in std_logic_vector (N-1 downto 0);
           d100_in         : in std_logic_vector (N-1 downto 0);
           d101_in         : in std_logic_vector (N-1 downto 0);
           d102_in         : in std_logic_vector (N-1 downto 0);
           d103_in         : in std_logic_vector (N-1 downto 0);
           d104_in         : in std_logic_vector (N-1 downto 0);
           d105_in         : in std_logic_vector (N-1 downto 0);
           d106_in         : in std_logic_vector (N-1 downto 0);
           d107_in         : in std_logic_vector (N-1 downto 0);
           d108_in         : in std_logic_vector (N-1 downto 0);
           d109_in         : in std_logic_vector (N-1 downto 0);
           d110_in         : in std_logic_vector (N-1 downto 0);
           d111_in         : in std_logic_vector (N-1 downto 0);
           d112_in         : in std_logic_vector (N-1 downto 0);
           d113_in         : in std_logic_vector (N-1 downto 0);
           d114_in         : in std_logic_vector (N-1 downto 0);
           d115_in         : in std_logic_vector (N-1 downto 0);
           d116_in         : in std_logic_vector (N-1 downto 0);
           d117_in         : in std_logic_vector (N-1 downto 0);
           d118_in         : in std_logic_vector (N-1 downto 0);
           d119_in         : in std_logic_vector (N-1 downto 0);
           d120_in         : in std_logic_vector (N-1 downto 0);
           d121_in         : in std_logic_vector (N-1 downto 0);
           d122_in         : in std_logic_vector (N-1 downto 0);
           d123_in         : in std_logic_vector (N-1 downto 0);
           d124_in         : in std_logic_vector (N-1 downto 0);
           d125_in         : in std_logic_vector (N-1 downto 0);
           d126_in         : in std_logic_vector (N-1 downto 0);
           d127_in         : in std_logic_vector (N-1 downto 0);
           d128_in         : in std_logic_vector (N-1 downto 0);

  	       en_in         : in  std_logic;
  	       sof_in        : in  std_logic;                         -- start of frame
           eof_in        : in  std_logic;                         -- end of frame

           buf_rd        : in  std_logic;
           buf_num       : in  std_logic_vector (6      downto 0);
           d_out         : out std_logic_vector (Wb  -1 downto 0);
           en_out        : out std_logic_vector (128  -1 downto 0);
           eof_out       : out std_logic);                        -- huffman code output
end Huffman128;

architecture a of Huffman128 is


component Huffman is
  generic (
           N             : integer := 4; -- input data width
           M             : integer := 8; -- max code width
           W             : integer := 10 -- output data width (Note W>=M)
           );
  port    (
           clk           : in  std_logic;
           rst           : in  std_logic; 

           init_en       : in  std_logic;                         -- initialising convert table
           alpha_data    : in  std_logic_vector(N-1 downto 0);    
           alpha_code    : in  std_logic_vector(M-1 downto 0);    
           alpha_width   : in  std_logic_vector(  3 downto 0);

           d_in          : in  std_logic_vector (N-1 downto 0);   -- data to convert
           en_in         : in  std_logic;
           sof_in        : in  std_logic;                         -- start of frame
           eof_in        : in  std_logic;                         -- end of frame

           d_out         : out std_logic_vector (W-1 downto 0);
           en_out        : out std_logic;
           eof_out       : out std_logic);                        -- huffman codde output
end component;

component fifo is
generic (depth   : integer := 16 ;
         burst   : integer := 10 ;  -- indication for burst read (Note, depth>burst) 
         Win     : integer := 16 ;
         Wout    : integer := 64 );  --depth of fifo
port (    clk        : in std_logic;
          rst        : in std_logic;
          enr        : in std_logic;   --enable read,should be '0' when not in use.
          enw        : in std_logic;    --enable write,should be '0' when not in use.
          data_in    : in std_logic_vector  (Win -1 downto 0);     --input data
          data_out   : out std_logic_vector(Wout-1 downto 0);    --output data
          burst_r    : out std_logic;   --set as '1' when the queue is ready for burst transaction
          fifo_empty : out std_logic;   --set as '1' when the queue is empty
          fifo_full  : out std_logic     --set as '1' when the queue is full
         );
end component;

signal h01_out, h65_out     : std_logic_vector(Wh-1 downto 0);
signal h02_out, h66_out     : std_logic_vector(Wh-1 downto 0);
signal h03_out, h67_out     : std_logic_vector(Wh-1 downto 0);
signal h04_out, h68_out     : std_logic_vector(Wh-1 downto 0);
signal h05_out, h69_out     : std_logic_vector(Wh-1 downto 0);
signal h06_out, h70_out     : std_logic_vector(Wh-1 downto 0);
signal h07_out, h71_out     : std_logic_vector(Wh-1 downto 0);
signal h08_out, h72_out     : std_logic_vector(Wh-1 downto 0);
signal h09_out, h73_out     : std_logic_vector(Wh-1 downto 0);
signal h10_out, h74_out     : std_logic_vector(Wh-1 downto 0);
signal h11_out, h75_out     : std_logic_vector(Wh-1 downto 0);
signal h12_out, h76_out     : std_logic_vector(Wh-1 downto 0);
signal h13_out, h77_out     : std_logic_vector(Wh-1 downto 0);
signal h14_out, h78_out     : std_logic_vector(Wh-1 downto 0);
signal h15_out, h79_out     : std_logic_vector(Wh-1 downto 0);
signal h16_out, h80_out     : std_logic_vector(Wh-1 downto 0);
signal h17_out, h81_out     : std_logic_vector(Wh-1 downto 0);
signal h18_out, h82_out     : std_logic_vector(Wh-1 downto 0);
signal h19_out, h83_out     : std_logic_vector(Wh-1 downto 0);
signal h20_out, h84_out     : std_logic_vector(Wh-1 downto 0);
signal h21_out, h85_out     : std_logic_vector(Wh-1 downto 0);
signal h22_out, h86_out     : std_logic_vector(Wh-1 downto 0);
signal h23_out, h87_out     : std_logic_vector(Wh-1 downto 0);
signal h24_out, h88_out     : std_logic_vector(Wh-1 downto 0);
signal h25_out, h89_out     : std_logic_vector(Wh-1 downto 0);
signal h26_out, h90_out     : std_logic_vector(Wh-1 downto 0);
signal h27_out, h91_out     : std_logic_vector(Wh-1 downto 0);
signal h28_out, h92_out     : std_logic_vector(Wh-1 downto 0);
signal h29_out, h93_out     : std_logic_vector(Wh-1 downto 0);
signal h30_out, h94_out     : std_logic_vector(Wh-1 downto 0);
signal h31_out, h95_out     : std_logic_vector(Wh-1 downto 0);
signal h32_out, h96_out     : std_logic_vector(Wh-1 downto 0);
signal h33_out, h97_out     : std_logic_vector(Wh-1 downto 0);
signal h34_out, h98_out     : std_logic_vector(Wh-1 downto 0);
signal h35_out, h99_out     : std_logic_vector(Wh-1 downto 0);
signal h36_out, h100_out    : std_logic_vector(Wh-1 downto 0);
signal h37_out, h101_out    : std_logic_vector(Wh-1 downto 0);
signal h38_out, h102_out    : std_logic_vector(Wh-1 downto 0);
signal h39_out, h103_out    : std_logic_vector(Wh-1 downto 0);
signal h40_out, h104_out    : std_logic_vector(Wh-1 downto 0);
signal h41_out, h105_out    : std_logic_vector(Wh-1 downto 0);
signal h42_out, h106_out    : std_logic_vector(Wh-1 downto 0);
signal h43_out, h107_out    : std_logic_vector(Wh-1 downto 0);
signal h44_out, h108_out    : std_logic_vector(Wh-1 downto 0);
signal h45_out, h109_out    : std_logic_vector(Wh-1 downto 0);
signal h46_out, h110_out    : std_logic_vector(Wh-1 downto 0);
signal h47_out, h111_out    : std_logic_vector(Wh-1 downto 0);
signal h48_out, h112_out    : std_logic_vector(Wh-1 downto 0);
signal h49_out, h113_out    : std_logic_vector(Wh-1 downto 0);
signal h50_out, h114_out    : std_logic_vector(Wh-1 downto 0);
signal h51_out, h115_out    : std_logic_vector(Wh-1 downto 0);
signal h52_out, h116_out    : std_logic_vector(Wh-1 downto 0);
signal h53_out, h117_out    : std_logic_vector(Wh-1 downto 0);
signal h54_out, h118_out    : std_logic_vector(Wh-1 downto 0);
signal h55_out, h119_out    : std_logic_vector(Wh-1 downto 0);
signal h56_out, h120_out    : std_logic_vector(Wh-1 downto 0);
signal h57_out, h121_out    : std_logic_vector(Wh-1 downto 0);
signal h58_out, h122_out    : std_logic_vector(Wh-1 downto 0);
signal h59_out, h123_out    : std_logic_vector(Wh-1 downto 0);
signal h60_out, h124_out    : std_logic_vector(Wh-1 downto 0);
signal h61_out, h125_out    : std_logic_vector(Wh-1 downto 0);
signal h62_out, h126_out    : std_logic_vector(Wh-1 downto 0);
signal h63_out, h127_out    : std_logic_vector(Wh-1 downto 0);
signal h64_out, h128_out    : std_logic_vector(Wh-1 downto 0);

signal h01_en, h65_en     : std_logic;
signal h02_en, h66_en     : std_logic;
signal h03_en, h67_en     : std_logic;
signal h04_en, h68_en     : std_logic;
signal h05_en, h69_en     : std_logic;
signal h06_en, h70_en     : std_logic;
signal h07_en, h71_en     : std_logic;
signal h08_en, h72_en     : std_logic;
signal h09_en, h73_en     : std_logic;
signal h10_en, h74_en     : std_logic;
signal h11_en, h75_en     : std_logic;
signal h12_en, h76_en     : std_logic;
signal h13_en, h77_en     : std_logic;
signal h14_en, h78_en     : std_logic;
signal h15_en, h79_en     : std_logic;
signal h16_en, h80_en     : std_logic;
signal h17_en, h81_en     : std_logic;
signal h18_en, h82_en     : std_logic;
signal h19_en, h83_en     : std_logic;
signal h20_en, h84_en     : std_logic;
signal h21_en, h85_en     : std_logic;
signal h22_en, h86_en     : std_logic;
signal h23_en, h87_en     : std_logic;
signal h24_en, h88_en     : std_logic;
signal h25_en, h89_en     : std_logic;
signal h26_en, h90_en     : std_logic;
signal h27_en, h91_en     : std_logic;
signal h28_en, h92_en     : std_logic;
signal h29_en, h93_en     : std_logic;
signal h30_en, h94_en     : std_logic;
signal h31_en, h95_en     : std_logic;
signal h32_en, h96_en     : std_logic;
signal h33_en, h97_en     : std_logic;
signal h34_en, h98_en     : std_logic;
signal h35_en, h99_en     : std_logic;
signal h36_en, h100_en    : std_logic;
signal h37_en, h101_en    : std_logic;
signal h38_en, h102_en    : std_logic;
signal h39_en, h103_en    : std_logic;
signal h40_en, h104_en    : std_logic;
signal h41_en, h105_en    : std_logic;
signal h42_en, h106_en    : std_logic;
signal h43_en, h107_en    : std_logic;
signal h44_en, h108_en    : std_logic;
signal h45_en, h109_en    : std_logic;
signal h46_en, h110_en    : std_logic;
signal h47_en, h111_en    : std_logic;
signal h48_en, h112_en    : std_logic;
signal h49_en, h113_en    : std_logic;
signal h50_en, h114_en    : std_logic;
signal h51_en, h115_en    : std_logic;
signal h52_en, h116_en    : std_logic;
signal h53_en, h117_en    : std_logic;
signal h54_en, h118_en    : std_logic;
signal h55_en, h119_en    : std_logic;
signal h56_en, h120_en    : std_logic;
signal h57_en, h121_en    : std_logic;
signal h58_en, h122_en    : std_logic;
signal h59_en, h123_en    : std_logic;
signal h60_en, h124_en    : std_logic;
signal h61_en, h125_en    : std_logic;
signal h62_en, h126_en    : std_logic;
signal h63_en, h127_en    : std_logic;
signal h64_en, h128_en    : std_logic;

signal buff01_out, buff02_out, buff03_out, buff04_out, buff05_out, buff06_out, buff07_out, buff08_out, buff09_out, buff10_out, buff11_out, buff12_out, buff13_out, buff14_out, buff15_out, buff16_out, buff17_out, buff18_out, buff19_out, buff20_out, buff21_out, buff22_out, buff23_out, buff24_out, buff25_out, buff26_out, buff27_out, buff28_out, buff29_out, buff30_out, buff31_out, buff32_out : std_logic_vector(Wb-1 downto 0);
signal buff33_out, buff34_out, buff35_out, buff36_out, buff37_out, buff38_out, buff39_out, buff40_out, buff41_out, buff42_out, buff43_out, buff44_out, buff45_out, buff46_out, buff47_out, buff48_out, buff49_out, buff50_out, buff51_out, buff52_out, buff53_out, buff54_out, buff55_out, buff56_out, buff57_out, buff58_out, buff59_out, buff60_out, buff61_out, buff62_out, buff63_out, buff64_out : std_logic_vector(Wb-1 downto 0);
signal buff65_out, buff66_out, buff67_out, buff68_out, buff69_out, buff70_out, buff71_out, buff72_out, buff73_out, buff74_out, buff75_out, buff76_out, buff77_out, buff78_out, buff79_out, buff80_out, buff81_out, buff82_out, buff83_out, buff84_out, buff85_out, buff86_out, buff87_out, buff88_out, buff89_out, buff90_out, buff91_out, buff92_out, buff93_out, buff94_out, buff95_out, buff96_out : std_logic_vector(Wb-1 downto 0);
signal buff97_out, buff98_out, buff99_out, buff100_out, buff101_out, buff102_out, buff103_out, buff104_out, buff105_out, buff106_out, buff107_out, buff108_out, buff109_out, buff110_out, buff111_out, buff112_out, buff113_out, buff114_out, buff115_out, buff116_out, buff117_out, buff118_out, buff119_out, buff120_out, buff121_out, buff122_out, buff123_out, buff124_out, buff125_out, buff126_out, buff127_out, buff128_out : std_logic_vector(Wb-1 downto 0);

signal b_rd : std_logic_vector (128-1 downto 0);

begin

g_Huff_enc_en: if Huff_enc_en = TRUE generate
   Huf01 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d01_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h01_out, en_out => h01_en, eof_out => eof_out);
   Huf02 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d02_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h02_out, en_out => h02_en, eof_out => open);
   Huf03 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d03_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h03_out, en_out => h03_en, eof_out => open);
   Huf04 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d04_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h04_out, en_out => h04_en, eof_out => open);
   Huf05 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d05_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h05_out, en_out => h05_en, eof_out => open);
   Huf06 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d06_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h06_out, en_out => h06_en, eof_out => open);
   Huf07 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d07_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h07_out, en_out => h07_en, eof_out => open);
   Huf08 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d08_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h08_out, en_out => h08_en, eof_out => open);
   Huf09 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d09_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h09_out, en_out => h09_en, eof_out => open);
   Huf10 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d10_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h10_out, en_out => h10_en, eof_out => open);
   Huf11 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d11_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h11_out, en_out => h11_en, eof_out => open);
   Huf12 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d12_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h12_out, en_out => h12_en, eof_out => open);
   Huf13 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d13_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h13_out, en_out => h13_en, eof_out => open);
   Huf14 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d14_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h14_out, en_out => h14_en, eof_out => open);
   Huf15 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d15_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h15_out, en_out => h15_en, eof_out => open);
   Huf16 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d16_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h16_out, en_out => h16_en, eof_out => open);
   Huf17 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d17_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h17_out, en_out => h17_en, eof_out => open);
   Huf18 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d18_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h18_out, en_out => h18_en, eof_out => open);
   Huf19 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d19_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h19_out, en_out => h19_en, eof_out => open);
   Huf20 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d20_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h20_out, en_out => h20_en, eof_out => open);
   Huf21 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d21_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h21_out, en_out => h21_en, eof_out => open);
   Huf22 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d22_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h22_out, en_out => h22_en, eof_out => open);
   Huf23 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d23_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h23_out, en_out => h23_en, eof_out => open);
   Huf24 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d24_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h24_out, en_out => h24_en, eof_out => open);
   Huf25 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d25_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h25_out, en_out => h25_en, eof_out => open);
   Huf26 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d26_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h26_out, en_out => h26_en, eof_out => open);
   Huf27 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d27_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h27_out, en_out => h27_en, eof_out => open);
   Huf28 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d28_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h28_out, en_out => h28_en, eof_out => open);
   Huf29 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d29_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h29_out, en_out => h29_en, eof_out => open);
   Huf30 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d30_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h30_out, en_out => h30_en, eof_out => open);
   Huf31 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d31_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h31_out, en_out => h31_en, eof_out => open);
   Huf32 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d32_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h32_out, en_out => h32_en, eof_out => open);
   Huf33 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d33_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h33_out, en_out => h33_en, eof_out => open);
   Huf34 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d34_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h34_out, en_out => h34_en, eof_out => open);
   Huf35 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d35_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h35_out, en_out => h35_en, eof_out => open);
   Huf36 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d36_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h36_out, en_out => h36_en, eof_out => open);
   Huf37 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d37_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h37_out, en_out => h37_en, eof_out => open);
   Huf38 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d38_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h38_out, en_out => h38_en, eof_out => open);
   Huf39 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d39_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h39_out, en_out => h39_en, eof_out => open);
   Huf40 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d40_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h40_out, en_out => h40_en, eof_out => open);
   Huf41 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d41_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h41_out, en_out => h41_en, eof_out => open);
   Huf42 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d42_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h42_out, en_out => h42_en, eof_out => open);
   Huf43 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d43_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h43_out, en_out => h43_en, eof_out => open);
   Huf44 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d44_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h44_out, en_out => h44_en, eof_out => open);
   Huf45 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d45_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h45_out, en_out => h45_en, eof_out => open);
   Huf46 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d46_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h46_out, en_out => h46_en, eof_out => open);
   Huf47 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d47_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h47_out, en_out => h47_en, eof_out => open);
   Huf48 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d48_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h48_out, en_out => h48_en, eof_out => open);
   Huf49 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d49_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h49_out, en_out => h49_en, eof_out => open);
   Huf50 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d50_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h50_out, en_out => h50_en, eof_out => open);
   Huf51 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d51_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h51_out, en_out => h51_en, eof_out => open);
   Huf52 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d52_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h52_out, en_out => h52_en, eof_out => open);
   Huf53 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d53_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h53_out, en_out => h53_en, eof_out => open);
   Huf54 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d54_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h54_out, en_out => h54_en, eof_out => open);
   Huf55 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d55_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h55_out, en_out => h55_en, eof_out => open);
   Huf56 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d56_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h56_out, en_out => h56_en, eof_out => open);
   Huf57 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d57_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h57_out, en_out => h57_en, eof_out => open);
   Huf58 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d58_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h58_out, en_out => h58_en, eof_out => open);
   Huf59 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d59_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h59_out, en_out => h59_en, eof_out => open);
   Huf60 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d60_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h60_out, en_out => h60_en, eof_out => open);
   Huf61 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d61_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h61_out, en_out => h61_en, eof_out => open);
   Huf62 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d62_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h62_out, en_out => h62_en, eof_out => open);
   Huf63 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d63_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h63_out, en_out => h63_en, eof_out => open);
   Huf64 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d64_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h64_out, en_out => h64_en, eof_out => open);

   Huf65 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d65_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h65_out , en_out => h65_en , eof_out => open);
   Huf66 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d66_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h66_out , en_out => h66_en , eof_out => open);
   Huf67 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d67_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h67_out , en_out => h67_en , eof_out => open);
   Huf68 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d68_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h68_out , en_out => h68_en , eof_out => open);
   Huf69 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d69_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h69_out , en_out => h69_en , eof_out => open);
   Huf70 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d70_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h70_out , en_out => h70_en , eof_out => open);
   Huf71 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d71_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h71_out , en_out => h71_en , eof_out => open);
   Huf72 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d72_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h72_out , en_out => h72_en , eof_out => open);
   Huf73 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d73_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h73_out , en_out => h73_en , eof_out => open);
   Huf74 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d74_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h74_out , en_out => h74_en , eof_out => open);
   Huf75 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d75_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h75_out , en_out => h75_en , eof_out => open);
   Huf76 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d76_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h76_out , en_out => h76_en , eof_out => open);
   Huf77 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d77_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h77_out , en_out => h77_en , eof_out => open);
   Huf78 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d78_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h78_out , en_out => h78_en , eof_out => open);
   Huf79 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d79_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h79_out , en_out => h79_en , eof_out => open);
   Huf80 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d80_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h80_out , en_out => h80_en , eof_out => open);
   Huf81 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d81_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h81_out , en_out => h81_en , eof_out => open);
   Huf82 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d82_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h82_out , en_out => h82_en , eof_out => open);
   Huf83 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d83_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h83_out , en_out => h83_en , eof_out => open);
   Huf84 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d84_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h84_out , en_out => h84_en , eof_out => open);
   Huf85 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d85_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h85_out , en_out => h85_en , eof_out => open);
   Huf86 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d86_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h86_out , en_out => h86_en , eof_out => open);
   Huf87 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d87_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h87_out , en_out => h87_en , eof_out => open);
   Huf88 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d88_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h88_out , en_out => h88_en , eof_out => open);
   Huf89 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d89_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h89_out , en_out => h89_en , eof_out => open);
   Huf90 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d90_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h90_out , en_out => h90_en , eof_out => open);
   Huf91 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d91_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h91_out , en_out => h91_en , eof_out => open);
   Huf92 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d92_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h92_out , en_out => h92_en , eof_out => open);
   Huf93 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d93_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h93_out , en_out => h93_en , eof_out => open);
   Huf94 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d94_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h94_out , en_out => h94_en , eof_out => open);
   Huf95 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d95_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h95_out , en_out => h95_en , eof_out => open);
   Huf96 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d96_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h96_out , en_out => h96_en , eof_out => open);
   Huf97 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d97_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h97_out , en_out => h97_en , eof_out => open);
   Huf98 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d98_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h98_out , en_out => h98_en , eof_out => open);
   Huf99 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d99_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h99_out , en_out => h99_en , eof_out => open);
   Huf100: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d100_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h100_out, en_out => h100_en, eof_out => open);
   Huf101: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d101_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h101_out, en_out => h101_en, eof_out => open);
   Huf102: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d102_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h102_out, en_out => h102_en, eof_out => open);
   Huf103: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d103_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h103_out, en_out => h103_en, eof_out => open);
   Huf104: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d104_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h104_out, en_out => h104_en, eof_out => open);
   Huf105: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d105_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h105_out, en_out => h105_en, eof_out => open);
   Huf106: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d106_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h106_out, en_out => h106_en, eof_out => open);
   Huf107: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d107_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h107_out, en_out => h107_en, eof_out => open);
   Huf108: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d108_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h108_out, en_out => h108_en, eof_out => open);
   Huf109: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d109_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h109_out, en_out => h109_en, eof_out => open);
   Huf110: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d110_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h110_out, en_out => h110_en, eof_out => open);
   Huf111: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d111_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h111_out, en_out => h111_en, eof_out => open);
   Huf112: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d112_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h112_out, en_out => h112_en, eof_out => open);
   Huf113: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d113_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h113_out, en_out => h113_en, eof_out => open);
   Huf114: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d114_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h114_out, en_out => h114_en, eof_out => open);
   Huf115: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d115_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h115_out, en_out => h115_en, eof_out => open);
   Huf116: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d116_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h116_out, en_out => h116_en, eof_out => open);
   Huf117: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d117_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h117_out, en_out => h117_en, eof_out => open);
   Huf118: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d118_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h118_out, en_out => h118_en, eof_out => open);
   Huf119: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d119_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h119_out, en_out => h119_en, eof_out => open);
   Huf120: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d120_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h120_out, en_out => h120_en, eof_out => open);
   Huf121: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d121_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h121_out, en_out => h121_en, eof_out => open);
   Huf122: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d122_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h122_out, en_out => h122_en, eof_out => open);
   Huf123: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d123_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h123_out, en_out => h123_en, eof_out => open);
   Huf124: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d124_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h124_out, en_out => h124_en, eof_out => open);
   Huf125: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d125_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h125_out, en_out => h125_en, eof_out => open);
   Huf126: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d126_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h126_out, en_out => h126_en, eof_out => open);
   Huf127: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d127_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h127_out, en_out => h127_en, eof_out => open);
   Huf128: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d128_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h128_out, en_out => h128_en, eof_out => open);
end generate g_Huff_enc_en;

g_Huff_enc_dis: if Huff_enc_en = FALSE generate
   h01_out(h01_out'left downto d01_in'left + 1) <= (others => '0');   h01_out(d01_in'left downto 0) <= d01_in;   h01_en <= en_in;
   h02_out(h02_out'left downto d02_in'left + 1) <= (others => '0');   h02_out(d02_in'left downto 0) <= d02_in;   h02_en <= en_in;
   h03_out(h03_out'left downto d03_in'left + 1) <= (others => '0');   h03_out(d03_in'left downto 0) <= d03_in;   h03_en <= en_in;
   h04_out(h04_out'left downto d04_in'left + 1) <= (others => '0');   h04_out(d04_in'left downto 0) <= d04_in;   h04_en <= en_in;
   h05_out(h05_out'left downto d05_in'left + 1) <= (others => '0');   h05_out(d05_in'left downto 0) <= d05_in;   h05_en <= en_in;
   h06_out(h06_out'left downto d06_in'left + 1) <= (others => '0');   h06_out(d06_in'left downto 0) <= d06_in;   h06_en <= en_in;
   h07_out(h07_out'left downto d07_in'left + 1) <= (others => '0');   h07_out(d07_in'left downto 0) <= d07_in;   h07_en <= en_in;
   h08_out(h08_out'left downto d08_in'left + 1) <= (others => '0');   h08_out(d08_in'left downto 0) <= d08_in;   h08_en <= en_in;
   h09_out(h09_out'left downto d09_in'left + 1) <= (others => '0');   h09_out(d09_in'left downto 0) <= d09_in;   h09_en <= en_in;
   h10_out(h10_out'left downto d10_in'left + 1) <= (others => '0');   h10_out(d10_in'left downto 0) <= d10_in;   h10_en <= en_in;
   h11_out(h11_out'left downto d11_in'left + 1) <= (others => '0');   h11_out(d11_in'left downto 0) <= d11_in;   h11_en <= en_in;
   h12_out(h12_out'left downto d12_in'left + 1) <= (others => '0');   h12_out(d12_in'left downto 0) <= d12_in;   h12_en <= en_in;
   h13_out(h13_out'left downto d13_in'left + 1) <= (others => '0');   h13_out(d13_in'left downto 0) <= d13_in;   h13_en <= en_in;
   h14_out(h14_out'left downto d14_in'left + 1) <= (others => '0');   h14_out(d14_in'left downto 0) <= d14_in;   h14_en <= en_in;
   h15_out(h15_out'left downto d15_in'left + 1) <= (others => '0');   h15_out(d15_in'left downto 0) <= d15_in;   h15_en <= en_in;
   h16_out(h16_out'left downto d16_in'left + 1) <= (others => '0');   h16_out(d16_in'left downto 0) <= d16_in;   h16_en <= en_in;
   h17_out(h17_out'left downto d17_in'left + 1) <= (others => '0');   h17_out(d17_in'left downto 0) <= d17_in;   h17_en <= en_in;
   h18_out(h18_out'left downto d18_in'left + 1) <= (others => '0');   h18_out(d18_in'left downto 0) <= d18_in;   h18_en <= en_in;
   h19_out(h19_out'left downto d19_in'left + 1) <= (others => '0');   h19_out(d19_in'left downto 0) <= d19_in;   h19_en <= en_in;
   h20_out(h20_out'left downto d20_in'left + 1) <= (others => '0');   h20_out(d20_in'left downto 0) <= d20_in;   h20_en <= en_in;
   h21_out(h21_out'left downto d21_in'left + 1) <= (others => '0');   h21_out(d21_in'left downto 0) <= d21_in;   h21_en <= en_in;
   h22_out(h22_out'left downto d22_in'left + 1) <= (others => '0');   h22_out(d22_in'left downto 0) <= d22_in;   h22_en <= en_in;
   h23_out(h23_out'left downto d23_in'left + 1) <= (others => '0');   h23_out(d23_in'left downto 0) <= d23_in;   h23_en <= en_in;
   h24_out(h24_out'left downto d24_in'left + 1) <= (others => '0');   h24_out(d24_in'left downto 0) <= d24_in;   h24_en <= en_in;
   h25_out(h25_out'left downto d25_in'left + 1) <= (others => '0');   h25_out(d25_in'left downto 0) <= d25_in;   h25_en <= en_in;
   h26_out(h26_out'left downto d26_in'left + 1) <= (others => '0');   h26_out(d26_in'left downto 0) <= d26_in;   h26_en <= en_in;
   h27_out(h27_out'left downto d27_in'left + 1) <= (others => '0');   h27_out(d27_in'left downto 0) <= d27_in;   h27_en <= en_in;
   h28_out(h28_out'left downto d28_in'left + 1) <= (others => '0');   h28_out(d28_in'left downto 0) <= d28_in;   h28_en <= en_in;
   h29_out(h29_out'left downto d29_in'left + 1) <= (others => '0');   h29_out(d29_in'left downto 0) <= d29_in;   h29_en <= en_in;
   h30_out(h30_out'left downto d30_in'left + 1) <= (others => '0');   h30_out(d30_in'left downto 0) <= d30_in;   h30_en <= en_in;
   h31_out(h31_out'left downto d31_in'left + 1) <= (others => '0');   h31_out(d31_in'left downto 0) <= d31_in;   h31_en <= en_in;
   h32_out(h32_out'left downto d32_in'left + 1) <= (others => '0');   h32_out(d32_in'left downto 0) <= d32_in;   h32_en <= en_in;
   h33_out(h33_out'left downto d33_in'left + 1) <= (others => '0');   h33_out(d33_in'left downto 0) <= d33_in;   h33_en <= en_in;
   h34_out(h34_out'left downto d34_in'left + 1) <= (others => '0');   h34_out(d34_in'left downto 0) <= d34_in;   h34_en <= en_in;
   h35_out(h35_out'left downto d35_in'left + 1) <= (others => '0');   h35_out(d35_in'left downto 0) <= d35_in;   h35_en <= en_in;
   h36_out(h36_out'left downto d36_in'left + 1) <= (others => '0');   h36_out(d36_in'left downto 0) <= d36_in;   h36_en <= en_in;
   h37_out(h37_out'left downto d37_in'left + 1) <= (others => '0');   h37_out(d37_in'left downto 0) <= d37_in;   h37_en <= en_in;
   h38_out(h38_out'left downto d38_in'left + 1) <= (others => '0');   h38_out(d38_in'left downto 0) <= d38_in;   h38_en <= en_in;
   h39_out(h39_out'left downto d39_in'left + 1) <= (others => '0');   h39_out(d39_in'left downto 0) <= d39_in;   h39_en <= en_in;
   h40_out(h40_out'left downto d40_in'left + 1) <= (others => '0');   h40_out(d40_in'left downto 0) <= d40_in;   h40_en <= en_in;
   h41_out(h41_out'left downto d41_in'left + 1) <= (others => '0');   h41_out(d41_in'left downto 0) <= d41_in;   h41_en <= en_in;
   h42_out(h42_out'left downto d42_in'left + 1) <= (others => '0');   h42_out(d42_in'left downto 0) <= d42_in;   h42_en <= en_in;
   h43_out(h43_out'left downto d43_in'left + 1) <= (others => '0');   h43_out(d43_in'left downto 0) <= d43_in;   h43_en <= en_in;
   h44_out(h44_out'left downto d44_in'left + 1) <= (others => '0');   h44_out(d44_in'left downto 0) <= d44_in;   h44_en <= en_in;
   h45_out(h45_out'left downto d45_in'left + 1) <= (others => '0');   h45_out(d45_in'left downto 0) <= d45_in;   h45_en <= en_in;
   h46_out(h46_out'left downto d46_in'left + 1) <= (others => '0');   h46_out(d46_in'left downto 0) <= d46_in;   h46_en <= en_in;
   h47_out(h47_out'left downto d47_in'left + 1) <= (others => '0');   h47_out(d47_in'left downto 0) <= d47_in;   h47_en <= en_in;
   h48_out(h48_out'left downto d48_in'left + 1) <= (others => '0');   h48_out(d48_in'left downto 0) <= d48_in;   h48_en <= en_in;
   h49_out(h49_out'left downto d49_in'left + 1) <= (others => '0');   h49_out(d49_in'left downto 0) <= d49_in;   h49_en <= en_in;
   h50_out(h50_out'left downto d50_in'left + 1) <= (others => '0');   h50_out(d50_in'left downto 0) <= d50_in;   h50_en <= en_in;
   h51_out(h51_out'left downto d51_in'left + 1) <= (others => '0');   h51_out(d51_in'left downto 0) <= d51_in;   h51_en <= en_in;
   h52_out(h52_out'left downto d52_in'left + 1) <= (others => '0');   h52_out(d52_in'left downto 0) <= d52_in;   h52_en <= en_in;
   h53_out(h53_out'left downto d53_in'left + 1) <= (others => '0');   h53_out(d53_in'left downto 0) <= d53_in;   h53_en <= en_in;
   h54_out(h54_out'left downto d54_in'left + 1) <= (others => '0');   h54_out(d54_in'left downto 0) <= d54_in;   h54_en <= en_in;
   h55_out(h55_out'left downto d55_in'left + 1) <= (others => '0');   h55_out(d55_in'left downto 0) <= d55_in;   h55_en <= en_in;
   h56_out(h56_out'left downto d56_in'left + 1) <= (others => '0');   h56_out(d56_in'left downto 0) <= d56_in;   h56_en <= en_in;
   h57_out(h57_out'left downto d57_in'left + 1) <= (others => '0');   h57_out(d57_in'left downto 0) <= d57_in;   h57_en <= en_in;
   h58_out(h58_out'left downto d58_in'left + 1) <= (others => '0');   h58_out(d58_in'left downto 0) <= d58_in;   h58_en <= en_in;
   h59_out(h59_out'left downto d59_in'left + 1) <= (others => '0');   h59_out(d59_in'left downto 0) <= d59_in;   h59_en <= en_in;
   h60_out(h60_out'left downto d60_in'left + 1) <= (others => '0');   h60_out(d60_in'left downto 0) <= d60_in;   h60_en <= en_in;
   h61_out(h61_out'left downto d61_in'left + 1) <= (others => '0');   h61_out(d61_in'left downto 0) <= d61_in;   h61_en <= en_in;
   h62_out(h62_out'left downto d62_in'left + 1) <= (others => '0');   h62_out(d62_in'left downto 0) <= d62_in;   h62_en <= en_in;
   h63_out(h63_out'left downto d63_in'left + 1) <= (others => '0');   h63_out(d63_in'left downto 0) <= d63_in;   h63_en <= en_in;
   h64_out(h64_out'left downto d64_in'left + 1) <= (others => '0');   h64_out(d64_in'left downto 0) <= d64_in;   h64_en <= en_in;


   h65_out (h65_out 'left downto d65_in'left  + 1) <= (others => '0');   h65_out (d65_in 'left downto 0) <= d65_in;   h65_en  <= en_in;
   h66_out (h66_out 'left downto d66_in'left  + 1) <= (others => '0');   h66_out (d66_in 'left downto 0) <= d66_in;   h66_en  <= en_in;
   h67_out (h67_out 'left downto d67_in'left  + 1) <= (others => '0');   h67_out (d67_in 'left downto 0) <= d67_in;   h67_en  <= en_in;
   h68_out (h68_out 'left downto d68_in'left  + 1) <= (others => '0');   h68_out (d68_in 'left downto 0) <= d68_in;   h68_en  <= en_in;
   h69_out (h69_out 'left downto d69_in'left  + 1) <= (others => '0');   h69_out (d69_in 'left downto 0) <= d69_in;   h69_en  <= en_in;
   h70_out (h70_out 'left downto d70_in'left  + 1) <= (others => '0');   h70_out (d70_in 'left downto 0) <= d70_in;   h70_en  <= en_in;
   h71_out (h71_out 'left downto d71_in'left  + 1) <= (others => '0');   h71_out (d71_in 'left downto 0) <= d71_in;   h71_en  <= en_in;
   h72_out (h72_out 'left downto d72_in'left  + 1) <= (others => '0');   h72_out (d72_in 'left downto 0) <= d72_in;   h72_en  <= en_in;
   h73_out (h73_out 'left downto d73_in'left  + 1) <= (others => '0');   h73_out (d73_in 'left downto 0) <= d73_in;   h73_en  <= en_in;
   h74_out (h74_out 'left downto d74_in'left  + 1) <= (others => '0');   h74_out (d74_in 'left downto 0) <= d74_in;   h74_en  <= en_in;
   h75_out (h75_out 'left downto d75_in'left  + 1) <= (others => '0');   h75_out (d75_in 'left downto 0) <= d75_in;   h75_en  <= en_in;
   h76_out (h76_out 'left downto d76_in'left  + 1) <= (others => '0');   h76_out (d76_in 'left downto 0) <= d76_in;   h76_en  <= en_in;
   h77_out (h77_out 'left downto d77_in'left  + 1) <= (others => '0');   h77_out (d77_in 'left downto 0) <= d77_in;   h77_en  <= en_in;
   h78_out (h78_out 'left downto d78_in'left  + 1) <= (others => '0');   h78_out (d78_in 'left downto 0) <= d78_in;   h78_en  <= en_in;
   h79_out (h79_out 'left downto d79_in'left  + 1) <= (others => '0');   h79_out (d79_in 'left downto 0) <= d79_in;   h79_en  <= en_in;
   h80_out (h80_out 'left downto d80_in'left  + 1) <= (others => '0');   h80_out (d80_in 'left downto 0) <= d80_in;   h80_en  <= en_in;
   h81_out (h81_out 'left downto d81_in'left  + 1) <= (others => '0');   h81_out (d81_in 'left downto 0) <= d81_in;   h81_en  <= en_in;
   h82_out (h82_out 'left downto d82_in'left  + 1) <= (others => '0');   h82_out (d82_in 'left downto 0) <= d82_in;   h82_en  <= en_in;
   h83_out (h83_out 'left downto d83_in'left  + 1) <= (others => '0');   h83_out (d83_in 'left downto 0) <= d83_in;   h83_en  <= en_in;
   h84_out (h84_out 'left downto d84_in'left  + 1) <= (others => '0');   h84_out (d84_in 'left downto 0) <= d84_in;   h84_en  <= en_in;
   h85_out (h85_out 'left downto d85_in'left  + 1) <= (others => '0');   h85_out (d85_in 'left downto 0) <= d85_in;   h85_en  <= en_in;
   h86_out (h86_out 'left downto d86_in'left  + 1) <= (others => '0');   h86_out (d86_in 'left downto 0) <= d86_in;   h86_en  <= en_in;
   h87_out (h87_out 'left downto d87_in'left  + 1) <= (others => '0');   h87_out (d87_in 'left downto 0) <= d87_in;   h87_en  <= en_in;
   h88_out (h88_out 'left downto d88_in'left  + 1) <= (others => '0');   h88_out (d88_in 'left downto 0) <= d88_in;   h88_en  <= en_in;
   h89_out (h89_out 'left downto d89_in'left  + 1) <= (others => '0');   h89_out (d89_in 'left downto 0) <= d89_in;   h89_en  <= en_in;
   h90_out (h90_out 'left downto d90_in'left  + 1) <= (others => '0');   h90_out (d90_in 'left downto 0) <= d90_in;   h90_en  <= en_in;
   h91_out (h91_out 'left downto d91_in'left  + 1) <= (others => '0');   h91_out (d91_in 'left downto 0) <= d91_in;   h91_en  <= en_in;
   h92_out (h92_out 'left downto d92_in'left  + 1) <= (others => '0');   h92_out (d92_in 'left downto 0) <= d92_in;   h92_en  <= en_in;
   h93_out (h93_out 'left downto d93_in'left  + 1) <= (others => '0');   h93_out (d93_in 'left downto 0) <= d93_in;   h93_en  <= en_in;
   h94_out (h94_out 'left downto d94_in'left  + 1) <= (others => '0');   h94_out (d94_in 'left downto 0) <= d94_in;   h94_en  <= en_in;
   h95_out (h95_out 'left downto d95_in'left  + 1) <= (others => '0');   h95_out (d95_in 'left downto 0) <= d95_in;   h95_en  <= en_in;
   h96_out (h96_out 'left downto d96_in'left  + 1) <= (others => '0');   h96_out (d96_in 'left downto 0) <= d96_in;   h96_en  <= en_in;
   h97_out (h97_out 'left downto d97_in'left  + 1) <= (others => '0');   h97_out (d97_in 'left downto 0) <= d97_in;   h97_en  <= en_in;
   h98_out (h98_out 'left downto d98_in'left  + 1) <= (others => '0');   h98_out (d98_in 'left downto 0) <= d98_in;   h98_en  <= en_in;
   h99_out (h99_out 'left downto d99_in'left  + 1) <= (others => '0');   h99_out (d99_in 'left downto 0) <= d99_in;   h99_en  <= en_in;
   h100_out(h100_out'left downto d100_in'left + 1) <= (others => '0');   h100_out(d100_in'left downto 0) <= d100_in;  h100_en <= en_in;
   h101_out(h101_out'left downto d101_in'left + 1) <= (others => '0');   h101_out(d101_in'left downto 0) <= d101_in;  h101_en <= en_in;
   h102_out(h102_out'left downto d102_in'left + 1) <= (others => '0');   h102_out(d102_in'left downto 0) <= d102_in;  h102_en <= en_in;
   h103_out(h103_out'left downto d103_in'left + 1) <= (others => '0');   h103_out(d103_in'left downto 0) <= d103_in;  h103_en <= en_in;
   h104_out(h104_out'left downto d104_in'left + 1) <= (others => '0');   h104_out(d104_in'left downto 0) <= d104_in;  h104_en <= en_in;
   h105_out(h105_out'left downto d105_in'left + 1) <= (others => '0');   h105_out(d105_in'left downto 0) <= d105_in;  h105_en <= en_in;
   h106_out(h106_out'left downto d106_in'left + 1) <= (others => '0');   h106_out(d106_in'left downto 0) <= d106_in;  h106_en <= en_in;
   h107_out(h107_out'left downto d107_in'left + 1) <= (others => '0');   h107_out(d107_in'left downto 0) <= d107_in;  h107_en <= en_in;
   h108_out(h108_out'left downto d108_in'left + 1) <= (others => '0');   h108_out(d108_in'left downto 0) <= d108_in;  h108_en <= en_in;
   h109_out(h109_out'left downto d109_in'left + 1) <= (others => '0');   h109_out(d109_in'left downto 0) <= d109_in;  h109_en <= en_in;
   h110_out(h110_out'left downto d110_in'left + 1) <= (others => '0');   h110_out(d110_in'left downto 0) <= d110_in;  h110_en <= en_in;
   h111_out(h111_out'left downto d111_in'left + 1) <= (others => '0');   h111_out(d111_in'left downto 0) <= d111_in;  h111_en <= en_in;
   h112_out(h112_out'left downto d112_in'left + 1) <= (others => '0');   h112_out(d112_in'left downto 0) <= d112_in;  h112_en <= en_in;
   h113_out(h113_out'left downto d113_in'left + 1) <= (others => '0');   h113_out(d113_in'left downto 0) <= d113_in;  h113_en <= en_in;
   h114_out(h114_out'left downto d114_in'left + 1) <= (others => '0');   h114_out(d114_in'left downto 0) <= d114_in;  h114_en <= en_in;
   h115_out(h115_out'left downto d115_in'left + 1) <= (others => '0');   h115_out(d115_in'left downto 0) <= d115_in;  h115_en <= en_in;
   h116_out(h116_out'left downto d116_in'left + 1) <= (others => '0');   h116_out(d116_in'left downto 0) <= d116_in;  h116_en <= en_in;
   h117_out(h117_out'left downto d117_in'left + 1) <= (others => '0');   h117_out(d117_in'left downto 0) <= d117_in;  h117_en <= en_in;
   h118_out(h118_out'left downto d118_in'left + 1) <= (others => '0');   h118_out(d118_in'left downto 0) <= d118_in;  h118_en <= en_in;
   h119_out(h119_out'left downto d119_in'left + 1) <= (others => '0');   h119_out(d119_in'left downto 0) <= d119_in;  h119_en <= en_in;
   h120_out(h120_out'left downto d120_in'left + 1) <= (others => '0');   h120_out(d120_in'left downto 0) <= d120_in;  h120_en <= en_in;
   h121_out(h121_out'left downto d121_in'left + 1) <= (others => '0');   h121_out(d121_in'left downto 0) <= d121_in;  h121_en <= en_in;
   h122_out(h122_out'left downto d122_in'left + 1) <= (others => '0');   h122_out(d122_in'left downto 0) <= d122_in;  h122_en <= en_in;
   h123_out(h123_out'left downto d123_in'left + 1) <= (others => '0');   h123_out(d123_in'left downto 0) <= d123_in;  h123_en <= en_in;
   h124_out(h124_out'left downto d124_in'left + 1) <= (others => '0');   h124_out(d124_in'left downto 0) <= d124_in;  h124_en <= en_in;
   h125_out(h125_out'left downto d125_in'left + 1) <= (others => '0');   h125_out(d125_in'left downto 0) <= d125_in;  h125_en <= en_in;
   h126_out(h126_out'left downto d126_in'left + 1) <= (others => '0');   h126_out(d126_in'left downto 0) <= d126_in;  h126_en <= en_in;
   h127_out(h127_out'left downto d127_in'left + 1) <= (others => '0');   h127_out(d127_in'left downto 0) <= d127_in;  h127_en <= en_in;
   h128_out(h128_out'left downto d128_in'left + 1) <= (others => '0');   h128_out(d128_in'left downto 0) <= d128_in;  h128_en <= en_in;
end generate g_Huff_enc_dis;  
                                                                                                  
Buf01 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 0), enw=>h01_en, data_in=>h01_out, data_out=>buff01_out, burst_r=>en_out( 0), fifo_empty=> open, fifo_full=> open ); 
Buf02 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 1), enw=>h02_en, data_in=>h02_out, data_out=>buff02_out, burst_r=>en_out( 1), fifo_empty=> open, fifo_full=> open ); 
Buf03 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 2), enw=>h03_en, data_in=>h03_out, data_out=>buff03_out, burst_r=>en_out( 2), fifo_empty=> open, fifo_full=> open ); 
Buf04 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 3), enw=>h04_en, data_in=>h04_out, data_out=>buff04_out, burst_r=>en_out( 3), fifo_empty=> open, fifo_full=> open ); 
Buf05 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 4), enw=>h05_en, data_in=>h05_out, data_out=>buff05_out, burst_r=>en_out( 4), fifo_empty=> open, fifo_full=> open ); 
Buf06 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 5), enw=>h06_en, data_in=>h06_out, data_out=>buff06_out, burst_r=>en_out( 5), fifo_empty=> open, fifo_full=> open ); 
Buf07 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 6), enw=>h07_en, data_in=>h07_out, data_out=>buff07_out, burst_r=>en_out( 6), fifo_empty=> open, fifo_full=> open ); 
Buf08 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 7), enw=>h08_en, data_in=>h08_out, data_out=>buff08_out, burst_r=>en_out( 7), fifo_empty=> open, fifo_full=> open ); 
Buf09 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 8), enw=>h09_en, data_in=>h09_out, data_out=>buff09_out, burst_r=>en_out( 8), fifo_empty=> open, fifo_full=> open ); 
Buf10 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 9), enw=>h10_en, data_in=>h10_out, data_out=>buff10_out, burst_r=>en_out( 9), fifo_empty=> open, fifo_full=> open ); 
Buf11 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(10), enw=>h11_en, data_in=>h11_out, data_out=>buff11_out, burst_r=>en_out(10), fifo_empty=> open, fifo_full=> open ); 
Buf12 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(11), enw=>h12_en, data_in=>h12_out, data_out=>buff12_out, burst_r=>en_out(11), fifo_empty=> open, fifo_full=> open ); 
Buf13 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(12), enw=>h13_en, data_in=>h13_out, data_out=>buff13_out, burst_r=>en_out(12), fifo_empty=> open, fifo_full=> open ); 
Buf14 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(13), enw=>h14_en, data_in=>h14_out, data_out=>buff14_out, burst_r=>en_out(13), fifo_empty=> open, fifo_full=> open ); 
Buf15 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(14), enw=>h15_en, data_in=>h15_out, data_out=>buff15_out, burst_r=>en_out(14), fifo_empty=> open, fifo_full=> open ); 
Buf16 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(15), enw=>h16_en, data_in=>h16_out, data_out=>buff16_out, burst_r=>en_out(15), fifo_empty=> open, fifo_full=> open ); 
Buf17 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(16), enw=>h17_en, data_in=>h17_out, data_out=>buff17_out, burst_r=>en_out(16), fifo_empty=> open, fifo_full=> open ); 
Buf18 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(17), enw=>h18_en, data_in=>h18_out, data_out=>buff18_out, burst_r=>en_out(17), fifo_empty=> open, fifo_full=> open ); 
Buf19 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(18), enw=>h19_en, data_in=>h19_out, data_out=>buff19_out, burst_r=>en_out(18), fifo_empty=> open, fifo_full=> open ); 
Buf20 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(19), enw=>h20_en, data_in=>h20_out, data_out=>buff20_out, burst_r=>en_out(19), fifo_empty=> open, fifo_full=> open ); 
Buf21 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(20), enw=>h21_en, data_in=>h21_out, data_out=>buff21_out, burst_r=>en_out(20), fifo_empty=> open, fifo_full=> open ); 
Buf22 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(21), enw=>h22_en, data_in=>h22_out, data_out=>buff22_out, burst_r=>en_out(21), fifo_empty=> open, fifo_full=> open ); 
Buf23 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(22), enw=>h23_en, data_in=>h23_out, data_out=>buff23_out, burst_r=>en_out(22), fifo_empty=> open, fifo_full=> open ); 
Buf24 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(23), enw=>h24_en, data_in=>h24_out, data_out=>buff24_out, burst_r=>en_out(23), fifo_empty=> open, fifo_full=> open ); 
Buf25 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(24), enw=>h25_en, data_in=>h25_out, data_out=>buff25_out, burst_r=>en_out(24), fifo_empty=> open, fifo_full=> open ); 
Buf26 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(25), enw=>h26_en, data_in=>h26_out, data_out=>buff26_out, burst_r=>en_out(25), fifo_empty=> open, fifo_full=> open ); 
Buf27 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(26), enw=>h27_en, data_in=>h27_out, data_out=>buff27_out, burst_r=>en_out(26), fifo_empty=> open, fifo_full=> open ); 
Buf28 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(27), enw=>h28_en, data_in=>h28_out, data_out=>buff28_out, burst_r=>en_out(27), fifo_empty=> open, fifo_full=> open ); 
Buf29 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(28), enw=>h29_en, data_in=>h29_out, data_out=>buff29_out, burst_r=>en_out(28), fifo_empty=> open, fifo_full=> open ); 
Buf30 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(29), enw=>h30_en, data_in=>h30_out, data_out=>buff30_out, burst_r=>en_out(29), fifo_empty=> open, fifo_full=> open ); 
Buf31 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(30), enw=>h31_en, data_in=>h31_out, data_out=>buff31_out, burst_r=>en_out(30), fifo_empty=> open, fifo_full=> open ); 
Buf32 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(31), enw=>h32_en, data_in=>h32_out, data_out=>buff32_out, burst_r=>en_out(31), fifo_empty=> open, fifo_full=> open ); 
Buf33 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(32), enw=>h33_en, data_in=>h33_out, data_out=>buff33_out, burst_r=>en_out(32), fifo_empty=> open, fifo_full=> open ); 
Buf34 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(33), enw=>h34_en, data_in=>h34_out, data_out=>buff34_out, burst_r=>en_out(33), fifo_empty=> open, fifo_full=> open ); 
Buf35 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(34), enw=>h35_en, data_in=>h35_out, data_out=>buff35_out, burst_r=>en_out(34), fifo_empty=> open, fifo_full=> open ); 
Buf36 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(35), enw=>h36_en, data_in=>h36_out, data_out=>buff36_out, burst_r=>en_out(35), fifo_empty=> open, fifo_full=> open ); 
Buf37 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(36), enw=>h37_en, data_in=>h37_out, data_out=>buff37_out, burst_r=>en_out(36), fifo_empty=> open, fifo_full=> open ); 
Buf38 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(37), enw=>h38_en, data_in=>h38_out, data_out=>buff38_out, burst_r=>en_out(37), fifo_empty=> open, fifo_full=> open ); 
Buf39 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(38), enw=>h39_en, data_in=>h39_out, data_out=>buff39_out, burst_r=>en_out(38), fifo_empty=> open, fifo_full=> open ); 
Buf40 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(39), enw=>h40_en, data_in=>h40_out, data_out=>buff40_out, burst_r=>en_out(39), fifo_empty=> open, fifo_full=> open ); 
Buf41 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(40), enw=>h41_en, data_in=>h41_out, data_out=>buff41_out, burst_r=>en_out(40), fifo_empty=> open, fifo_full=> open ); 
Buf42 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(41), enw=>h42_en, data_in=>h42_out, data_out=>buff42_out, burst_r=>en_out(41), fifo_empty=> open, fifo_full=> open ); 
Buf43 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(42), enw=>h43_en, data_in=>h43_out, data_out=>buff43_out, burst_r=>en_out(42), fifo_empty=> open, fifo_full=> open ); 
Buf44 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(43), enw=>h44_en, data_in=>h44_out, data_out=>buff44_out, burst_r=>en_out(43), fifo_empty=> open, fifo_full=> open ); 
Buf45 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(44), enw=>h45_en, data_in=>h45_out, data_out=>buff45_out, burst_r=>en_out(44), fifo_empty=> open, fifo_full=> open ); 
Buf46 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(45), enw=>h46_en, data_in=>h46_out, data_out=>buff46_out, burst_r=>en_out(45), fifo_empty=> open, fifo_full=> open ); 
Buf47 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(46), enw=>h47_en, data_in=>h47_out, data_out=>buff47_out, burst_r=>en_out(46), fifo_empty=> open, fifo_full=> open ); 
Buf48 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(47), enw=>h48_en, data_in=>h48_out, data_out=>buff48_out, burst_r=>en_out(47), fifo_empty=> open, fifo_full=> open ); 
Buf49 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(48), enw=>h49_en, data_in=>h49_out, data_out=>buff49_out, burst_r=>en_out(48), fifo_empty=> open, fifo_full=> open ); 
Buf50 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(49), enw=>h50_en, data_in=>h50_out, data_out=>buff50_out, burst_r=>en_out(49), fifo_empty=> open, fifo_full=> open ); 
Buf51 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(50), enw=>h51_en, data_in=>h51_out, data_out=>buff51_out, burst_r=>en_out(50), fifo_empty=> open, fifo_full=> open ); 
Buf52 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(51), enw=>h52_en, data_in=>h52_out, data_out=>buff52_out, burst_r=>en_out(51), fifo_empty=> open, fifo_full=> open ); 
Buf53 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(52), enw=>h53_en, data_in=>h53_out, data_out=>buff53_out, burst_r=>en_out(52), fifo_empty=> open, fifo_full=> open ); 
Buf54 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(53), enw=>h54_en, data_in=>h54_out, data_out=>buff54_out, burst_r=>en_out(53), fifo_empty=> open, fifo_full=> open ); 
Buf55 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(54), enw=>h55_en, data_in=>h55_out, data_out=>buff55_out, burst_r=>en_out(54), fifo_empty=> open, fifo_full=> open ); 
Buf56 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(55), enw=>h56_en, data_in=>h56_out, data_out=>buff56_out, burst_r=>en_out(55), fifo_empty=> open, fifo_full=> open ); 
Buf57 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(56), enw=>h57_en, data_in=>h57_out, data_out=>buff57_out, burst_r=>en_out(56), fifo_empty=> open, fifo_full=> open ); 
Buf58 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(57), enw=>h58_en, data_in=>h58_out, data_out=>buff58_out, burst_r=>en_out(57), fifo_empty=> open, fifo_full=> open ); 
Buf59 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(58), enw=>h59_en, data_in=>h59_out, data_out=>buff59_out, burst_r=>en_out(58), fifo_empty=> open, fifo_full=> open ); 
Buf60 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(59), enw=>h60_en, data_in=>h60_out, data_out=>buff60_out, burst_r=>en_out(59), fifo_empty=> open, fifo_full=> open ); 
Buf61 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(60), enw=>h61_en, data_in=>h61_out, data_out=>buff61_out, burst_r=>en_out(60), fifo_empty=> open, fifo_full=> open ); 
Buf62 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(61), enw=>h62_en, data_in=>h62_out, data_out=>buff62_out, burst_r=>en_out(61), fifo_empty=> open, fifo_full=> open ); 
Buf63 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(62), enw=>h63_en, data_in=>h63_out, data_out=>buff63_out, burst_r=>en_out(62), fifo_empty=> open, fifo_full=> open ); 
Buf64 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(63), enw=>h64_en, data_in=>h64_out, data_out=>buff64_out, burst_r=>en_out(63), fifo_empty=> open, fifo_full=> open ); 

Buf65  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 64), enw=>h65_en , data_in=>h65_out , data_out=>buff65_out , burst_r=>en_out( 64), fifo_empty=> open, fifo_full=> open ); 
Buf66  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 65), enw=>h66_en , data_in=>h66_out , data_out=>buff66_out , burst_r=>en_out( 65), fifo_empty=> open, fifo_full=> open ); 
Buf67  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 66), enw=>h67_en , data_in=>h67_out , data_out=>buff67_out , burst_r=>en_out( 66), fifo_empty=> open, fifo_full=> open ); 
Buf68  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 67), enw=>h68_en , data_in=>h68_out , data_out=>buff68_out , burst_r=>en_out( 67), fifo_empty=> open, fifo_full=> open ); 
Buf69  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 68), enw=>h69_en , data_in=>h69_out , data_out=>buff69_out , burst_r=>en_out( 68), fifo_empty=> open, fifo_full=> open ); 
Buf70  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 69), enw=>h70_en , data_in=>h70_out , data_out=>buff70_out , burst_r=>en_out( 69), fifo_empty=> open, fifo_full=> open ); 
Buf71  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 70), enw=>h71_en , data_in=>h71_out , data_out=>buff71_out , burst_r=>en_out( 70), fifo_empty=> open, fifo_full=> open ); 
Buf72  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 71), enw=>h72_en , data_in=>h72_out , data_out=>buff72_out , burst_r=>en_out( 71), fifo_empty=> open, fifo_full=> open ); 
Buf73  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 72), enw=>h73_en , data_in=>h73_out , data_out=>buff73_out , burst_r=>en_out( 72), fifo_empty=> open, fifo_full=> open ); 
Buf74  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 73), enw=>h74_en , data_in=>h74_out , data_out=>buff74_out , burst_r=>en_out( 73), fifo_empty=> open, fifo_full=> open ); 
Buf75  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 74), enw=>h75_en , data_in=>h75_out , data_out=>buff75_out , burst_r=>en_out( 74), fifo_empty=> open, fifo_full=> open ); 
Buf76  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 75), enw=>h76_en , data_in=>h76_out , data_out=>buff76_out , burst_r=>en_out( 75), fifo_empty=> open, fifo_full=> open ); 
Buf77  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 76), enw=>h77_en , data_in=>h77_out , data_out=>buff77_out , burst_r=>en_out( 76), fifo_empty=> open, fifo_full=> open ); 
Buf78  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 77), enw=>h78_en , data_in=>h78_out , data_out=>buff78_out , burst_r=>en_out( 77), fifo_empty=> open, fifo_full=> open ); 
Buf79  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 78), enw=>h79_en , data_in=>h79_out , data_out=>buff79_out , burst_r=>en_out( 78), fifo_empty=> open, fifo_full=> open ); 
Buf80  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 79), enw=>h80_en , data_in=>h80_out , data_out=>buff80_out , burst_r=>en_out( 79), fifo_empty=> open, fifo_full=> open ); 
Buf81  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 80), enw=>h81_en , data_in=>h81_out , data_out=>buff81_out , burst_r=>en_out( 80), fifo_empty=> open, fifo_full=> open ); 
Buf82  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 81), enw=>h82_en , data_in=>h82_out , data_out=>buff82_out , burst_r=>en_out( 81), fifo_empty=> open, fifo_full=> open ); 
Buf83  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 82), enw=>h83_en , data_in=>h83_out , data_out=>buff83_out , burst_r=>en_out( 82), fifo_empty=> open, fifo_full=> open ); 
Buf84  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 83), enw=>h84_en , data_in=>h84_out , data_out=>buff84_out , burst_r=>en_out( 83), fifo_empty=> open, fifo_full=> open ); 
Buf85  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 84), enw=>h85_en , data_in=>h85_out , data_out=>buff85_out , burst_r=>en_out( 84), fifo_empty=> open, fifo_full=> open ); 
Buf86  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 85), enw=>h86_en , data_in=>h86_out , data_out=>buff86_out , burst_r=>en_out( 85), fifo_empty=> open, fifo_full=> open ); 
Buf87  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 86), enw=>h87_en , data_in=>h87_out , data_out=>buff87_out , burst_r=>en_out( 86), fifo_empty=> open, fifo_full=> open ); 
Buf88  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 87), enw=>h88_en , data_in=>h88_out , data_out=>buff88_out , burst_r=>en_out( 87), fifo_empty=> open, fifo_full=> open ); 
Buf89  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 88), enw=>h89_en , data_in=>h89_out , data_out=>buff89_out , burst_r=>en_out( 88), fifo_empty=> open, fifo_full=> open ); 
Buf90  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 89), enw=>h90_en , data_in=>h90_out , data_out=>buff90_out , burst_r=>en_out( 89), fifo_empty=> open, fifo_full=> open ); 
Buf91  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 90), enw=>h91_en , data_in=>h91_out , data_out=>buff91_out , burst_r=>en_out( 90), fifo_empty=> open, fifo_full=> open ); 
Buf92  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 91), enw=>h92_en , data_in=>h92_out , data_out=>buff92_out , burst_r=>en_out( 91), fifo_empty=> open, fifo_full=> open ); 
Buf93  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 92), enw=>h93_en , data_in=>h93_out , data_out=>buff93_out , burst_r=>en_out( 92), fifo_empty=> open, fifo_full=> open ); 
Buf94  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 93), enw=>h94_en , data_in=>h94_out , data_out=>buff94_out , burst_r=>en_out( 93), fifo_empty=> open, fifo_full=> open ); 
Buf95  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 94), enw=>h95_en , data_in=>h95_out , data_out=>buff95_out , burst_r=>en_out( 94), fifo_empty=> open, fifo_full=> open ); 
Buf96  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 95), enw=>h96_en , data_in=>h96_out , data_out=>buff96_out , burst_r=>en_out( 95), fifo_empty=> open, fifo_full=> open ); 
Buf97  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 96), enw=>h97_en , data_in=>h97_out , data_out=>buff97_out , burst_r=>en_out( 96), fifo_empty=> open, fifo_full=> open ); 
Buf98  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 97), enw=>h98_en , data_in=>h98_out , data_out=>buff98_out , burst_r=>en_out( 97), fifo_empty=> open, fifo_full=> open ); 
Buf99  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 98), enw=>h99_en , data_in=>h99_out , data_out=>buff99_out , burst_r=>en_out( 98), fifo_empty=> open, fifo_full=> open ); 
Buf100 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 99), enw=>h100_en, data_in=>h100_out, data_out=>buff100_out, burst_r=>en_out( 99), fifo_empty=> open, fifo_full=> open ); 
Buf101 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(100), enw=>h101_en, data_in=>h101_out, data_out=>buff101_out, burst_r=>en_out(100), fifo_empty=> open, fifo_full=> open ); 
Buf102 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(101), enw=>h102_en, data_in=>h102_out, data_out=>buff102_out, burst_r=>en_out(101), fifo_empty=> open, fifo_full=> open ); 
Buf103 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(102), enw=>h103_en, data_in=>h103_out, data_out=>buff103_out, burst_r=>en_out(102), fifo_empty=> open, fifo_full=> open ); 
Buf104 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(103), enw=>h104_en, data_in=>h104_out, data_out=>buff104_out, burst_r=>en_out(103), fifo_empty=> open, fifo_full=> open ); 
Buf105 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(104), enw=>h105_en, data_in=>h105_out, data_out=>buff105_out, burst_r=>en_out(104), fifo_empty=> open, fifo_full=> open ); 
Buf106 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(105), enw=>h106_en, data_in=>h106_out, data_out=>buff106_out, burst_r=>en_out(105), fifo_empty=> open, fifo_full=> open ); 
Buf107 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(106), enw=>h107_en, data_in=>h107_out, data_out=>buff107_out, burst_r=>en_out(106), fifo_empty=> open, fifo_full=> open ); 
Buf108 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(107), enw=>h108_en, data_in=>h108_out, data_out=>buff108_out, burst_r=>en_out(107), fifo_empty=> open, fifo_full=> open ); 
Buf109 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(108), enw=>h109_en, data_in=>h109_out, data_out=>buff109_out, burst_r=>en_out(108), fifo_empty=> open, fifo_full=> open ); 
Buf110 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(109), enw=>h110_en, data_in=>h110_out, data_out=>buff110_out, burst_r=>en_out(109), fifo_empty=> open, fifo_full=> open ); 
Buf111 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(110), enw=>h111_en, data_in=>h111_out, data_out=>buff111_out, burst_r=>en_out(110), fifo_empty=> open, fifo_full=> open ); 
Buf112 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(111), enw=>h112_en, data_in=>h112_out, data_out=>buff112_out, burst_r=>en_out(111), fifo_empty=> open, fifo_full=> open ); 
Buf113 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(112), enw=>h113_en, data_in=>h113_out, data_out=>buff113_out, burst_r=>en_out(112), fifo_empty=> open, fifo_full=> open ); 
Buf114 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(113), enw=>h114_en, data_in=>h114_out, data_out=>buff114_out, burst_r=>en_out(113), fifo_empty=> open, fifo_full=> open ); 
Buf115 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(114), enw=>h115_en, data_in=>h115_out, data_out=>buff115_out, burst_r=>en_out(114), fifo_empty=> open, fifo_full=> open ); 
Buf116 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(115), enw=>h116_en, data_in=>h116_out, data_out=>buff116_out, burst_r=>en_out(115), fifo_empty=> open, fifo_full=> open ); 
Buf117 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(116), enw=>h117_en, data_in=>h117_out, data_out=>buff117_out, burst_r=>en_out(116), fifo_empty=> open, fifo_full=> open ); 
Buf118 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(117), enw=>h118_en, data_in=>h118_out, data_out=>buff118_out, burst_r=>en_out(117), fifo_empty=> open, fifo_full=> open ); 
Buf119 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(118), enw=>h119_en, data_in=>h119_out, data_out=>buff119_out, burst_r=>en_out(118), fifo_empty=> open, fifo_full=> open ); 
Buf120 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(119), enw=>h120_en, data_in=>h120_out, data_out=>buff120_out, burst_r=>en_out(119), fifo_empty=> open, fifo_full=> open ); 
Buf121 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(120), enw=>h121_en, data_in=>h121_out, data_out=>buff121_out, burst_r=>en_out(120), fifo_empty=> open, fifo_full=> open ); 
Buf122 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(121), enw=>h122_en, data_in=>h122_out, data_out=>buff122_out, burst_r=>en_out(121), fifo_empty=> open, fifo_full=> open ); 
Buf123 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(122), enw=>h123_en, data_in=>h123_out, data_out=>buff123_out, burst_r=>en_out(122), fifo_empty=> open, fifo_full=> open ); 
Buf124 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(123), enw=>h124_en, data_in=>h124_out, data_out=>buff124_out, burst_r=>en_out(123), fifo_empty=> open, fifo_full=> open ); 
Buf125 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(124), enw=>h125_en, data_in=>h125_out, data_out=>buff125_out, burst_r=>en_out(124), fifo_empty=> open, fifo_full=> open ); 
Buf126 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(125), enw=>h126_en, data_in=>h126_out, data_out=>buff126_out, burst_r=>en_out(125), fifo_empty=> open, fifo_full=> open ); 
Buf127 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(126), enw=>h127_en, data_in=>h127_out, data_out=>buff127_out, burst_r=>en_out(126), fifo_empty=> open, fifo_full=> open ); 
Buf128 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(127), enw=>h128_en, data_in=>h128_out, data_out=>buff128_out, burst_r=>en_out(127), fifo_empty=> open, fifo_full=> open ); 

--b_rd <= x"0000000000000001"; -- one Huffman
--d_out <= buff01_out;         -- one Huffman
p_rd_ctr :     process (clk, rst)
begin
   if ( rst = '1') then
      b_rd <= conv_std_logic_vector(0, b_rd'length);
   elsif(rising_edge(clk)) then   
      if buf_rd = '1' then
         --case
         if conv_integer('0' & buf_num) =    0 then b_rd <= x"00000000000000000000000000000001"; end if;
         if conv_integer('0' & buf_num) =    1 then b_rd <= x"00000000000000000000000000000002"; end if;
         if conv_integer('0' & buf_num) =    2 then b_rd <= x"00000000000000000000000000000004"; end if;
         if conv_integer('0' & buf_num) =    3 then b_rd <= x"00000000000000000000000000000008"; end if;
         if conv_integer('0' & buf_num) =    4 then b_rd <= x"00000000000000000000000000000010"; end if;
         if conv_integer('0' & buf_num) =    5 then b_rd <= x"00000000000000000000000000000020"; end if;
         if conv_integer('0' & buf_num) =    6 then b_rd <= x"00000000000000000000000000000040"; end if;
         if conv_integer('0' & buf_num) =    7 then b_rd <= x"00000000000000000000000000000080"; end if;
         if conv_integer('0' & buf_num) =    8 then b_rd <= x"00000000000000000000000000000100"; end if;
         if conv_integer('0' & buf_num) =    9 then b_rd <= x"00000000000000000000000000000200"; end if;
         if conv_integer('0' & buf_num) =   10 then b_rd <= x"00000000000000000000000000000400"; end if;
         if conv_integer('0' & buf_num) =   11 then b_rd <= x"00000000000000000000000000000800"; end if;
         if conv_integer('0' & buf_num) =   12 then b_rd <= x"00000000000000000000000000001000"; end if;
         if conv_integer('0' & buf_num) =   13 then b_rd <= x"00000000000000000000000000002000"; end if;
         if conv_integer('0' & buf_num) =   14 then b_rd <= x"00000000000000000000000000004000"; end if;
         if conv_integer('0' & buf_num) =   15 then b_rd <= x"00000000000000000000000000008000"; end if;
         if conv_integer('0' & buf_num) =   16 then b_rd <= x"00000000000000000000000000010000"; end if;
         if conv_integer('0' & buf_num) =   17 then b_rd <= x"00000000000000000000000000020000"; end if;
         if conv_integer('0' & buf_num) =   18 then b_rd <= x"00000000000000000000000000040000"; end if;
         if conv_integer('0' & buf_num) =   19 then b_rd <= x"00000000000000000000000000080000"; end if;
         if conv_integer('0' & buf_num) =   20 then b_rd <= x"00000000000000000000000000100000"; end if;
         if conv_integer('0' & buf_num) =   21 then b_rd <= x"00000000000000000000000000200000"; end if;
         if conv_integer('0' & buf_num) =   22 then b_rd <= x"00000000000000000000000000400000"; end if;
         if conv_integer('0' & buf_num) =   23 then b_rd <= x"00000000000000000000000000800000"; end if;
         if conv_integer('0' & buf_num) =   24 then b_rd <= x"00000000000000000000000001000000"; end if;
         if conv_integer('0' & buf_num) =   25 then b_rd <= x"00000000000000000000000002000000"; end if;
         if conv_integer('0' & buf_num) =   26 then b_rd <= x"00000000000000000000000004000000"; end if;
         if conv_integer('0' & buf_num) =   27 then b_rd <= x"00000000000000000000000008000000"; end if;
         if conv_integer('0' & buf_num) =   28 then b_rd <= x"00000000000000000000000010000000"; end if;
         if conv_integer('0' & buf_num) =   29 then b_rd <= x"00000000000000000000000020000000"; end if;
         if conv_integer('0' & buf_num) =   30 then b_rd <= x"00000000000000000000000040000000"; end if;
         if conv_integer('0' & buf_num) =   31 then b_rd <= x"00000000000000000000000080000000"; end if;
         if conv_integer('0' & buf_num) =   32 then b_rd <= x"00000000000000000000000100000000"; end if;
         if conv_integer('0' & buf_num) =   33 then b_rd <= x"00000000000000000000000200000000"; end if;
         if conv_integer('0' & buf_num) =   34 then b_rd <= x"00000000000000000000000400000000"; end if;
         if conv_integer('0' & buf_num) =   35 then b_rd <= x"00000000000000000000000800000000"; end if;
         if conv_integer('0' & buf_num) =   36 then b_rd <= x"00000000000000000000001000000000"; end if;
         if conv_integer('0' & buf_num) =   37 then b_rd <= x"00000000000000000000002000000000"; end if;
         if conv_integer('0' & buf_num) =   38 then b_rd <= x"00000000000000000000004000000000"; end if;
         if conv_integer('0' & buf_num) =   39 then b_rd <= x"00000000000000000000008000000000"; end if;
         if conv_integer('0' & buf_num) =   40 then b_rd <= x"00000000000000000000010000000000"; end if;
         if conv_integer('0' & buf_num) =   41 then b_rd <= x"00000000000000000000020000000000"; end if;
         if conv_integer('0' & buf_num) =   42 then b_rd <= x"00000000000000000000040000000000"; end if;
         if conv_integer('0' & buf_num) =   43 then b_rd <= x"00000000000000000000080000000000"; end if;
         if conv_integer('0' & buf_num) =   44 then b_rd <= x"00000000000000000000100000000000"; end if;
         if conv_integer('0' & buf_num) =   45 then b_rd <= x"00000000000000000000200000000000"; end if;
         if conv_integer('0' & buf_num) =   46 then b_rd <= x"00000000000000000000400000000000"; end if;
         if conv_integer('0' & buf_num) =   47 then b_rd <= x"00000000000000000000800000000000"; end if;
         if conv_integer('0' & buf_num) =   48 then b_rd <= x"00000000000000000001000000000000"; end if;
         if conv_integer('0' & buf_num) =   49 then b_rd <= x"00000000000000000002000000000000"; end if;
         if conv_integer('0' & buf_num) =   50 then b_rd <= x"00000000000000000004000000000000"; end if;
         if conv_integer('0' & buf_num) =   51 then b_rd <= x"00000000000000000008000000000000"; end if;
         if conv_integer('0' & buf_num) =   52 then b_rd <= x"00000000000000000010000000000000"; end if;
         if conv_integer('0' & buf_num) =   53 then b_rd <= x"00000000000000000020000000000000"; end if;
         if conv_integer('0' & buf_num) =   54 then b_rd <= x"00000000000000000040000000000000"; end if;
         if conv_integer('0' & buf_num) =   55 then b_rd <= x"00000000000000000080000000000000"; end if;
         if conv_integer('0' & buf_num) =   56 then b_rd <= x"00000000000000000100000000000000"; end if;
         if conv_integer('0' & buf_num) =   57 then b_rd <= x"00000000000000000200000000000000"; end if;
         if conv_integer('0' & buf_num) =   58 then b_rd <= x"00000000000000000400000000000000"; end if;
         if conv_integer('0' & buf_num) =   59 then b_rd <= x"00000000000000000800000000000000"; end if;
         if conv_integer('0' & buf_num) =   60 then b_rd <= x"00000000000000001000000000000000"; end if;
         if conv_integer('0' & buf_num) =   61 then b_rd <= x"00000000000000002000000000000000"; end if;
         if conv_integer('0' & buf_num) =   62 then b_rd <= x"00000000000000004000000000000000"; end if;
         if conv_integer('0' & buf_num) =   63 then b_rd <= x"00000000000000008000000000000000"; end if;

         if conv_integer('0' & buf_num) =   65  then b_rd <= x"00000000000000010000000000000000"; end if;
         if conv_integer('0' & buf_num) =   66  then b_rd <= x"00000000000000020000000000000000"; end if;
         if conv_integer('0' & buf_num) =   67  then b_rd <= x"00000000000000040000000000000000"; end if;
         if conv_integer('0' & buf_num) =   68  then b_rd <= x"00000000000000080000000000000000"; end if;
         if conv_integer('0' & buf_num) =   69  then b_rd <= x"00000000000000100000000000000000"; end if;
         if conv_integer('0' & buf_num) =   70  then b_rd <= x"00000000000000200000000000000000"; end if;
         if conv_integer('0' & buf_num) =   71  then b_rd <= x"00000000000000400000000000000000"; end if;
         if conv_integer('0' & buf_num) =   72  then b_rd <= x"00000000000000800000000000000000"; end if;
         if conv_integer('0' & buf_num) =   73  then b_rd <= x"00000000000001000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   74  then b_rd <= x"00000000000002000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   75  then b_rd <= x"00000000000004000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   76  then b_rd <= x"00000000000008000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   77  then b_rd <= x"00000000000010000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   78  then b_rd <= x"00000000000020000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   79  then b_rd <= x"00000000000040000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   80  then b_rd <= x"00000000000080000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   81  then b_rd <= x"00000000000100000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   82  then b_rd <= x"00000000000200000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   83  then b_rd <= x"00000000000400000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   84  then b_rd <= x"00000000000800000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   85  then b_rd <= x"00000000001000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   86  then b_rd <= x"00000000002000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   87  then b_rd <= x"00000000004000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   88  then b_rd <= x"00000000008000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   89  then b_rd <= x"00000000010000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   90  then b_rd <= x"00000000020000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   91  then b_rd <= x"00000000040000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   92  then b_rd <= x"00000000080000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   93  then b_rd <= x"00000000100000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   94  then b_rd <= x"00000000200000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   95  then b_rd <= x"00000000400000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   96  then b_rd <= x"00000000800000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   97  then b_rd <= x"00000001000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   98  then b_rd <= x"00000002000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   99  then b_rd <= x"00000004000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  100  then b_rd <= x"00000008000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  101  then b_rd <= x"00000010000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  102  then b_rd <= x"00000020000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  103  then b_rd <= x"00000040000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  104  then b_rd <= x"00000080000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  105  then b_rd <= x"00000100000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  106  then b_rd <= x"00000200000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  107  then b_rd <= x"00000400000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  108  then b_rd <= x"00000800000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  109  then b_rd <= x"00001000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  110  then b_rd <= x"00002000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  111  then b_rd <= x"00004000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  112  then b_rd <= x"00008000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  113  then b_rd <= x"00010000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  114  then b_rd <= x"00020000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  115  then b_rd <= x"00040000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  116  then b_rd <= x"00080000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  117  then b_rd <= x"00100000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  118  then b_rd <= x"00200000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  119  then b_rd <= x"00400000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  120  then b_rd <= x"00800000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  121  then b_rd <= x"01000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  122  then b_rd <= x"02000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  123  then b_rd <= x"04000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  124  then b_rd <= x"08000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  125  then b_rd <= x"10000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  126  then b_rd <= x"20000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  127  then b_rd <= x"40000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  128  then b_rd <= x"80000000000000000000000000000000"; end if;
            --for i in 0 to (2**C_INPUT_SIZE)-1 generate
            ----begin
            --    when (i = conv_integer(buf_num)) => b_rd <= conv_std_logic_vector((i*2), b_rd'length);        
            --end generate;
            --when others => b_rd <= conv_std_logic_vector(0, b_rd'length);
         --end case;
      end if;
      if conv_integer('0' & buf_num) =  0 then d_out <= buff01_out; end if;
      if conv_integer('0' & buf_num) =  1 then d_out <= buff02_out; end if;
      if conv_integer('0' & buf_num) =  2 then d_out <= buff03_out; end if;
      if conv_integer('0' & buf_num) =  3 then d_out <= buff04_out; end if;
      if conv_integer('0' & buf_num) =  4 then d_out <= buff05_out; end if;
      if conv_integer('0' & buf_num) =  5 then d_out <= buff06_out; end if;
      if conv_integer('0' & buf_num) =  6 then d_out <= buff07_out; end if;
      if conv_integer('0' & buf_num) =  7 then d_out <= buff08_out; end if;
      if conv_integer('0' & buf_num) =  8 then d_out <= buff09_out; end if;
      if conv_integer('0' & buf_num) =  9 then d_out <= buff10_out; end if;
      if conv_integer('0' & buf_num) = 10 then d_out <= buff11_out; end if;
      if conv_integer('0' & buf_num) = 11 then d_out <= buff12_out; end if;
      if conv_integer('0' & buf_num) = 12 then d_out <= buff13_out; end if;
      if conv_integer('0' & buf_num) = 13 then d_out <= buff14_out; end if;
      if conv_integer('0' & buf_num) = 14 then d_out <= buff15_out; end if;
      if conv_integer('0' & buf_num) = 15 then d_out <= buff16_out; end if;
      if conv_integer('0' & buf_num) = 16 then d_out <= buff17_out; end if;
      if conv_integer('0' & buf_num) = 17 then d_out <= buff18_out; end if;
      if conv_integer('0' & buf_num) = 18 then d_out <= buff19_out; end if;
      if conv_integer('0' & buf_num) = 19 then d_out <= buff20_out; end if;
      if conv_integer('0' & buf_num) = 20 then d_out <= buff21_out; end if;
      if conv_integer('0' & buf_num) = 21 then d_out <= buff22_out; end if;
      if conv_integer('0' & buf_num) = 22 then d_out <= buff23_out; end if;
      if conv_integer('0' & buf_num) = 23 then d_out <= buff24_out; end if;
      if conv_integer('0' & buf_num) = 24 then d_out <= buff25_out; end if;
      if conv_integer('0' & buf_num) = 25 then d_out <= buff26_out; end if;
      if conv_integer('0' & buf_num) = 26 then d_out <= buff27_out; end if;
      if conv_integer('0' & buf_num) = 27 then d_out <= buff28_out; end if;
      if conv_integer('0' & buf_num) = 28 then d_out <= buff29_out; end if;
      if conv_integer('0' & buf_num) = 29 then d_out <= buff30_out; end if;
      if conv_integer('0' & buf_num) = 30 then d_out <= buff31_out; end if;
      if conv_integer('0' & buf_num) = 31 then d_out <= buff32_out; end if;
      if conv_integer('0' & buf_num) = 32 then d_out <= buff33_out; end if;
      if conv_integer('0' & buf_num) = 33 then d_out <= buff34_out; end if;
      if conv_integer('0' & buf_num) = 34 then d_out <= buff35_out; end if;
      if conv_integer('0' & buf_num) = 35 then d_out <= buff36_out; end if;
      if conv_integer('0' & buf_num) = 36 then d_out <= buff37_out; end if;
      if conv_integer('0' & buf_num) = 37 then d_out <= buff38_out; end if;
      if conv_integer('0' & buf_num) = 38 then d_out <= buff39_out; end if;
      if conv_integer('0' & buf_num) = 39 then d_out <= buff40_out; end if;
      if conv_integer('0' & buf_num) = 40 then d_out <= buff41_out; end if;
      if conv_integer('0' & buf_num) = 41 then d_out <= buff42_out; end if;
      if conv_integer('0' & buf_num) = 42 then d_out <= buff43_out; end if;
      if conv_integer('0' & buf_num) = 43 then d_out <= buff44_out; end if;
      if conv_integer('0' & buf_num) = 44 then d_out <= buff45_out; end if;
      if conv_integer('0' & buf_num) = 45 then d_out <= buff46_out; end if;
      if conv_integer('0' & buf_num) = 46 then d_out <= buff47_out; end if;
      if conv_integer('0' & buf_num) = 47 then d_out <= buff48_out; end if;
      if conv_integer('0' & buf_num) = 48 then d_out <= buff49_out; end if;
      if conv_integer('0' & buf_num) = 49 then d_out <= buff50_out; end if;
      if conv_integer('0' & buf_num) = 50 then d_out <= buff51_out; end if;
      if conv_integer('0' & buf_num) = 51 then d_out <= buff52_out; end if;
      if conv_integer('0' & buf_num) = 52 then d_out <= buff53_out; end if;
      if conv_integer('0' & buf_num) = 53 then d_out <= buff54_out; end if;
      if conv_integer('0' & buf_num) = 54 then d_out <= buff55_out; end if;
      if conv_integer('0' & buf_num) = 55 then d_out <= buff56_out; end if;
      if conv_integer('0' & buf_num) = 56 then d_out <= buff57_out; end if;
      if conv_integer('0' & buf_num) = 57 then d_out <= buff58_out; end if;
      if conv_integer('0' & buf_num) = 58 then d_out <= buff59_out; end if;
      if conv_integer('0' & buf_num) = 59 then d_out <= buff60_out; end if;
      if conv_integer('0' & buf_num) = 60 then d_out <= buff61_out; end if;
      if conv_integer('0' & buf_num) = 61 then d_out <= buff62_out; end if;
      if conv_integer('0' & buf_num) = 62 then d_out <= buff63_out; end if;
      if conv_integer('0' & buf_num) = 63 then d_out <= buff64_out; end if;

      if conv_integer('0' & buf_num) = 65  then d_out <= buff65_out ; end if;
      if conv_integer('0' & buf_num) = 66  then d_out <= buff66_out ; end if;
      if conv_integer('0' & buf_num) = 67  then d_out <= buff67_out ; end if;
      if conv_integer('0' & buf_num) = 68  then d_out <= buff68_out ; end if;
      if conv_integer('0' & buf_num) = 69  then d_out <= buff69_out ; end if;
      if conv_integer('0' & buf_num) = 70  then d_out <= buff70_out ; end if;
      if conv_integer('0' & buf_num) = 71  then d_out <= buff71_out ; end if;
      if conv_integer('0' & buf_num) = 72  then d_out <= buff72_out ; end if;
      if conv_integer('0' & buf_num) = 73  then d_out <= buff73_out ; end if;
      if conv_integer('0' & buf_num) = 74  then d_out <= buff74_out ; end if;
      if conv_integer('0' & buf_num) = 75  then d_out <= buff75_out ; end if;
      if conv_integer('0' & buf_num) = 76  then d_out <= buff76_out ; end if;
      if conv_integer('0' & buf_num) = 77  then d_out <= buff77_out ; end if;
      if conv_integer('0' & buf_num) = 78  then d_out <= buff78_out ; end if;
      if conv_integer('0' & buf_num) = 79  then d_out <= buff79_out ; end if;
      if conv_integer('0' & buf_num) = 80  then d_out <= buff80_out ; end if;
      if conv_integer('0' & buf_num) = 81  then d_out <= buff81_out ; end if;
      if conv_integer('0' & buf_num) = 82  then d_out <= buff82_out ; end if;
      if conv_integer('0' & buf_num) = 83  then d_out <= buff83_out ; end if;
      if conv_integer('0' & buf_num) = 84  then d_out <= buff84_out ; end if;
      if conv_integer('0' & buf_num) = 85  then d_out <= buff85_out ; end if;
      if conv_integer('0' & buf_num) = 86  then d_out <= buff86_out ; end if;
      if conv_integer('0' & buf_num) = 87  then d_out <= buff87_out ; end if;
      if conv_integer('0' & buf_num) = 88  then d_out <= buff88_out ; end if;
      if conv_integer('0' & buf_num) = 89  then d_out <= buff89_out ; end if;
      if conv_integer('0' & buf_num) = 90  then d_out <= buff90_out ; end if;
      if conv_integer('0' & buf_num) = 91  then d_out <= buff91_out ; end if;
      if conv_integer('0' & buf_num) = 92  then d_out <= buff92_out ; end if;
      if conv_integer('0' & buf_num) = 93  then d_out <= buff93_out ; end if;
      if conv_integer('0' & buf_num) = 94  then d_out <= buff94_out ; end if;
      if conv_integer('0' & buf_num) = 95  then d_out <= buff95_out ; end if;
      if conv_integer('0' & buf_num) = 96  then d_out <= buff96_out ; end if;
      if conv_integer('0' & buf_num) = 97  then d_out <= buff97_out ; end if;
      if conv_integer('0' & buf_num) = 98  then d_out <= buff98_out ; end if;
      if conv_integer('0' & buf_num) = 99  then d_out <= buff99_out ; end if;
      if conv_integer('0' & buf_num) =100  then d_out <= buff100_out; end if;
      if conv_integer('0' & buf_num) =101  then d_out <= buff101_out; end if;
      if conv_integer('0' & buf_num) =102  then d_out <= buff102_out; end if;
      if conv_integer('0' & buf_num) =103  then d_out <= buff103_out; end if;
      if conv_integer('0' & buf_num) =104  then d_out <= buff104_out; end if;
      if conv_integer('0' & buf_num) =105  then d_out <= buff105_out; end if;
      if conv_integer('0' & buf_num) =106  then d_out <= buff106_out; end if;
      if conv_integer('0' & buf_num) =107  then d_out <= buff107_out; end if;
      if conv_integer('0' & buf_num) =108  then d_out <= buff108_out; end if;
      if conv_integer('0' & buf_num) =109  then d_out <= buff109_out; end if;
      if conv_integer('0' & buf_num) =110  then d_out <= buff110_out; end if;
      if conv_integer('0' & buf_num) =111  then d_out <= buff111_out; end if;
      if conv_integer('0' & buf_num) =112  then d_out <= buff112_out; end if;
      if conv_integer('0' & buf_num) =113  then d_out <= buff113_out; end if;
      if conv_integer('0' & buf_num) =114  then d_out <= buff114_out; end if;
      if conv_integer('0' & buf_num) =115  then d_out <= buff115_out; end if;
      if conv_integer('0' & buf_num) =116  then d_out <= buff116_out; end if;
      if conv_integer('0' & buf_num) =117  then d_out <= buff117_out; end if;
      if conv_integer('0' & buf_num) =118  then d_out <= buff118_out; end if;
      if conv_integer('0' & buf_num) =119  then d_out <= buff119_out; end if;
      if conv_integer('0' & buf_num) =120  then d_out <= buff120_out; end if;
      if conv_integer('0' & buf_num) =121  then d_out <= buff121_out; end if;
      if conv_integer('0' & buf_num) =122  then d_out <= buff122_out; end if;
      if conv_integer('0' & buf_num) =123  then d_out <= buff123_out; end if;
      if conv_integer('0' & buf_num) =124  then d_out <= buff124_out; end if;
      if conv_integer('0' & buf_num) =125  then d_out <= buff125_out; end if;
      if conv_integer('0' & buf_num) =126  then d_out <= buff126_out; end if;
      if conv_integer('0' & buf_num) =127  then d_out <= buff127_out; end if;
      if conv_integer('0' & buf_num) =128  then d_out <= buff128_out; end if;
   end if;
end process p_rd_ctr;

end a;