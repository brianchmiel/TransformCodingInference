library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_SIGNED.ALL;

entity Huffman256 is
  generic (
           N             : integer := 4;  -- input data width
           M             : integer := 8;  -- max code width
           Wh            : integer := 16;  -- Huffman unit output data width (Note W>=M)
           Wb            : integer := 512; -- output buffer data width
           Huff_enc_en   : boolean := TRUE; -- Huffman encoder Enable/Bypass
           depth         : integer := 500; -- buffer depth
           burst         : integer := 10   -- buffer read burst
  	       );
  port    (
           clk           : in  std_logic;
           rst           : in  std_logic; 

           init_en       : in  std_logic;                         -- initialising convert table
           alpha_data    : in  std_logic_vector(N-1 downto 0);    
           alpha_code    : in  std_logic_vector(M-1 downto 0);    
           alpha_width   : in  std_logic_vector(  3 downto 0);

  	       d01_in, d65_in , d129_in, d193_in   : in std_logic_vector (N-1 downto 0);
           d02_in, d66_in , d130_in, d194_in   : in std_logic_vector (N-1 downto 0);
           d03_in, d67_in , d131_in, d195_in   : in std_logic_vector (N-1 downto 0);
           d04_in, d68_in , d132_in, d196_in   : in std_logic_vector (N-1 downto 0);
           d05_in, d69_in , d133_in, d197_in   : in std_logic_vector (N-1 downto 0);
           d06_in, d70_in , d134_in, d198_in   : in std_logic_vector (N-1 downto 0);
           d07_in, d71_in , d135_in, d199_in   : in std_logic_vector (N-1 downto 0);
           d08_in, d72_in , d136_in, d200_in   : in std_logic_vector (N-1 downto 0);
           d09_in, d73_in , d137_in, d201_in   : in std_logic_vector (N-1 downto 0);
           d10_in, d74_in , d138_in, d202_in   : in std_logic_vector (N-1 downto 0);
           d11_in, d75_in , d139_in, d203_in   : in std_logic_vector (N-1 downto 0);
           d12_in, d76_in , d140_in, d204_in   : in std_logic_vector (N-1 downto 0);
           d13_in, d77_in , d141_in, d205_in   : in std_logic_vector (N-1 downto 0);
           d14_in, d78_in , d142_in, d206_in   : in std_logic_vector (N-1 downto 0);
           d15_in, d79_in , d143_in, d207_in   : in std_logic_vector (N-1 downto 0);
           d16_in, d80_in , d144_in, d208_in   : in std_logic_vector (N-1 downto 0);
           d17_in, d81_in , d145_in, d209_in   : in std_logic_vector (N-1 downto 0);
           d18_in, d82_in , d146_in, d210_in   : in std_logic_vector (N-1 downto 0);
           d19_in, d83_in , d147_in, d211_in   : in std_logic_vector (N-1 downto 0);
           d20_in, d84_in , d148_in, d212_in   : in std_logic_vector (N-1 downto 0);
           d21_in, d85_in , d149_in, d213_in   : in std_logic_vector (N-1 downto 0);
           d22_in, d86_in , d150_in, d214_in   : in std_logic_vector (N-1 downto 0);
           d23_in, d87_in , d151_in, d215_in   : in std_logic_vector (N-1 downto 0);
           d24_in, d88_in , d152_in, d216_in   : in std_logic_vector (N-1 downto 0);
           d25_in, d89_in , d153_in, d217_in   : in std_logic_vector (N-1 downto 0);
           d26_in, d90_in , d154_in, d218_in   : in std_logic_vector (N-1 downto 0);
           d27_in, d91_in , d155_in, d219_in   : in std_logic_vector (N-1 downto 0);
           d28_in, d92_in , d156_in, d220_in   : in std_logic_vector (N-1 downto 0);
           d29_in, d93_in , d157_in, d221_in   : in std_logic_vector (N-1 downto 0);
           d30_in, d94_in , d158_in, d222_in   : in std_logic_vector (N-1 downto 0);
           d31_in, d95_in , d159_in, d223_in   : in std_logic_vector (N-1 downto 0);
           d32_in, d96_in , d160_in, d224_in   : in std_logic_vector (N-1 downto 0);
           d33_in, d97_in , d161_in, d225_in   : in std_logic_vector (N-1 downto 0);
           d34_in, d98_in , d162_in, d226_in   : in std_logic_vector (N-1 downto 0);
           d35_in, d99_in , d163_in, d227_in   : in std_logic_vector (N-1 downto 0);
           d36_in, d100_in, d164_in, d228_in   : in std_logic_vector (N-1 downto 0);
           d37_in, d101_in, d165_in, d229_in   : in std_logic_vector (N-1 downto 0);
           d38_in, d102_in, d166_in, d230_in   : in std_logic_vector (N-1 downto 0);
           d39_in, d103_in, d167_in, d231_in   : in std_logic_vector (N-1 downto 0);
           d40_in, d104_in, d168_in, d232_in   : in std_logic_vector (N-1 downto 0);
           d41_in, d105_in, d169_in, d233_in   : in std_logic_vector (N-1 downto 0);
           d42_in, d106_in, d170_in, d234_in   : in std_logic_vector (N-1 downto 0);
           d43_in, d107_in, d171_in, d235_in   : in std_logic_vector (N-1 downto 0);
           d44_in, d108_in, d172_in, d236_in   : in std_logic_vector (N-1 downto 0);
           d45_in, d109_in, d173_in, d237_in   : in std_logic_vector (N-1 downto 0);
           d46_in, d110_in, d174_in, d238_in   : in std_logic_vector (N-1 downto 0);
           d47_in, d111_in, d175_in, d239_in   : in std_logic_vector (N-1 downto 0);
           d48_in, d112_in, d176_in, d240_in   : in std_logic_vector (N-1 downto 0);
           d49_in, d113_in, d177_in, d241_in   : in std_logic_vector (N-1 downto 0);
           d50_in, d114_in, d178_in, d242_in   : in std_logic_vector (N-1 downto 0);
           d51_in, d115_in, d179_in, d243_in   : in std_logic_vector (N-1 downto 0);
           d52_in, d116_in, d180_in, d244_in   : in std_logic_vector (N-1 downto 0);
           d53_in, d117_in, d181_in, d245_in   : in std_logic_vector (N-1 downto 0);
           d54_in, d118_in, d182_in, d246_in   : in std_logic_vector (N-1 downto 0);
           d55_in, d119_in, d183_in, d247_in   : in std_logic_vector (N-1 downto 0);
           d56_in, d120_in, d184_in, d248_in   : in std_logic_vector (N-1 downto 0);
           d57_in, d121_in, d185_in, d249_in   : in std_logic_vector (N-1 downto 0);
           d58_in, d122_in, d186_in, d250_in   : in std_logic_vector (N-1 downto 0);
           d59_in, d123_in, d187_in, d251_in   : in std_logic_vector (N-1 downto 0);
           d60_in, d124_in, d188_in, d252_in   : in std_logic_vector (N-1 downto 0);
           d61_in, d125_in, d189_in, d253_in   : in std_logic_vector (N-1 downto 0);
           d62_in, d126_in, d190_in, d254_in   : in std_logic_vector (N-1 downto 0);
           d63_in, d127_in, d191_in, d255_in   : in std_logic_vector (N-1 downto 0);
           d64_in, d128_in, d192_in, d256_in   : in std_logic_vector (N-1 downto 0);

  	       en_in         : in  std_logic;
  	       sof_in        : in  std_logic;                         -- start of frame
           eof_in        : in  std_logic;                         -- end of frame

           buf_rd        : in  std_logic;
           buf_num       : in  std_logic_vector (7      downto 0);
           d_out         : out std_logic_vector (Wb  -1 downto 0);
           en_out        : out std_logic_vector (256  -1 downto 0);
           eof_out       : out std_logic);                        -- huffman code output
end Huffman256;

architecture a of Huffman256 is


component Huffman is
  generic (
           N             : integer := 4; -- input data width
           M             : integer := 8; -- max code width
           W             : integer := 10 -- output data width (Note W>=M)
           );
  port    (
           clk           : in  std_logic;
           rst           : in  std_logic; 

           init_en       : in  std_logic;                         -- initialising convert table
           alpha_data    : in  std_logic_vector(N-1 downto 0);    
           alpha_code    : in  std_logic_vector(M-1 downto 0);    
           alpha_width   : in  std_logic_vector(  3 downto 0);

           d_in          : in  std_logic_vector (N-1 downto 0);   -- data to convert
           en_in         : in  std_logic;
           sof_in        : in  std_logic;                         -- start of frame
           eof_in        : in  std_logic;                         -- end of frame

           d_out         : out std_logic_vector (W-1 downto 0);
           en_out        : out std_logic;
           eof_out       : out std_logic);                        -- huffman codde output
end component;

component fifo is
generic (depth   : integer := 16 ;
         burst   : integer := 10 ;  -- indication for burst read (Note, depth>burst) 
         Win     : integer := 16 ;
         Wout    : integer := 64 );  --depth of fifo
port (    clk        : in std_logic;
          rst        : in std_logic;
          enr        : in std_logic;   --enable read,should be '0' when not in use.
          enw        : in std_logic;    --enable write,should be '0' when not in use.
          data_in    : in std_logic_vector  (Win -1 downto 0);     --input data
          data_out   : out std_logic_vector(Wout-1 downto 0);    --output data
          burst_r    : out std_logic;   --set as '1' when the queue is ready for burst transaction
          fifo_empty : out std_logic;   --set as '1' when the queue is empty
          fifo_full  : out std_logic     --set as '1' when the queue is full
         );
end component;

signal h01_out, h65_out , h129_out, h193_out    : std_logic_vector(Wh-1 downto 0);
signal h02_out, h66_out , h130_out, h194_out    : std_logic_vector(Wh-1 downto 0);
signal h03_out, h67_out , h131_out, h195_out    : std_logic_vector(Wh-1 downto 0);
signal h04_out, h68_out , h132_out, h196_out    : std_logic_vector(Wh-1 downto 0);
signal h05_out, h69_out , h133_out, h197_out    : std_logic_vector(Wh-1 downto 0);
signal h06_out, h70_out , h134_out, h198_out    : std_logic_vector(Wh-1 downto 0);
signal h07_out, h71_out , h135_out, h199_out    : std_logic_vector(Wh-1 downto 0);
signal h08_out, h72_out , h136_out, h200_out    : std_logic_vector(Wh-1 downto 0);
signal h09_out, h73_out , h137_out, h201_out    : std_logic_vector(Wh-1 downto 0);
signal h10_out, h74_out , h138_out, h202_out    : std_logic_vector(Wh-1 downto 0);
signal h11_out, h75_out , h139_out, h203_out    : std_logic_vector(Wh-1 downto 0);
signal h12_out, h76_out , h140_out, h204_out    : std_logic_vector(Wh-1 downto 0);
signal h13_out, h77_out , h141_out, h205_out    : std_logic_vector(Wh-1 downto 0);
signal h14_out, h78_out , h142_out, h206_out    : std_logic_vector(Wh-1 downto 0);
signal h15_out, h79_out , h143_out, h207_out    : std_logic_vector(Wh-1 downto 0);
signal h16_out, h80_out , h144_out, h208_out    : std_logic_vector(Wh-1 downto 0);
signal h17_out, h81_out , h145_out, h209_out    : std_logic_vector(Wh-1 downto 0);
signal h18_out, h82_out , h146_out, h210_out    : std_logic_vector(Wh-1 downto 0);
signal h19_out, h83_out , h147_out, h211_out    : std_logic_vector(Wh-1 downto 0);
signal h20_out, h84_out , h148_out, h212_out    : std_logic_vector(Wh-1 downto 0);
signal h21_out, h85_out , h149_out, h213_out    : std_logic_vector(Wh-1 downto 0);
signal h22_out, h86_out , h150_out, h214_out    : std_logic_vector(Wh-1 downto 0);
signal h23_out, h87_out , h151_out, h215_out    : std_logic_vector(Wh-1 downto 0);
signal h24_out, h88_out , h152_out, h216_out    : std_logic_vector(Wh-1 downto 0);
signal h25_out, h89_out , h153_out, h217_out    : std_logic_vector(Wh-1 downto 0);
signal h26_out, h90_out , h154_out, h218_out    : std_logic_vector(Wh-1 downto 0);
signal h27_out, h91_out , h155_out, h219_out    : std_logic_vector(Wh-1 downto 0);
signal h28_out, h92_out , h156_out, h220_out    : std_logic_vector(Wh-1 downto 0);
signal h29_out, h93_out , h157_out, h221_out    : std_logic_vector(Wh-1 downto 0);
signal h30_out, h94_out , h158_out, h222_out    : std_logic_vector(Wh-1 downto 0);
signal h31_out, h95_out , h159_out, h223_out    : std_logic_vector(Wh-1 downto 0);
signal h32_out, h96_out , h160_out, h224_out    : std_logic_vector(Wh-1 downto 0);
signal h33_out, h97_out , h161_out, h225_out    : std_logic_vector(Wh-1 downto 0);
signal h34_out, h98_out , h162_out, h226_out    : std_logic_vector(Wh-1 downto 0);
signal h35_out, h99_out , h163_out, h227_out    : std_logic_vector(Wh-1 downto 0);
signal h36_out, h100_out, h164_out, h228_out    : std_logic_vector(Wh-1 downto 0);
signal h37_out, h101_out, h165_out, h229_out    : std_logic_vector(Wh-1 downto 0);
signal h38_out, h102_out, h166_out, h230_out    : std_logic_vector(Wh-1 downto 0);
signal h39_out, h103_out, h167_out, h231_out    : std_logic_vector(Wh-1 downto 0);
signal h40_out, h104_out, h168_out, h232_out    : std_logic_vector(Wh-1 downto 0);
signal h41_out, h105_out, h169_out, h233_out    : std_logic_vector(Wh-1 downto 0);
signal h42_out, h106_out, h170_out, h234_out    : std_logic_vector(Wh-1 downto 0);
signal h43_out, h107_out, h171_out, h235_out    : std_logic_vector(Wh-1 downto 0);
signal h44_out, h108_out, h172_out, h236_out    : std_logic_vector(Wh-1 downto 0);
signal h45_out, h109_out, h173_out, h237_out    : std_logic_vector(Wh-1 downto 0);
signal h46_out, h110_out, h174_out, h238_out    : std_logic_vector(Wh-1 downto 0);
signal h47_out, h111_out, h175_out, h239_out    : std_logic_vector(Wh-1 downto 0);
signal h48_out, h112_out, h176_out, h240_out    : std_logic_vector(Wh-1 downto 0);
signal h49_out, h113_out, h177_out, h241_out    : std_logic_vector(Wh-1 downto 0);
signal h50_out, h114_out, h178_out, h242_out    : std_logic_vector(Wh-1 downto 0);
signal h51_out, h115_out, h179_out, h243_out    : std_logic_vector(Wh-1 downto 0);
signal h52_out, h116_out, h180_out, h244_out    : std_logic_vector(Wh-1 downto 0);
signal h53_out, h117_out, h181_out, h245_out    : std_logic_vector(Wh-1 downto 0);
signal h54_out, h118_out, h182_out, h246_out    : std_logic_vector(Wh-1 downto 0);
signal h55_out, h119_out, h183_out, h247_out    : std_logic_vector(Wh-1 downto 0);
signal h56_out, h120_out, h184_out, h248_out    : std_logic_vector(Wh-1 downto 0);
signal h57_out, h121_out, h185_out, h249_out    : std_logic_vector(Wh-1 downto 0);
signal h58_out, h122_out, h186_out, h250_out    : std_logic_vector(Wh-1 downto 0);
signal h59_out, h123_out, h187_out, h251_out    : std_logic_vector(Wh-1 downto 0);
signal h60_out, h124_out, h188_out, h252_out    : std_logic_vector(Wh-1 downto 0);
signal h61_out, h125_out, h189_out, h253_out    : std_logic_vector(Wh-1 downto 0);
signal h62_out, h126_out, h190_out, h254_out    : std_logic_vector(Wh-1 downto 0);
signal h63_out, h127_out, h191_out, h255_out    : std_logic_vector(Wh-1 downto 0);
signal h64_out, h128_out, h192_out, h256_out    : std_logic_vector(Wh-1 downto 0);

signal h01_en, h65_en , h129_en, h193_en    : std_logic;
signal h02_en, h66_en , h130_en, h194_en    : std_logic;
signal h03_en, h67_en , h131_en, h195_en    : std_logic;
signal h04_en, h68_en , h132_en, h196_en    : std_logic;
signal h05_en, h69_en , h133_en, h197_en    : std_logic;
signal h06_en, h70_en , h134_en, h198_en    : std_logic;
signal h07_en, h71_en , h135_en, h199_en    : std_logic;
signal h08_en, h72_en , h136_en, h200_en    : std_logic;
signal h09_en, h73_en , h137_en, h201_en    : std_logic;
signal h10_en, h74_en , h138_en, h202_en    : std_logic;
signal h11_en, h75_en , h139_en, h203_en    : std_logic;
signal h12_en, h76_en , h140_en, h204_en    : std_logic;
signal h13_en, h77_en , h141_en, h205_en    : std_logic;
signal h14_en, h78_en , h142_en, h206_en    : std_logic;
signal h15_en, h79_en , h143_en, h207_en    : std_logic;
signal h16_en, h80_en , h144_en, h208_en    : std_logic;
signal h17_en, h81_en , h145_en, h209_en    : std_logic;
signal h18_en, h82_en , h146_en, h210_en    : std_logic;
signal h19_en, h83_en , h147_en, h211_en    : std_logic;
signal h20_en, h84_en , h148_en, h212_en    : std_logic;
signal h21_en, h85_en , h149_en, h213_en    : std_logic;
signal h22_en, h86_en , h150_en, h214_en    : std_logic;
signal h23_en, h87_en , h151_en, h215_en    : std_logic;
signal h24_en, h88_en , h152_en, h216_en    : std_logic;
signal h25_en, h89_en , h153_en, h217_en    : std_logic;
signal h26_en, h90_en , h154_en, h218_en    : std_logic;
signal h27_en, h91_en , h155_en, h219_en    : std_logic;
signal h28_en, h92_en , h156_en, h220_en    : std_logic;
signal h29_en, h93_en , h157_en, h221_en    : std_logic;
signal h30_en, h94_en , h158_en, h222_en    : std_logic;
signal h31_en, h95_en , h159_en, h223_en    : std_logic;
signal h32_en, h96_en , h160_en, h224_en    : std_logic;
signal h33_en, h97_en , h161_en, h225_en    : std_logic;
signal h34_en, h98_en , h162_en, h226_en    : std_logic;
signal h35_en, h99_en , h163_en, h227_en    : std_logic;
signal h36_en, h100_en, h164_en, h228_en    : std_logic;
signal h37_en, h101_en, h165_en, h229_en    : std_logic;
signal h38_en, h102_en, h166_en, h230_en    : std_logic;
signal h39_en, h103_en, h167_en, h231_en    : std_logic;
signal h40_en, h104_en, h168_en, h232_en    : std_logic;
signal h41_en, h105_en, h169_en, h233_en    : std_logic;
signal h42_en, h106_en, h170_en, h234_en    : std_logic;
signal h43_en, h107_en, h171_en, h235_en    : std_logic;
signal h44_en, h108_en, h172_en, h236_en    : std_logic;
signal h45_en, h109_en, h173_en, h237_en    : std_logic;
signal h46_en, h110_en, h174_en, h238_en    : std_logic;
signal h47_en, h111_en, h175_en, h239_en    : std_logic;
signal h48_en, h112_en, h176_en, h240_en    : std_logic;
signal h49_en, h113_en, h177_en, h241_en    : std_logic;
signal h50_en, h114_en, h178_en, h242_en    : std_logic;
signal h51_en, h115_en, h179_en, h243_en    : std_logic;
signal h52_en, h116_en, h180_en, h244_en    : std_logic;
signal h53_en, h117_en, h181_en, h245_en    : std_logic;
signal h54_en, h118_en, h182_en, h246_en    : std_logic;
signal h55_en, h119_en, h183_en, h247_en    : std_logic;
signal h56_en, h120_en, h184_en, h248_en    : std_logic;
signal h57_en, h121_en, h185_en, h249_en    : std_logic;
signal h58_en, h122_en, h186_en, h250_en    : std_logic;
signal h59_en, h123_en, h187_en, h251_en    : std_logic;
signal h60_en, h124_en, h188_en, h252_en    : std_logic;
signal h61_en, h125_en, h189_en, h253_en    : std_logic;
signal h62_en, h126_en, h190_en, h254_en    : std_logic;
signal h63_en, h127_en, h191_en, h255_en    : std_logic;
signal h64_en, h128_en, h192_en, h256_en    : std_logic;

signal buff01_out, buff02_out, buff03_out, buff04_out, buff05_out, buff06_out, buff07_out, buff08_out, buff09_out, buff10_out, buff11_out, buff12_out, buff13_out, buff14_out, buff15_out, buff16_out, buff17_out, buff18_out, buff19_out, buff20_out, buff21_out, buff22_out, buff23_out, buff24_out, buff25_out, buff26_out, buff27_out, buff28_out, buff29_out, buff30_out, buff31_out, buff32_out : std_logic_vector(Wb-1 downto 0);
signal buff33_out, buff34_out, buff35_out, buff36_out, buff37_out, buff38_out, buff39_out, buff40_out, buff41_out, buff42_out, buff43_out, buff44_out, buff45_out, buff46_out, buff47_out, buff48_out, buff49_out, buff50_out, buff51_out, buff52_out, buff53_out, buff54_out, buff55_out, buff56_out, buff57_out, buff58_out, buff59_out, buff60_out, buff61_out, buff62_out, buff63_out, buff64_out : std_logic_vector(Wb-1 downto 0);
signal buff65_out, buff66_out, buff67_out, buff68_out, buff69_out, buff70_out, buff71_out, buff72_out, buff73_out, buff74_out, buff75_out, buff76_out, buff77_out, buff78_out, buff79_out, buff80_out, buff81_out, buff82_out, buff83_out, buff84_out, buff85_out, buff86_out, buff87_out, buff88_out, buff89_out, buff90_out, buff91_out, buff92_out, buff93_out, buff94_out, buff95_out, buff96_out : std_logic_vector(Wb-1 downto 0);
signal buff97_out, buff98_out, buff99_out, buff100_out, buff101_out, buff102_out, buff103_out, buff104_out, buff105_out, buff106_out, buff107_out, buff108_out, buff109_out, buff110_out, buff111_out, buff112_out, buff113_out, buff114_out, buff115_out, buff116_out, buff117_out, buff118_out, buff119_out, buff120_out, buff121_out, buff122_out, buff123_out, buff124_out, buff125_out, buff126_out, buff127_out, buff128_out : std_logic_vector(Wb-1 downto 0);
signal buff129_out,buff130_out,buff131_out,buff132_out,buff133_out,buff134_out,buff135_out,buff136_out,buff137_out,buff138_out,buff139_out,buff140_out,buff141_out,buff142_out,buff143_out,buff144_out,buff145_out,buff146_out,buff147_out,buff148_out,buff149_out,buff150_out,buff151_out,buff152_out,buff153_out,buff154_out,buff155_out,buff156_out,buff157_out,buff158_out,buff159_out,buff160_out: std_logic_vector(Wb-1 downto 0);
signal buff161_out,buff162_out,buff163_out,buff164_out,buff165_out,buff166_out,buff167_out,buff168_out,buff169_out,buff170_out,buff171_out,buff172_out,buff173_out,buff174_out,buff175_out,buff176_out,buff177_out,buff178_out,buff179_out,buff180_out,buff181_out,buff182_out,buff183_out,buff184_out,buff185_out,buff186_out,buff187_out,buff188_out,buff189_out,buff190_out,buff191_out,buff192_out: std_logic_vector(Wb-1 downto 0);
signal buff193_out,buff194_out,buff195_out,buff196_out,buff197_out,buff198_out,buff199_out,buff200_out,buff201_out,buff202_out,buff203_out,buff204_out,buff205_out,buff206_out,buff207_out,buff208_out,buff209_out,buff210_out,buff211_out,buff212_out,buff213_out,buff214_out,buff215_out,buff216_out,buff217_out,buff218_out,buff219_out,buff220_out,buff221_out,buff222_out,buff223_out,buff224_out: std_logic_vector(Wb-1 downto 0);
signal buff225_out,buff226_out,buff227_out,buff228_out,buff229_out,buff230_out,buff231_out,buff232_out,buff233_out,buff234_out,buff235_out,buff236_out,buff237_out,buff238_out,buff239_out,buff240_out,buff241_out,buff242_out,buff243_out,buff244_out,buff245_out,buff246_out,buff247_out,buff248_out,buff249_out,buff250_out,buff251_out,buff252_out,buff253_out,buff254_out,buff255_out,buff256_out: std_logic_vector(Wb-1 downto 0);


signal b_rd : std_logic_vector (256-1 downto 0);

begin

g_Huff_enc_en: if Huff_enc_en = TRUE generate
   Huf01 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d01_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h01_out, en_out => h01_en, eof_out => eof_out);
   Huf02 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d02_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h02_out, en_out => h02_en, eof_out => open);
   Huf03 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d03_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h03_out, en_out => h03_en, eof_out => open);
   Huf04 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d04_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h04_out, en_out => h04_en, eof_out => open);
   Huf05 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d05_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h05_out, en_out => h05_en, eof_out => open);
   Huf06 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d06_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h06_out, en_out => h06_en, eof_out => open);
   Huf07 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d07_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h07_out, en_out => h07_en, eof_out => open);
   Huf08 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d08_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h08_out, en_out => h08_en, eof_out => open);
   Huf09 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d09_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h09_out, en_out => h09_en, eof_out => open);
   Huf10 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d10_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h10_out, en_out => h10_en, eof_out => open);
   Huf11 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d11_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h11_out, en_out => h11_en, eof_out => open);
   Huf12 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d12_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h12_out, en_out => h12_en, eof_out => open);
   Huf13 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d13_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h13_out, en_out => h13_en, eof_out => open);
   Huf14 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d14_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h14_out, en_out => h14_en, eof_out => open);
   Huf15 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d15_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h15_out, en_out => h15_en, eof_out => open);
   Huf16 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d16_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h16_out, en_out => h16_en, eof_out => open);
   Huf17 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d17_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h17_out, en_out => h17_en, eof_out => open);
   Huf18 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d18_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h18_out, en_out => h18_en, eof_out => open);
   Huf19 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d19_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h19_out, en_out => h19_en, eof_out => open);
   Huf20 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d20_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h20_out, en_out => h20_en, eof_out => open);
   Huf21 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d21_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h21_out, en_out => h21_en, eof_out => open);
   Huf22 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d22_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h22_out, en_out => h22_en, eof_out => open);
   Huf23 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d23_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h23_out, en_out => h23_en, eof_out => open);
   Huf24 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d24_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h24_out, en_out => h24_en, eof_out => open);
   Huf25 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d25_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h25_out, en_out => h25_en, eof_out => open);
   Huf26 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d26_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h26_out, en_out => h26_en, eof_out => open);
   Huf27 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d27_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h27_out, en_out => h27_en, eof_out => open);
   Huf28 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d28_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h28_out, en_out => h28_en, eof_out => open);
   Huf29 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d29_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h29_out, en_out => h29_en, eof_out => open);
   Huf30 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d30_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h30_out, en_out => h30_en, eof_out => open);
   Huf31 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d31_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h31_out, en_out => h31_en, eof_out => open);
   Huf32 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d32_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h32_out, en_out => h32_en, eof_out => open);
   Huf33 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d33_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h33_out, en_out => h33_en, eof_out => open);
   Huf34 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d34_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h34_out, en_out => h34_en, eof_out => open);
   Huf35 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d35_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h35_out, en_out => h35_en, eof_out => open);
   Huf36 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d36_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h36_out, en_out => h36_en, eof_out => open);
   Huf37 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d37_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h37_out, en_out => h37_en, eof_out => open);
   Huf38 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d38_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h38_out, en_out => h38_en, eof_out => open);
   Huf39 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d39_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h39_out, en_out => h39_en, eof_out => open);
   Huf40 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d40_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h40_out, en_out => h40_en, eof_out => open);
   Huf41 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d41_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h41_out, en_out => h41_en, eof_out => open);
   Huf42 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d42_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h42_out, en_out => h42_en, eof_out => open);
   Huf43 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d43_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h43_out, en_out => h43_en, eof_out => open);
   Huf44 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d44_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h44_out, en_out => h44_en, eof_out => open);
   Huf45 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d45_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h45_out, en_out => h45_en, eof_out => open);
   Huf46 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d46_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h46_out, en_out => h46_en, eof_out => open);
   Huf47 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d47_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h47_out, en_out => h47_en, eof_out => open);
   Huf48 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d48_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h48_out, en_out => h48_en, eof_out => open);
   Huf49 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d49_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h49_out, en_out => h49_en, eof_out => open);
   Huf50 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d50_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h50_out, en_out => h50_en, eof_out => open);
   Huf51 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d51_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h51_out, en_out => h51_en, eof_out => open);
   Huf52 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d52_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h52_out, en_out => h52_en, eof_out => open);
   Huf53 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d53_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h53_out, en_out => h53_en, eof_out => open);
   Huf54 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d54_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h54_out, en_out => h54_en, eof_out => open);
   Huf55 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d55_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h55_out, en_out => h55_en, eof_out => open);
   Huf56 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d56_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h56_out, en_out => h56_en, eof_out => open);
   Huf57 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d57_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h57_out, en_out => h57_en, eof_out => open);
   Huf58 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d58_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h58_out, en_out => h58_en, eof_out => open);
   Huf59 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d59_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h59_out, en_out => h59_en, eof_out => open);
   Huf60 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d60_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h60_out, en_out => h60_en, eof_out => open);
   Huf61 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d61_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h61_out, en_out => h61_en, eof_out => open);
   Huf62 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d62_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h62_out, en_out => h62_en, eof_out => open);
   Huf63 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d63_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h63_out, en_out => h63_en, eof_out => open);
   Huf64 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d64_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h64_out, en_out => h64_en, eof_out => open);

   Huf65 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d65_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h65_out , en_out => h65_en , eof_out => open);
   Huf66 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d66_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h66_out , en_out => h66_en , eof_out => open);
   Huf67 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d67_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h67_out , en_out => h67_en , eof_out => open);
   Huf68 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d68_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h68_out , en_out => h68_en , eof_out => open);
   Huf69 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d69_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h69_out , en_out => h69_en , eof_out => open);
   Huf70 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d70_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h70_out , en_out => h70_en , eof_out => open);
   Huf71 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d71_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h71_out , en_out => h71_en , eof_out => open);
   Huf72 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d72_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h72_out , en_out => h72_en , eof_out => open);
   Huf73 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d73_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h73_out , en_out => h73_en , eof_out => open);
   Huf74 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d74_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h74_out , en_out => h74_en , eof_out => open);
   Huf75 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d75_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h75_out , en_out => h75_en , eof_out => open);
   Huf76 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d76_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h76_out , en_out => h76_en , eof_out => open);
   Huf77 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d77_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h77_out , en_out => h77_en , eof_out => open);
   Huf78 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d78_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h78_out , en_out => h78_en , eof_out => open);
   Huf79 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d79_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h79_out , en_out => h79_en , eof_out => open);
   Huf80 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d80_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h80_out , en_out => h80_en , eof_out => open);
   Huf81 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d81_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h81_out , en_out => h81_en , eof_out => open);
   Huf82 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d82_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h82_out , en_out => h82_en , eof_out => open);
   Huf83 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d83_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h83_out , en_out => h83_en , eof_out => open);
   Huf84 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d84_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h84_out , en_out => h84_en , eof_out => open);
   Huf85 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d85_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h85_out , en_out => h85_en , eof_out => open);
   Huf86 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d86_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h86_out , en_out => h86_en , eof_out => open);
   Huf87 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d87_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h87_out , en_out => h87_en , eof_out => open);
   Huf88 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d88_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h88_out , en_out => h88_en , eof_out => open);
   Huf89 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d89_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h89_out , en_out => h89_en , eof_out => open);
   Huf90 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d90_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h90_out , en_out => h90_en , eof_out => open);
   Huf91 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d91_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h91_out , en_out => h91_en , eof_out => open);
   Huf92 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d92_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h92_out , en_out => h92_en , eof_out => open);
   Huf93 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d93_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h93_out , en_out => h93_en , eof_out => open);
   Huf94 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d94_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h94_out , en_out => h94_en , eof_out => open);
   Huf95 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d95_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h95_out , en_out => h95_en , eof_out => open);
   Huf96 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d96_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h96_out , en_out => h96_en , eof_out => open);
   Huf97 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d97_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h97_out , en_out => h97_en , eof_out => open);
   Huf98 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d98_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h98_out , en_out => h98_en , eof_out => open);
   Huf99 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d99_in , en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h99_out , en_out => h99_en , eof_out => open);
   Huf100: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d100_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h100_out, en_out => h100_en, eof_out => open);
   Huf101: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d101_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h101_out, en_out => h101_en, eof_out => open);
   Huf102: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d102_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h102_out, en_out => h102_en, eof_out => open);
   Huf103: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d103_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h103_out, en_out => h103_en, eof_out => open);
   Huf104: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d104_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h104_out, en_out => h104_en, eof_out => open);
   Huf105: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d105_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h105_out, en_out => h105_en, eof_out => open);
   Huf106: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d106_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h106_out, en_out => h106_en, eof_out => open);
   Huf107: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d107_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h107_out, en_out => h107_en, eof_out => open);
   Huf108: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d108_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h108_out, en_out => h108_en, eof_out => open);
   Huf109: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d109_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h109_out, en_out => h109_en, eof_out => open);
   Huf110: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d110_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h110_out, en_out => h110_en, eof_out => open);
   Huf111: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d111_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h111_out, en_out => h111_en, eof_out => open);
   Huf112: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d112_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h112_out, en_out => h112_en, eof_out => open);
   Huf113: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d113_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h113_out, en_out => h113_en, eof_out => open);
   Huf114: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d114_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h114_out, en_out => h114_en, eof_out => open);
   Huf115: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d115_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h115_out, en_out => h115_en, eof_out => open);
   Huf116: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d116_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h116_out, en_out => h116_en, eof_out => open);
   Huf117: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d117_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h117_out, en_out => h117_en, eof_out => open);
   Huf118: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d118_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h118_out, en_out => h118_en, eof_out => open);
   Huf119: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d119_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h119_out, en_out => h119_en, eof_out => open);
   Huf120: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d120_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h120_out, en_out => h120_en, eof_out => open);
   Huf121: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d121_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h121_out, en_out => h121_en, eof_out => open);
   Huf122: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d122_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h122_out, en_out => h122_en, eof_out => open);
   Huf123: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d123_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h123_out, en_out => h123_en, eof_out => open);
   Huf124: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d124_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h124_out, en_out => h124_en, eof_out => open);
   Huf125: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d125_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h125_out, en_out => h125_en, eof_out => open);
   Huf126: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d126_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h126_out, en_out => h126_en, eof_out => open);
   Huf127: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d127_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h127_out, en_out => h127_en, eof_out => open);
   Huf128: Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d128_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h128_out, en_out => h128_en, eof_out => open);

   Huf129 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d129_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h129_out, en_out => h129_en, eof_out => open);
   Huf130 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d130_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h130_out, en_out => h130_en, eof_out => open);
   Huf131 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d131_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h131_out, en_out => h131_en, eof_out => open);
   Huf132 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d132_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h132_out, en_out => h132_en, eof_out => open);
   Huf133 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d133_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h133_out, en_out => h133_en, eof_out => open);
   Huf134 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d134_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h134_out, en_out => h134_en, eof_out => open);
   Huf135 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d135_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h135_out, en_out => h135_en, eof_out => open);
   Huf136 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d136_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h136_out, en_out => h136_en, eof_out => open);
   Huf137 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d137_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h137_out, en_out => h137_en, eof_out => open);
   Huf138 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d138_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h138_out, en_out => h138_en, eof_out => open);
   Huf139 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d139_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h139_out, en_out => h139_en, eof_out => open);
   Huf140 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d140_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h140_out, en_out => h140_en, eof_out => open);
   Huf141 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d141_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h141_out, en_out => h141_en, eof_out => open);
   Huf142 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d142_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h142_out, en_out => h142_en, eof_out => open);
   Huf143 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d143_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h143_out, en_out => h143_en, eof_out => open);
   Huf144 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d144_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h144_out, en_out => h144_en, eof_out => open);
   Huf145 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d145_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h145_out, en_out => h145_en, eof_out => open);
   Huf146 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d146_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h146_out, en_out => h146_en, eof_out => open);
   Huf147 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d147_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h147_out, en_out => h147_en, eof_out => open);
   Huf148 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d148_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h148_out, en_out => h148_en, eof_out => open);
   Huf149 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d149_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h149_out, en_out => h149_en, eof_out => open);
   Huf150 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d150_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h150_out, en_out => h150_en, eof_out => open);
   Huf151 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d151_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h151_out, en_out => h151_en, eof_out => open);
   Huf152 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d152_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h152_out, en_out => h152_en, eof_out => open);
   Huf153 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d153_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h153_out, en_out => h153_en, eof_out => open);
   Huf154 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d154_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h154_out, en_out => h154_en, eof_out => open);
   Huf155 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d155_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h155_out, en_out => h155_en, eof_out => open);
   Huf156 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d156_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h156_out, en_out => h156_en, eof_out => open);
   Huf157 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d157_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h157_out, en_out => h157_en, eof_out => open);
   Huf158 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d158_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h158_out, en_out => h158_en, eof_out => open);
   Huf159 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d159_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h159_out, en_out => h159_en, eof_out => open);
   Huf160 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d160_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h160_out, en_out => h160_en, eof_out => open);
   Huf161 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d161_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h161_out, en_out => h161_en, eof_out => open);
   Huf162 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d162_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h162_out, en_out => h162_en, eof_out => open);
   Huf163 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d163_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h163_out, en_out => h163_en, eof_out => open);
   Huf164 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d164_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h164_out, en_out => h164_en, eof_out => open);
   Huf165 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d165_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h165_out, en_out => h165_en, eof_out => open);
   Huf166 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d166_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h166_out, en_out => h166_en, eof_out => open);
   Huf167 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d167_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h167_out, en_out => h167_en, eof_out => open);
   Huf168 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d168_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h168_out, en_out => h168_en, eof_out => open);
   Huf169 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d169_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h169_out, en_out => h169_en, eof_out => open);
   Huf170 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d170_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h170_out, en_out => h170_en, eof_out => open);
   Huf171 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d171_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h171_out, en_out => h171_en, eof_out => open);
   Huf172 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d172_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h172_out, en_out => h172_en, eof_out => open);
   Huf173 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d173_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h173_out, en_out => h173_en, eof_out => open);
   Huf174 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d174_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h174_out, en_out => h174_en, eof_out => open);
   Huf175 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d175_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h175_out, en_out => h175_en, eof_out => open);
   Huf176 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d176_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h176_out, en_out => h176_en, eof_out => open);
   Huf177 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d177_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h177_out, en_out => h177_en, eof_out => open);
   Huf178 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d178_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h178_out, en_out => h178_en, eof_out => open);
   Huf179 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d179_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h179_out, en_out => h179_en, eof_out => open);
   Huf180 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d180_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h180_out, en_out => h180_en, eof_out => open);
   Huf181 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d181_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h181_out, en_out => h181_en, eof_out => open);
   Huf182 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d182_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h182_out, en_out => h182_en, eof_out => open);
   Huf183 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d183_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h183_out, en_out => h183_en, eof_out => open);
   Huf184 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d184_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h184_out, en_out => h184_en, eof_out => open);
   Huf185 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d185_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h185_out, en_out => h185_en, eof_out => open);
   Huf186 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d186_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h186_out, en_out => h186_en, eof_out => open);
   Huf187 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d187_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h187_out, en_out => h187_en, eof_out => open);
   Huf188 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d188_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h188_out, en_out => h188_en, eof_out => open);
   Huf189 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d189_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h189_out, en_out => h189_en, eof_out => open);
   Huf190 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d190_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h190_out, en_out => h190_en, eof_out => open);
   Huf191 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d191_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h191_out, en_out => h191_en, eof_out => open);
   Huf192 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d192_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h192_out, en_out => h192_en, eof_out => open);

   Huf193 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d193_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h193_out, en_out => h193_en, eof_out => open);
   Huf194 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d194_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h194_out, en_out => h194_en, eof_out => open);
   Huf195 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d195_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h195_out, en_out => h195_en, eof_out => open);
   Huf196 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d196_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h196_out, en_out => h196_en, eof_out => open);
   Huf197 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d197_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h197_out, en_out => h197_en, eof_out => open);
   Huf198 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d198_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h198_out, en_out => h198_en, eof_out => open);
   Huf199 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d199_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h199_out, en_out => h199_en, eof_out => open);
   Huf200 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d200_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h200_out, en_out => h200_en, eof_out => open);
   Huf201 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d201_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h201_out, en_out => h201_en, eof_out => open);
   Huf202 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d202_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h202_out, en_out => h202_en, eof_out => open);
   Huf203 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d203_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h203_out, en_out => h203_en, eof_out => open);
   Huf204 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d204_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h204_out, en_out => h204_en, eof_out => open);
   Huf205 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d205_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h205_out, en_out => h205_en, eof_out => open);
   Huf206 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d206_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h206_out, en_out => h206_en, eof_out => open);
   Huf207 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d207_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h207_out, en_out => h207_en, eof_out => open);
   Huf208 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d208_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h208_out, en_out => h208_en, eof_out => open);
   Huf209 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d209_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h209_out, en_out => h209_en, eof_out => open);
   Huf210 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d210_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h210_out, en_out => h210_en, eof_out => open);
   Huf211 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d211_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h211_out, en_out => h211_en, eof_out => open);
   Huf212 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d212_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h212_out, en_out => h212_en, eof_out => open);
   Huf213 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d213_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h213_out, en_out => h213_en, eof_out => open);
   Huf214 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d214_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h214_out, en_out => h214_en, eof_out => open);
   Huf215 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d215_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h215_out, en_out => h215_en, eof_out => open);
   Huf216 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d216_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h216_out, en_out => h216_en, eof_out => open);
   Huf217 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d217_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h217_out, en_out => h217_en, eof_out => open);
   Huf218 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d218_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h218_out, en_out => h218_en, eof_out => open);
   Huf219 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d219_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h219_out, en_out => h219_en, eof_out => open);
   Huf220 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d220_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h220_out, en_out => h220_en, eof_out => open);
   Huf221 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d221_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h221_out, en_out => h221_en, eof_out => open);
   Huf222 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d222_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h222_out, en_out => h222_en, eof_out => open);
   Huf223 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d223_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h223_out, en_out => h223_en, eof_out => open);
   Huf224 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d224_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h224_out, en_out => h224_en, eof_out => open);
   Huf225 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d225_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h225_out, en_out => h225_en, eof_out => open);
   Huf226 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d226_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h226_out, en_out => h226_en, eof_out => open);
   Huf227 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d227_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h227_out, en_out => h227_en, eof_out => open);
   Huf228 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d228_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h228_out, en_out => h228_en, eof_out => open);
   Huf229 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d229_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h229_out, en_out => h229_en, eof_out => open);
   Huf230 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d230_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h230_out, en_out => h230_en, eof_out => open);
   Huf231 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d231_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h231_out, en_out => h231_en, eof_out => open);
   Huf232 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d232_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h232_out, en_out => h232_en, eof_out => open);
   Huf233 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d233_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h233_out, en_out => h233_en, eof_out => open);
   Huf234 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d234_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h234_out, en_out => h234_en, eof_out => open);
   Huf235 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d235_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h235_out, en_out => h235_en, eof_out => open);
   Huf236 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d236_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h236_out, en_out => h236_en, eof_out => open);
   Huf237 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d237_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h237_out, en_out => h237_en, eof_out => open);
   Huf238 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d238_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h238_out, en_out => h238_en, eof_out => open);
   Huf239 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d239_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h239_out, en_out => h239_en, eof_out => open);
   Huf240 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d240_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h240_out, en_out => h240_en, eof_out => open);
   Huf241 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d241_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h241_out, en_out => h241_en, eof_out => open);
   Huf242 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d242_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h242_out, en_out => h242_en, eof_out => open);
   Huf243 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d243_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h243_out, en_out => h243_en, eof_out => open);
   Huf244 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d244_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h244_out, en_out => h244_en, eof_out => open);
   Huf245 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d245_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h245_out, en_out => h245_en, eof_out => open);
   Huf246 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d246_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h246_out, en_out => h246_en, eof_out => open);
   Huf247 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d247_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h247_out, en_out => h247_en, eof_out => open);
   Huf248 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d248_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h248_out, en_out => h248_en, eof_out => open);
   Huf249 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d249_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h249_out, en_out => h249_en, eof_out => open);
   Huf250 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d250_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h250_out, en_out => h250_en, eof_out => open);
   Huf251 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d251_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h251_out, en_out => h251_en, eof_out => open);
   Huf252 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d252_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h252_out, en_out => h252_en, eof_out => open);
   Huf253 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d253_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h253_out, en_out => h253_en, eof_out => open);
   Huf254 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d254_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h254_out, en_out => h254_en, eof_out => open);
   Huf255 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d255_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h255_out, en_out => h255_en, eof_out => open);
   Huf256 : Huffman generic map(N => N, M => M, W => Wh) port map( clk =>clk, rst =>rst , init_en => init_en, alpha_data => alpha_data, alpha_code => alpha_code, alpha_width => alpha_width, d_in  => d256_in, en_in => en_in, sof_in=> sof_in, eof_in=> eof_in, d_out => h256_out, en_out => h256_en, eof_out => open);


end generate g_Huff_enc_en;

g_Huff_enc_dis: if Huff_enc_en = FALSE generate
   h01_out(h01_out'left downto d01_in'left + 1) <= (others => '0');   h01_out(d01_in'left downto 0) <= d01_in;   h01_en <= en_in;
   h02_out(h02_out'left downto d02_in'left + 1) <= (others => '0');   h02_out(d02_in'left downto 0) <= d02_in;   h02_en <= en_in;
   h03_out(h03_out'left downto d03_in'left + 1) <= (others => '0');   h03_out(d03_in'left downto 0) <= d03_in;   h03_en <= en_in;
   h04_out(h04_out'left downto d04_in'left + 1) <= (others => '0');   h04_out(d04_in'left downto 0) <= d04_in;   h04_en <= en_in;
   h05_out(h05_out'left downto d05_in'left + 1) <= (others => '0');   h05_out(d05_in'left downto 0) <= d05_in;   h05_en <= en_in;
   h06_out(h06_out'left downto d06_in'left + 1) <= (others => '0');   h06_out(d06_in'left downto 0) <= d06_in;   h06_en <= en_in;
   h07_out(h07_out'left downto d07_in'left + 1) <= (others => '0');   h07_out(d07_in'left downto 0) <= d07_in;   h07_en <= en_in;
   h08_out(h08_out'left downto d08_in'left + 1) <= (others => '0');   h08_out(d08_in'left downto 0) <= d08_in;   h08_en <= en_in;
   h09_out(h09_out'left downto d09_in'left + 1) <= (others => '0');   h09_out(d09_in'left downto 0) <= d09_in;   h09_en <= en_in;
   h10_out(h10_out'left downto d10_in'left + 1) <= (others => '0');   h10_out(d10_in'left downto 0) <= d10_in;   h10_en <= en_in;
   h11_out(h11_out'left downto d11_in'left + 1) <= (others => '0');   h11_out(d11_in'left downto 0) <= d11_in;   h11_en <= en_in;
   h12_out(h12_out'left downto d12_in'left + 1) <= (others => '0');   h12_out(d12_in'left downto 0) <= d12_in;   h12_en <= en_in;
   h13_out(h13_out'left downto d13_in'left + 1) <= (others => '0');   h13_out(d13_in'left downto 0) <= d13_in;   h13_en <= en_in;
   h14_out(h14_out'left downto d14_in'left + 1) <= (others => '0');   h14_out(d14_in'left downto 0) <= d14_in;   h14_en <= en_in;
   h15_out(h15_out'left downto d15_in'left + 1) <= (others => '0');   h15_out(d15_in'left downto 0) <= d15_in;   h15_en <= en_in;
   h16_out(h16_out'left downto d16_in'left + 1) <= (others => '0');   h16_out(d16_in'left downto 0) <= d16_in;   h16_en <= en_in;
   h17_out(h17_out'left downto d17_in'left + 1) <= (others => '0');   h17_out(d17_in'left downto 0) <= d17_in;   h17_en <= en_in;
   h18_out(h18_out'left downto d18_in'left + 1) <= (others => '0');   h18_out(d18_in'left downto 0) <= d18_in;   h18_en <= en_in;
   h19_out(h19_out'left downto d19_in'left + 1) <= (others => '0');   h19_out(d19_in'left downto 0) <= d19_in;   h19_en <= en_in;
   h20_out(h20_out'left downto d20_in'left + 1) <= (others => '0');   h20_out(d20_in'left downto 0) <= d20_in;   h20_en <= en_in;
   h21_out(h21_out'left downto d21_in'left + 1) <= (others => '0');   h21_out(d21_in'left downto 0) <= d21_in;   h21_en <= en_in;
   h22_out(h22_out'left downto d22_in'left + 1) <= (others => '0');   h22_out(d22_in'left downto 0) <= d22_in;   h22_en <= en_in;
   h23_out(h23_out'left downto d23_in'left + 1) <= (others => '0');   h23_out(d23_in'left downto 0) <= d23_in;   h23_en <= en_in;
   h24_out(h24_out'left downto d24_in'left + 1) <= (others => '0');   h24_out(d24_in'left downto 0) <= d24_in;   h24_en <= en_in;
   h25_out(h25_out'left downto d25_in'left + 1) <= (others => '0');   h25_out(d25_in'left downto 0) <= d25_in;   h25_en <= en_in;
   h26_out(h26_out'left downto d26_in'left + 1) <= (others => '0');   h26_out(d26_in'left downto 0) <= d26_in;   h26_en <= en_in;
   h27_out(h27_out'left downto d27_in'left + 1) <= (others => '0');   h27_out(d27_in'left downto 0) <= d27_in;   h27_en <= en_in;
   h28_out(h28_out'left downto d28_in'left + 1) <= (others => '0');   h28_out(d28_in'left downto 0) <= d28_in;   h28_en <= en_in;
   h29_out(h29_out'left downto d29_in'left + 1) <= (others => '0');   h29_out(d29_in'left downto 0) <= d29_in;   h29_en <= en_in;
   h30_out(h30_out'left downto d30_in'left + 1) <= (others => '0');   h30_out(d30_in'left downto 0) <= d30_in;   h30_en <= en_in;
   h31_out(h31_out'left downto d31_in'left + 1) <= (others => '0');   h31_out(d31_in'left downto 0) <= d31_in;   h31_en <= en_in;
   h32_out(h32_out'left downto d32_in'left + 1) <= (others => '0');   h32_out(d32_in'left downto 0) <= d32_in;   h32_en <= en_in;
   h33_out(h33_out'left downto d33_in'left + 1) <= (others => '0');   h33_out(d33_in'left downto 0) <= d33_in;   h33_en <= en_in;
   h34_out(h34_out'left downto d34_in'left + 1) <= (others => '0');   h34_out(d34_in'left downto 0) <= d34_in;   h34_en <= en_in;
   h35_out(h35_out'left downto d35_in'left + 1) <= (others => '0');   h35_out(d35_in'left downto 0) <= d35_in;   h35_en <= en_in;
   h36_out(h36_out'left downto d36_in'left + 1) <= (others => '0');   h36_out(d36_in'left downto 0) <= d36_in;   h36_en <= en_in;
   h37_out(h37_out'left downto d37_in'left + 1) <= (others => '0');   h37_out(d37_in'left downto 0) <= d37_in;   h37_en <= en_in;
   h38_out(h38_out'left downto d38_in'left + 1) <= (others => '0');   h38_out(d38_in'left downto 0) <= d38_in;   h38_en <= en_in;
   h39_out(h39_out'left downto d39_in'left + 1) <= (others => '0');   h39_out(d39_in'left downto 0) <= d39_in;   h39_en <= en_in;
   h40_out(h40_out'left downto d40_in'left + 1) <= (others => '0');   h40_out(d40_in'left downto 0) <= d40_in;   h40_en <= en_in;
   h41_out(h41_out'left downto d41_in'left + 1) <= (others => '0');   h41_out(d41_in'left downto 0) <= d41_in;   h41_en <= en_in;
   h42_out(h42_out'left downto d42_in'left + 1) <= (others => '0');   h42_out(d42_in'left downto 0) <= d42_in;   h42_en <= en_in;
   h43_out(h43_out'left downto d43_in'left + 1) <= (others => '0');   h43_out(d43_in'left downto 0) <= d43_in;   h43_en <= en_in;
   h44_out(h44_out'left downto d44_in'left + 1) <= (others => '0');   h44_out(d44_in'left downto 0) <= d44_in;   h44_en <= en_in;
   h45_out(h45_out'left downto d45_in'left + 1) <= (others => '0');   h45_out(d45_in'left downto 0) <= d45_in;   h45_en <= en_in;
   h46_out(h46_out'left downto d46_in'left + 1) <= (others => '0');   h46_out(d46_in'left downto 0) <= d46_in;   h46_en <= en_in;
   h47_out(h47_out'left downto d47_in'left + 1) <= (others => '0');   h47_out(d47_in'left downto 0) <= d47_in;   h47_en <= en_in;
   h48_out(h48_out'left downto d48_in'left + 1) <= (others => '0');   h48_out(d48_in'left downto 0) <= d48_in;   h48_en <= en_in;
   h49_out(h49_out'left downto d49_in'left + 1) <= (others => '0');   h49_out(d49_in'left downto 0) <= d49_in;   h49_en <= en_in;
   h50_out(h50_out'left downto d50_in'left + 1) <= (others => '0');   h50_out(d50_in'left downto 0) <= d50_in;   h50_en <= en_in;
   h51_out(h51_out'left downto d51_in'left + 1) <= (others => '0');   h51_out(d51_in'left downto 0) <= d51_in;   h51_en <= en_in;
   h52_out(h52_out'left downto d52_in'left + 1) <= (others => '0');   h52_out(d52_in'left downto 0) <= d52_in;   h52_en <= en_in;
   h53_out(h53_out'left downto d53_in'left + 1) <= (others => '0');   h53_out(d53_in'left downto 0) <= d53_in;   h53_en <= en_in;
   h54_out(h54_out'left downto d54_in'left + 1) <= (others => '0');   h54_out(d54_in'left downto 0) <= d54_in;   h54_en <= en_in;
   h55_out(h55_out'left downto d55_in'left + 1) <= (others => '0');   h55_out(d55_in'left downto 0) <= d55_in;   h55_en <= en_in;
   h56_out(h56_out'left downto d56_in'left + 1) <= (others => '0');   h56_out(d56_in'left downto 0) <= d56_in;   h56_en <= en_in;
   h57_out(h57_out'left downto d57_in'left + 1) <= (others => '0');   h57_out(d57_in'left downto 0) <= d57_in;   h57_en <= en_in;
   h58_out(h58_out'left downto d58_in'left + 1) <= (others => '0');   h58_out(d58_in'left downto 0) <= d58_in;   h58_en <= en_in;
   h59_out(h59_out'left downto d59_in'left + 1) <= (others => '0');   h59_out(d59_in'left downto 0) <= d59_in;   h59_en <= en_in;
   h60_out(h60_out'left downto d60_in'left + 1) <= (others => '0');   h60_out(d60_in'left downto 0) <= d60_in;   h60_en <= en_in;
   h61_out(h61_out'left downto d61_in'left + 1) <= (others => '0');   h61_out(d61_in'left downto 0) <= d61_in;   h61_en <= en_in;
   h62_out(h62_out'left downto d62_in'left + 1) <= (others => '0');   h62_out(d62_in'left downto 0) <= d62_in;   h62_en <= en_in;
   h63_out(h63_out'left downto d63_in'left + 1) <= (others => '0');   h63_out(d63_in'left downto 0) <= d63_in;   h63_en <= en_in;
   h64_out(h64_out'left downto d64_in'left + 1) <= (others => '0');   h64_out(d64_in'left downto 0) <= d64_in;   h64_en <= en_in;

   h65_out (h65_out 'left downto d65_in'left  + 1) <= (others => '0');   h65_out (d65_in 'left downto 0) <= d65_in;   h65_en  <= en_in;
   h66_out (h66_out 'left downto d66_in'left  + 1) <= (others => '0');   h66_out (d66_in 'left downto 0) <= d66_in;   h66_en  <= en_in;
   h67_out (h67_out 'left downto d67_in'left  + 1) <= (others => '0');   h67_out (d67_in 'left downto 0) <= d67_in;   h67_en  <= en_in;
   h68_out (h68_out 'left downto d68_in'left  + 1) <= (others => '0');   h68_out (d68_in 'left downto 0) <= d68_in;   h68_en  <= en_in;
   h69_out (h69_out 'left downto d69_in'left  + 1) <= (others => '0');   h69_out (d69_in 'left downto 0) <= d69_in;   h69_en  <= en_in;
   h70_out (h70_out 'left downto d70_in'left  + 1) <= (others => '0');   h70_out (d70_in 'left downto 0) <= d70_in;   h70_en  <= en_in;
   h71_out (h71_out 'left downto d71_in'left  + 1) <= (others => '0');   h71_out (d71_in 'left downto 0) <= d71_in;   h71_en  <= en_in;
   h72_out (h72_out 'left downto d72_in'left  + 1) <= (others => '0');   h72_out (d72_in 'left downto 0) <= d72_in;   h72_en  <= en_in;
   h73_out (h73_out 'left downto d73_in'left  + 1) <= (others => '0');   h73_out (d73_in 'left downto 0) <= d73_in;   h73_en  <= en_in;
   h74_out (h74_out 'left downto d74_in'left  + 1) <= (others => '0');   h74_out (d74_in 'left downto 0) <= d74_in;   h74_en  <= en_in;
   h75_out (h75_out 'left downto d75_in'left  + 1) <= (others => '0');   h75_out (d75_in 'left downto 0) <= d75_in;   h75_en  <= en_in;
   h76_out (h76_out 'left downto d76_in'left  + 1) <= (others => '0');   h76_out (d76_in 'left downto 0) <= d76_in;   h76_en  <= en_in;
   h77_out (h77_out 'left downto d77_in'left  + 1) <= (others => '0');   h77_out (d77_in 'left downto 0) <= d77_in;   h77_en  <= en_in;
   h78_out (h78_out 'left downto d78_in'left  + 1) <= (others => '0');   h78_out (d78_in 'left downto 0) <= d78_in;   h78_en  <= en_in;
   h79_out (h79_out 'left downto d79_in'left  + 1) <= (others => '0');   h79_out (d79_in 'left downto 0) <= d79_in;   h79_en  <= en_in;
   h80_out (h80_out 'left downto d80_in'left  + 1) <= (others => '0');   h80_out (d80_in 'left downto 0) <= d80_in;   h80_en  <= en_in;
   h81_out (h81_out 'left downto d81_in'left  + 1) <= (others => '0');   h81_out (d81_in 'left downto 0) <= d81_in;   h81_en  <= en_in;
   h82_out (h82_out 'left downto d82_in'left  + 1) <= (others => '0');   h82_out (d82_in 'left downto 0) <= d82_in;   h82_en  <= en_in;
   h83_out (h83_out 'left downto d83_in'left  + 1) <= (others => '0');   h83_out (d83_in 'left downto 0) <= d83_in;   h83_en  <= en_in;
   h84_out (h84_out 'left downto d84_in'left  + 1) <= (others => '0');   h84_out (d84_in 'left downto 0) <= d84_in;   h84_en  <= en_in;
   h85_out (h85_out 'left downto d85_in'left  + 1) <= (others => '0');   h85_out (d85_in 'left downto 0) <= d85_in;   h85_en  <= en_in;
   h86_out (h86_out 'left downto d86_in'left  + 1) <= (others => '0');   h86_out (d86_in 'left downto 0) <= d86_in;   h86_en  <= en_in;
   h87_out (h87_out 'left downto d87_in'left  + 1) <= (others => '0');   h87_out (d87_in 'left downto 0) <= d87_in;   h87_en  <= en_in;
   h88_out (h88_out 'left downto d88_in'left  + 1) <= (others => '0');   h88_out (d88_in 'left downto 0) <= d88_in;   h88_en  <= en_in;
   h89_out (h89_out 'left downto d89_in'left  + 1) <= (others => '0');   h89_out (d89_in 'left downto 0) <= d89_in;   h89_en  <= en_in;
   h90_out (h90_out 'left downto d90_in'left  + 1) <= (others => '0');   h90_out (d90_in 'left downto 0) <= d90_in;   h90_en  <= en_in;
   h91_out (h91_out 'left downto d91_in'left  + 1) <= (others => '0');   h91_out (d91_in 'left downto 0) <= d91_in;   h91_en  <= en_in;
   h92_out (h92_out 'left downto d92_in'left  + 1) <= (others => '0');   h92_out (d92_in 'left downto 0) <= d92_in;   h92_en  <= en_in;
   h93_out (h93_out 'left downto d93_in'left  + 1) <= (others => '0');   h93_out (d93_in 'left downto 0) <= d93_in;   h93_en  <= en_in;
   h94_out (h94_out 'left downto d94_in'left  + 1) <= (others => '0');   h94_out (d94_in 'left downto 0) <= d94_in;   h94_en  <= en_in;
   h95_out (h95_out 'left downto d95_in'left  + 1) <= (others => '0');   h95_out (d95_in 'left downto 0) <= d95_in;   h95_en  <= en_in;
   h96_out (h96_out 'left downto d96_in'left  + 1) <= (others => '0');   h96_out (d96_in 'left downto 0) <= d96_in;   h96_en  <= en_in;
   h97_out (h97_out 'left downto d97_in'left  + 1) <= (others => '0');   h97_out (d97_in 'left downto 0) <= d97_in;   h97_en  <= en_in;
   h98_out (h98_out 'left downto d98_in'left  + 1) <= (others => '0');   h98_out (d98_in 'left downto 0) <= d98_in;   h98_en  <= en_in;
   h99_out (h99_out 'left downto d99_in'left  + 1) <= (others => '0');   h99_out (d99_in 'left downto 0) <= d99_in;   h99_en  <= en_in;
   h100_out(h100_out'left downto d100_in'left + 1) <= (others => '0');   h100_out(d100_in'left downto 0) <= d100_in;  h100_en <= en_in;
   h101_out(h101_out'left downto d101_in'left + 1) <= (others => '0');   h101_out(d101_in'left downto 0) <= d101_in;  h101_en <= en_in;
   h102_out(h102_out'left downto d102_in'left + 1) <= (others => '0');   h102_out(d102_in'left downto 0) <= d102_in;  h102_en <= en_in;
   h103_out(h103_out'left downto d103_in'left + 1) <= (others => '0');   h103_out(d103_in'left downto 0) <= d103_in;  h103_en <= en_in;
   h104_out(h104_out'left downto d104_in'left + 1) <= (others => '0');   h104_out(d104_in'left downto 0) <= d104_in;  h104_en <= en_in;
   h105_out(h105_out'left downto d105_in'left + 1) <= (others => '0');   h105_out(d105_in'left downto 0) <= d105_in;  h105_en <= en_in;
   h106_out(h106_out'left downto d106_in'left + 1) <= (others => '0');   h106_out(d106_in'left downto 0) <= d106_in;  h106_en <= en_in;
   h107_out(h107_out'left downto d107_in'left + 1) <= (others => '0');   h107_out(d107_in'left downto 0) <= d107_in;  h107_en <= en_in;
   h108_out(h108_out'left downto d108_in'left + 1) <= (others => '0');   h108_out(d108_in'left downto 0) <= d108_in;  h108_en <= en_in;
   h109_out(h109_out'left downto d109_in'left + 1) <= (others => '0');   h109_out(d109_in'left downto 0) <= d109_in;  h109_en <= en_in;
   h110_out(h110_out'left downto d110_in'left + 1) <= (others => '0');   h110_out(d110_in'left downto 0) <= d110_in;  h110_en <= en_in;
   h111_out(h111_out'left downto d111_in'left + 1) <= (others => '0');   h111_out(d111_in'left downto 0) <= d111_in;  h111_en <= en_in;
   h112_out(h112_out'left downto d112_in'left + 1) <= (others => '0');   h112_out(d112_in'left downto 0) <= d112_in;  h112_en <= en_in;
   h113_out(h113_out'left downto d113_in'left + 1) <= (others => '0');   h113_out(d113_in'left downto 0) <= d113_in;  h113_en <= en_in;
   h114_out(h114_out'left downto d114_in'left + 1) <= (others => '0');   h114_out(d114_in'left downto 0) <= d114_in;  h114_en <= en_in;
   h115_out(h115_out'left downto d115_in'left + 1) <= (others => '0');   h115_out(d115_in'left downto 0) <= d115_in;  h115_en <= en_in;
   h116_out(h116_out'left downto d116_in'left + 1) <= (others => '0');   h116_out(d116_in'left downto 0) <= d116_in;  h116_en <= en_in;
   h117_out(h117_out'left downto d117_in'left + 1) <= (others => '0');   h117_out(d117_in'left downto 0) <= d117_in;  h117_en <= en_in;
   h118_out(h118_out'left downto d118_in'left + 1) <= (others => '0');   h118_out(d118_in'left downto 0) <= d118_in;  h118_en <= en_in;
   h119_out(h119_out'left downto d119_in'left + 1) <= (others => '0');   h119_out(d119_in'left downto 0) <= d119_in;  h119_en <= en_in;
   h120_out(h120_out'left downto d120_in'left + 1) <= (others => '0');   h120_out(d120_in'left downto 0) <= d120_in;  h120_en <= en_in;
   h121_out(h121_out'left downto d121_in'left + 1) <= (others => '0');   h121_out(d121_in'left downto 0) <= d121_in;  h121_en <= en_in;
   h122_out(h122_out'left downto d122_in'left + 1) <= (others => '0');   h122_out(d122_in'left downto 0) <= d122_in;  h122_en <= en_in;
   h123_out(h123_out'left downto d123_in'left + 1) <= (others => '0');   h123_out(d123_in'left downto 0) <= d123_in;  h123_en <= en_in;
   h124_out(h124_out'left downto d124_in'left + 1) <= (others => '0');   h124_out(d124_in'left downto 0) <= d124_in;  h124_en <= en_in;
   h125_out(h125_out'left downto d125_in'left + 1) <= (others => '0');   h125_out(d125_in'left downto 0) <= d125_in;  h125_en <= en_in;
   h126_out(h126_out'left downto d126_in'left + 1) <= (others => '0');   h126_out(d126_in'left downto 0) <= d126_in;  h126_en <= en_in;
   h127_out(h127_out'left downto d127_in'left + 1) <= (others => '0');   h127_out(d127_in'left downto 0) <= d127_in;  h127_en <= en_in;
   h128_out(h128_out'left downto d128_in'left + 1) <= (others => '0');   h128_out(d128_in'left downto 0) <= d128_in;  h128_en <= en_in;

   h129_out(h129_out'left downto d129_in'left + 1) <= (others => '0');   h129_out(d129_in'left downto 0) <= d129_in;   h129_en <= en_in;
   h130_out(h130_out'left downto d130_in'left + 1) <= (others => '0');   h130_out(d130_in'left downto 0) <= d130_in;   h130_en <= en_in;
   h131_out(h131_out'left downto d131_in'left + 1) <= (others => '0');   h131_out(d131_in'left downto 0) <= d131_in;   h131_en <= en_in;
   h132_out(h132_out'left downto d132_in'left + 1) <= (others => '0');   h132_out(d132_in'left downto 0) <= d132_in;   h132_en <= en_in;
   h133_out(h133_out'left downto d133_in'left + 1) <= (others => '0');   h133_out(d133_in'left downto 0) <= d133_in;   h133_en <= en_in;
   h134_out(h134_out'left downto d134_in'left + 1) <= (others => '0');   h134_out(d134_in'left downto 0) <= d134_in;   h134_en <= en_in;
   h135_out(h135_out'left downto d135_in'left + 1) <= (others => '0');   h135_out(d135_in'left downto 0) <= d135_in;   h135_en <= en_in;
   h136_out(h136_out'left downto d136_in'left + 1) <= (others => '0');   h136_out(d136_in'left downto 0) <= d136_in;   h136_en <= en_in;
   h137_out(h137_out'left downto d137_in'left + 1) <= (others => '0');   h137_out(d137_in'left downto 0) <= d137_in;   h137_en <= en_in;
   h138_out(h138_out'left downto d138_in'left + 1) <= (others => '0');   h138_out(d138_in'left downto 0) <= d138_in;   h138_en <= en_in;
   h139_out(h139_out'left downto d139_in'left + 1) <= (others => '0');   h139_out(d139_in'left downto 0) <= d139_in;   h139_en <= en_in;
   h140_out(h140_out'left downto d140_in'left + 1) <= (others => '0');   h140_out(d140_in'left downto 0) <= d140_in;   h140_en <= en_in;
   h141_out(h141_out'left downto d141_in'left + 1) <= (others => '0');   h141_out(d141_in'left downto 0) <= d141_in;   h141_en <= en_in;
   h142_out(h142_out'left downto d142_in'left + 1) <= (others => '0');   h142_out(d142_in'left downto 0) <= d142_in;   h142_en <= en_in;
   h143_out(h143_out'left downto d143_in'left + 1) <= (others => '0');   h143_out(d143_in'left downto 0) <= d143_in;   h143_en <= en_in;
   h144_out(h144_out'left downto d144_in'left + 1) <= (others => '0');   h144_out(d144_in'left downto 0) <= d144_in;   h144_en <= en_in;
   h145_out(h145_out'left downto d145_in'left + 1) <= (others => '0');   h145_out(d145_in'left downto 0) <= d145_in;   h145_en <= en_in;
   h146_out(h146_out'left downto d146_in'left + 1) <= (others => '0');   h146_out(d146_in'left downto 0) <= d146_in;   h146_en <= en_in;
   h147_out(h147_out'left downto d147_in'left + 1) <= (others => '0');   h147_out(d147_in'left downto 0) <= d147_in;   h147_en <= en_in;
   h148_out(h148_out'left downto d148_in'left + 1) <= (others => '0');   h148_out(d148_in'left downto 0) <= d148_in;   h148_en <= en_in;
   h149_out(h149_out'left downto d149_in'left + 1) <= (others => '0');   h149_out(d149_in'left downto 0) <= d149_in;   h149_en <= en_in;
   h150_out(h150_out'left downto d150_in'left + 1) <= (others => '0');   h150_out(d150_in'left downto 0) <= d150_in;   h150_en <= en_in;
   h151_out(h151_out'left downto d151_in'left + 1) <= (others => '0');   h151_out(d151_in'left downto 0) <= d151_in;   h151_en <= en_in;
   h152_out(h152_out'left downto d152_in'left + 1) <= (others => '0');   h152_out(d152_in'left downto 0) <= d152_in;   h152_en <= en_in;
   h153_out(h153_out'left downto d153_in'left + 1) <= (others => '0');   h153_out(d153_in'left downto 0) <= d153_in;   h153_en <= en_in;
   h154_out(h154_out'left downto d154_in'left + 1) <= (others => '0');   h154_out(d154_in'left downto 0) <= d154_in;   h154_en <= en_in;
   h155_out(h155_out'left downto d155_in'left + 1) <= (others => '0');   h155_out(d155_in'left downto 0) <= d155_in;   h155_en <= en_in;
   h156_out(h156_out'left downto d156_in'left + 1) <= (others => '0');   h156_out(d156_in'left downto 0) <= d156_in;   h156_en <= en_in;
   h157_out(h157_out'left downto d157_in'left + 1) <= (others => '0');   h157_out(d157_in'left downto 0) <= d157_in;   h157_en <= en_in;
   h158_out(h158_out'left downto d158_in'left + 1) <= (others => '0');   h158_out(d158_in'left downto 0) <= d158_in;   h158_en <= en_in;
   h159_out(h159_out'left downto d159_in'left + 1) <= (others => '0');   h159_out(d159_in'left downto 0) <= d159_in;   h159_en <= en_in;
   h160_out(h160_out'left downto d160_in'left + 1) <= (others => '0');   h160_out(d160_in'left downto 0) <= d160_in;   h160_en <= en_in;
   h161_out(h161_out'left downto d161_in'left + 1) <= (others => '0');   h161_out(d161_in'left downto 0) <= d161_in;   h161_en <= en_in;
   h162_out(h162_out'left downto d162_in'left + 1) <= (others => '0');   h162_out(d162_in'left downto 0) <= d162_in;   h162_en <= en_in;
   h163_out(h163_out'left downto d163_in'left + 1) <= (others => '0');   h163_out(d163_in'left downto 0) <= d163_in;   h163_en <= en_in;
   h164_out(h164_out'left downto d164_in'left + 1) <= (others => '0');   h164_out(d164_in'left downto 0) <= d164_in;   h164_en <= en_in;
   h165_out(h165_out'left downto d165_in'left + 1) <= (others => '0');   h165_out(d165_in'left downto 0) <= d165_in;   h165_en <= en_in;
   h166_out(h166_out'left downto d166_in'left + 1) <= (others => '0');   h166_out(d166_in'left downto 0) <= d166_in;   h166_en <= en_in;
   h167_out(h167_out'left downto d167_in'left + 1) <= (others => '0');   h167_out(d167_in'left downto 0) <= d167_in;   h167_en <= en_in;
   h168_out(h168_out'left downto d168_in'left + 1) <= (others => '0');   h168_out(d168_in'left downto 0) <= d168_in;   h168_en <= en_in;
   h169_out(h169_out'left downto d169_in'left + 1) <= (others => '0');   h169_out(d169_in'left downto 0) <= d169_in;   h169_en <= en_in;
   h170_out(h170_out'left downto d170_in'left + 1) <= (others => '0');   h170_out(d170_in'left downto 0) <= d170_in;   h170_en <= en_in;
   h171_out(h171_out'left downto d171_in'left + 1) <= (others => '0');   h171_out(d171_in'left downto 0) <= d171_in;   h171_en <= en_in;
   h172_out(h172_out'left downto d172_in'left + 1) <= (others => '0');   h172_out(d172_in'left downto 0) <= d172_in;   h172_en <= en_in;
   h173_out(h173_out'left downto d173_in'left + 1) <= (others => '0');   h173_out(d173_in'left downto 0) <= d173_in;   h173_en <= en_in;
   h174_out(h174_out'left downto d174_in'left + 1) <= (others => '0');   h174_out(d174_in'left downto 0) <= d174_in;   h174_en <= en_in;
   h175_out(h175_out'left downto d175_in'left + 1) <= (others => '0');   h175_out(d175_in'left downto 0) <= d175_in;   h175_en <= en_in;
   h176_out(h176_out'left downto d176_in'left + 1) <= (others => '0');   h176_out(d176_in'left downto 0) <= d176_in;   h176_en <= en_in;
   h177_out(h177_out'left downto d177_in'left + 1) <= (others => '0');   h177_out(d177_in'left downto 0) <= d177_in;   h177_en <= en_in;
   h178_out(h178_out'left downto d178_in'left + 1) <= (others => '0');   h178_out(d178_in'left downto 0) <= d178_in;   h178_en <= en_in;
   h179_out(h179_out'left downto d179_in'left + 1) <= (others => '0');   h179_out(d179_in'left downto 0) <= d179_in;   h179_en <= en_in;
   h180_out(h180_out'left downto d180_in'left + 1) <= (others => '0');   h180_out(d180_in'left downto 0) <= d180_in;   h180_en <= en_in;
   h181_out(h181_out'left downto d181_in'left + 1) <= (others => '0');   h181_out(d181_in'left downto 0) <= d181_in;   h181_en <= en_in;
   h182_out(h182_out'left downto d182_in'left + 1) <= (others => '0');   h182_out(d182_in'left downto 0) <= d182_in;   h182_en <= en_in;
   h183_out(h183_out'left downto d183_in'left + 1) <= (others => '0');   h183_out(d183_in'left downto 0) <= d183_in;   h183_en <= en_in;
   h184_out(h184_out'left downto d184_in'left + 1) <= (others => '0');   h184_out(d184_in'left downto 0) <= d184_in;   h184_en <= en_in;
   h185_out(h185_out'left downto d185_in'left + 1) <= (others => '0');   h185_out(d185_in'left downto 0) <= d185_in;   h185_en <= en_in;
   h186_out(h186_out'left downto d186_in'left + 1) <= (others => '0');   h186_out(d186_in'left downto 0) <= d186_in;   h186_en <= en_in;
   h187_out(h187_out'left downto d187_in'left + 1) <= (others => '0');   h187_out(d187_in'left downto 0) <= d187_in;   h187_en <= en_in;
   h188_out(h188_out'left downto d188_in'left + 1) <= (others => '0');   h188_out(d188_in'left downto 0) <= d188_in;   h188_en <= en_in;
   h189_out(h189_out'left downto d189_in'left + 1) <= (others => '0');   h189_out(d189_in'left downto 0) <= d189_in;   h189_en <= en_in;
   h190_out(h190_out'left downto d190_in'left + 1) <= (others => '0');   h190_out(d190_in'left downto 0) <= d190_in;   h190_en <= en_in;
   h191_out(h191_out'left downto d191_in'left + 1) <= (others => '0');   h191_out(d191_in'left downto 0) <= d191_in;   h191_en <= en_in;
   h192_out(h192_out'left downto d192_in'left + 1) <= (others => '0');   h192_out(d192_in'left downto 0) <= d192_in;   h192_en <= en_in;

   h193_out(h193_out'left downto d193_in'left + 1) <= (others => '0');   h193_out(d193_in'left downto 0) <= d193_in;   h193_en <= en_in;
   h194_out(h194_out'left downto d194_in'left + 1) <= (others => '0');   h194_out(d194_in'left downto 0) <= d194_in;   h194_en <= en_in;
   h195_out(h195_out'left downto d195_in'left + 1) <= (others => '0');   h195_out(d195_in'left downto 0) <= d195_in;   h195_en <= en_in;
   h196_out(h196_out'left downto d196_in'left + 1) <= (others => '0');   h196_out(d196_in'left downto 0) <= d196_in;   h196_en <= en_in;
   h197_out(h197_out'left downto d197_in'left + 1) <= (others => '0');   h197_out(d197_in'left downto 0) <= d197_in;   h197_en <= en_in;
   h198_out(h198_out'left downto d198_in'left + 1) <= (others => '0');   h198_out(d198_in'left downto 0) <= d198_in;   h198_en <= en_in;
   h199_out(h199_out'left downto d199_in'left + 1) <= (others => '0');   h199_out(d199_in'left downto 0) <= d199_in;   h199_en <= en_in;
   h200_out(h200_out'left downto d200_in'left + 1) <= (others => '0');   h200_out(d200_in'left downto 0) <= d200_in;   h200_en <= en_in;
   h201_out(h201_out'left downto d201_in'left + 1) <= (others => '0');   h201_out(d201_in'left downto 0) <= d201_in;   h201_en <= en_in;
   h202_out(h202_out'left downto d202_in'left + 1) <= (others => '0');   h202_out(d202_in'left downto 0) <= d202_in;   h202_en <= en_in;
   h203_out(h203_out'left downto d203_in'left + 1) <= (others => '0');   h203_out(d203_in'left downto 0) <= d203_in;   h203_en <= en_in;
   h204_out(h204_out'left downto d204_in'left + 1) <= (others => '0');   h204_out(d204_in'left downto 0) <= d204_in;   h204_en <= en_in;
   h205_out(h205_out'left downto d205_in'left + 1) <= (others => '0');   h205_out(d205_in'left downto 0) <= d205_in;   h205_en <= en_in;
   h206_out(h206_out'left downto d206_in'left + 1) <= (others => '0');   h206_out(d206_in'left downto 0) <= d206_in;   h206_en <= en_in;
   h207_out(h207_out'left downto d207_in'left + 1) <= (others => '0');   h207_out(d207_in'left downto 0) <= d207_in;   h207_en <= en_in;
   h208_out(h208_out'left downto d208_in'left + 1) <= (others => '0');   h208_out(d208_in'left downto 0) <= d208_in;   h208_en <= en_in;
   h209_out(h209_out'left downto d209_in'left + 1) <= (others => '0');   h209_out(d209_in'left downto 0) <= d209_in;   h209_en <= en_in;
   h210_out(h210_out'left downto d210_in'left + 1) <= (others => '0');   h210_out(d210_in'left downto 0) <= d210_in;   h210_en <= en_in;
   h211_out(h211_out'left downto d211_in'left + 1) <= (others => '0');   h211_out(d211_in'left downto 0) <= d211_in;   h211_en <= en_in;
   h212_out(h212_out'left downto d212_in'left + 1) <= (others => '0');   h212_out(d212_in'left downto 0) <= d212_in;   h212_en <= en_in;
   h213_out(h213_out'left downto d213_in'left + 1) <= (others => '0');   h213_out(d213_in'left downto 0) <= d213_in;   h213_en <= en_in;
   h214_out(h214_out'left downto d214_in'left + 1) <= (others => '0');   h214_out(d214_in'left downto 0) <= d214_in;   h214_en <= en_in;
   h215_out(h215_out'left downto d215_in'left + 1) <= (others => '0');   h215_out(d215_in'left downto 0) <= d215_in;   h215_en <= en_in;
   h216_out(h216_out'left downto d216_in'left + 1) <= (others => '0');   h216_out(d216_in'left downto 0) <= d216_in;   h216_en <= en_in;
   h217_out(h217_out'left downto d217_in'left + 1) <= (others => '0');   h217_out(d217_in'left downto 0) <= d217_in;   h217_en <= en_in;
   h218_out(h218_out'left downto d218_in'left + 1) <= (others => '0');   h218_out(d218_in'left downto 0) <= d218_in;   h218_en <= en_in;
   h219_out(h219_out'left downto d219_in'left + 1) <= (others => '0');   h219_out(d219_in'left downto 0) <= d219_in;   h219_en <= en_in;
   h220_out(h220_out'left downto d220_in'left + 1) <= (others => '0');   h220_out(d220_in'left downto 0) <= d220_in;   h220_en <= en_in;
   h221_out(h221_out'left downto d221_in'left + 1) <= (others => '0');   h221_out(d221_in'left downto 0) <= d221_in;   h221_en <= en_in;
   h222_out(h222_out'left downto d222_in'left + 1) <= (others => '0');   h222_out(d222_in'left downto 0) <= d222_in;   h222_en <= en_in;
   h223_out(h223_out'left downto d223_in'left + 1) <= (others => '0');   h223_out(d223_in'left downto 0) <= d223_in;   h223_en <= en_in;
   h224_out(h224_out'left downto d224_in'left + 1) <= (others => '0');   h224_out(d224_in'left downto 0) <= d224_in;   h224_en <= en_in;
   h225_out(h225_out'left downto d225_in'left + 1) <= (others => '0');   h225_out(d225_in'left downto 0) <= d225_in;   h225_en <= en_in;
   h226_out(h226_out'left downto d226_in'left + 1) <= (others => '0');   h226_out(d226_in'left downto 0) <= d226_in;   h226_en <= en_in;
   h227_out(h227_out'left downto d227_in'left + 1) <= (others => '0');   h227_out(d227_in'left downto 0) <= d227_in;   h227_en <= en_in;
   h228_out(h228_out'left downto d228_in'left + 1) <= (others => '0');   h228_out(d228_in'left downto 0) <= d228_in;   h228_en <= en_in;
   h229_out(h229_out'left downto d229_in'left + 1) <= (others => '0');   h229_out(d229_in'left downto 0) <= d229_in;   h229_en <= en_in;
   h230_out(h230_out'left downto d230_in'left + 1) <= (others => '0');   h230_out(d230_in'left downto 0) <= d230_in;   h230_en <= en_in;
   h231_out(h231_out'left downto d231_in'left + 1) <= (others => '0');   h231_out(d231_in'left downto 0) <= d231_in;   h231_en <= en_in;
   h232_out(h232_out'left downto d232_in'left + 1) <= (others => '0');   h232_out(d232_in'left downto 0) <= d232_in;   h232_en <= en_in;
   h233_out(h233_out'left downto d233_in'left + 1) <= (others => '0');   h233_out(d233_in'left downto 0) <= d233_in;   h233_en <= en_in;
   h234_out(h234_out'left downto d234_in'left + 1) <= (others => '0');   h234_out(d234_in'left downto 0) <= d234_in;   h234_en <= en_in;
   h235_out(h235_out'left downto d235_in'left + 1) <= (others => '0');   h235_out(d235_in'left downto 0) <= d235_in;   h235_en <= en_in;
   h236_out(h236_out'left downto d236_in'left + 1) <= (others => '0');   h236_out(d236_in'left downto 0) <= d236_in;   h236_en <= en_in;
   h237_out(h237_out'left downto d237_in'left + 1) <= (others => '0');   h237_out(d237_in'left downto 0) <= d237_in;   h237_en <= en_in;
   h238_out(h238_out'left downto d238_in'left + 1) <= (others => '0');   h238_out(d238_in'left downto 0) <= d238_in;   h238_en <= en_in;
   h239_out(h239_out'left downto d239_in'left + 1) <= (others => '0');   h239_out(d239_in'left downto 0) <= d239_in;   h239_en <= en_in;
   h240_out(h240_out'left downto d240_in'left + 1) <= (others => '0');   h240_out(d240_in'left downto 0) <= d240_in;   h240_en <= en_in;
   h241_out(h241_out'left downto d241_in'left + 1) <= (others => '0');   h241_out(d241_in'left downto 0) <= d241_in;   h241_en <= en_in;
   h242_out(h242_out'left downto d242_in'left + 1) <= (others => '0');   h242_out(d242_in'left downto 0) <= d242_in;   h242_en <= en_in;
   h243_out(h243_out'left downto d243_in'left + 1) <= (others => '0');   h243_out(d243_in'left downto 0) <= d243_in;   h243_en <= en_in;
   h244_out(h244_out'left downto d244_in'left + 1) <= (others => '0');   h244_out(d244_in'left downto 0) <= d244_in;   h244_en <= en_in;
   h245_out(h245_out'left downto d245_in'left + 1) <= (others => '0');   h245_out(d245_in'left downto 0) <= d245_in;   h245_en <= en_in;
   h246_out(h246_out'left downto d246_in'left + 1) <= (others => '0');   h246_out(d246_in'left downto 0) <= d246_in;   h246_en <= en_in;
   h247_out(h247_out'left downto d247_in'left + 1) <= (others => '0');   h247_out(d247_in'left downto 0) <= d247_in;   h247_en <= en_in;
   h248_out(h248_out'left downto d248_in'left + 1) <= (others => '0');   h248_out(d248_in'left downto 0) <= d248_in;   h248_en <= en_in;
   h249_out(h249_out'left downto d249_in'left + 1) <= (others => '0');   h249_out(d249_in'left downto 0) <= d249_in;   h249_en <= en_in;
   h250_out(h250_out'left downto d250_in'left + 1) <= (others => '0');   h250_out(d250_in'left downto 0) <= d250_in;   h250_en <= en_in;
   h251_out(h251_out'left downto d251_in'left + 1) <= (others => '0');   h251_out(d251_in'left downto 0) <= d251_in;   h251_en <= en_in;
   h252_out(h252_out'left downto d252_in'left + 1) <= (others => '0');   h252_out(d252_in'left downto 0) <= d252_in;   h252_en <= en_in;
   h253_out(h253_out'left downto d253_in'left + 1) <= (others => '0');   h253_out(d253_in'left downto 0) <= d253_in;   h253_en <= en_in;
   h254_out(h254_out'left downto d254_in'left + 1) <= (others => '0');   h254_out(d254_in'left downto 0) <= d254_in;   h254_en <= en_in;
   h255_out(h255_out'left downto d255_in'left + 1) <= (others => '0');   h255_out(d255_in'left downto 0) <= d255_in;   h255_en <= en_in;
   h256_out(h256_out'left downto d256_in'left + 1) <= (others => '0');   h256_out(d256_in'left downto 0) <= d256_in;   h256_en <= en_in;
end generate g_Huff_enc_dis;  
                                                                                                  
Buf01 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 0), enw=>h01_en, data_in=>h01_out, data_out=>buff01_out, burst_r=>en_out( 0), fifo_empty=> open, fifo_full=> open ); 
Buf02 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 1), enw=>h02_en, data_in=>h02_out, data_out=>buff02_out, burst_r=>en_out( 1), fifo_empty=> open, fifo_full=> open ); 
Buf03 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 2), enw=>h03_en, data_in=>h03_out, data_out=>buff03_out, burst_r=>en_out( 2), fifo_empty=> open, fifo_full=> open ); 
Buf04 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 3), enw=>h04_en, data_in=>h04_out, data_out=>buff04_out, burst_r=>en_out( 3), fifo_empty=> open, fifo_full=> open ); 
Buf05 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 4), enw=>h05_en, data_in=>h05_out, data_out=>buff05_out, burst_r=>en_out( 4), fifo_empty=> open, fifo_full=> open ); 
Buf06 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 5), enw=>h06_en, data_in=>h06_out, data_out=>buff06_out, burst_r=>en_out( 5), fifo_empty=> open, fifo_full=> open ); 
Buf07 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 6), enw=>h07_en, data_in=>h07_out, data_out=>buff07_out, burst_r=>en_out( 6), fifo_empty=> open, fifo_full=> open ); 
Buf08 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 7), enw=>h08_en, data_in=>h08_out, data_out=>buff08_out, burst_r=>en_out( 7), fifo_empty=> open, fifo_full=> open ); 
Buf09 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 8), enw=>h09_en, data_in=>h09_out, data_out=>buff09_out, burst_r=>en_out( 8), fifo_empty=> open, fifo_full=> open ); 
Buf10 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 9), enw=>h10_en, data_in=>h10_out, data_out=>buff10_out, burst_r=>en_out( 9), fifo_empty=> open, fifo_full=> open ); 
Buf11 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(10), enw=>h11_en, data_in=>h11_out, data_out=>buff11_out, burst_r=>en_out(10), fifo_empty=> open, fifo_full=> open ); 
Buf12 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(11), enw=>h12_en, data_in=>h12_out, data_out=>buff12_out, burst_r=>en_out(11), fifo_empty=> open, fifo_full=> open ); 
Buf13 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(12), enw=>h13_en, data_in=>h13_out, data_out=>buff13_out, burst_r=>en_out(12), fifo_empty=> open, fifo_full=> open ); 
Buf14 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(13), enw=>h14_en, data_in=>h14_out, data_out=>buff14_out, burst_r=>en_out(13), fifo_empty=> open, fifo_full=> open ); 
Buf15 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(14), enw=>h15_en, data_in=>h15_out, data_out=>buff15_out, burst_r=>en_out(14), fifo_empty=> open, fifo_full=> open ); 
Buf16 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(15), enw=>h16_en, data_in=>h16_out, data_out=>buff16_out, burst_r=>en_out(15), fifo_empty=> open, fifo_full=> open ); 
Buf17 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(16), enw=>h17_en, data_in=>h17_out, data_out=>buff17_out, burst_r=>en_out(16), fifo_empty=> open, fifo_full=> open ); 
Buf18 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(17), enw=>h18_en, data_in=>h18_out, data_out=>buff18_out, burst_r=>en_out(17), fifo_empty=> open, fifo_full=> open ); 
Buf19 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(18), enw=>h19_en, data_in=>h19_out, data_out=>buff19_out, burst_r=>en_out(18), fifo_empty=> open, fifo_full=> open ); 
Buf20 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(19), enw=>h20_en, data_in=>h20_out, data_out=>buff20_out, burst_r=>en_out(19), fifo_empty=> open, fifo_full=> open ); 
Buf21 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(20), enw=>h21_en, data_in=>h21_out, data_out=>buff21_out, burst_r=>en_out(20), fifo_empty=> open, fifo_full=> open ); 
Buf22 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(21), enw=>h22_en, data_in=>h22_out, data_out=>buff22_out, burst_r=>en_out(21), fifo_empty=> open, fifo_full=> open ); 
Buf23 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(22), enw=>h23_en, data_in=>h23_out, data_out=>buff23_out, burst_r=>en_out(22), fifo_empty=> open, fifo_full=> open ); 
Buf24 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(23), enw=>h24_en, data_in=>h24_out, data_out=>buff24_out, burst_r=>en_out(23), fifo_empty=> open, fifo_full=> open ); 
Buf25 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(24), enw=>h25_en, data_in=>h25_out, data_out=>buff25_out, burst_r=>en_out(24), fifo_empty=> open, fifo_full=> open ); 
Buf26 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(25), enw=>h26_en, data_in=>h26_out, data_out=>buff26_out, burst_r=>en_out(25), fifo_empty=> open, fifo_full=> open ); 
Buf27 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(26), enw=>h27_en, data_in=>h27_out, data_out=>buff27_out, burst_r=>en_out(26), fifo_empty=> open, fifo_full=> open ); 
Buf28 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(27), enw=>h28_en, data_in=>h28_out, data_out=>buff28_out, burst_r=>en_out(27), fifo_empty=> open, fifo_full=> open ); 
Buf29 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(28), enw=>h29_en, data_in=>h29_out, data_out=>buff29_out, burst_r=>en_out(28), fifo_empty=> open, fifo_full=> open ); 
Buf30 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(29), enw=>h30_en, data_in=>h30_out, data_out=>buff30_out, burst_r=>en_out(29), fifo_empty=> open, fifo_full=> open ); 
Buf31 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(30), enw=>h31_en, data_in=>h31_out, data_out=>buff31_out, burst_r=>en_out(30), fifo_empty=> open, fifo_full=> open ); 
Buf32 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(31), enw=>h32_en, data_in=>h32_out, data_out=>buff32_out, burst_r=>en_out(31), fifo_empty=> open, fifo_full=> open ); 
Buf33 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(32), enw=>h33_en, data_in=>h33_out, data_out=>buff33_out, burst_r=>en_out(32), fifo_empty=> open, fifo_full=> open ); 
Buf34 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(33), enw=>h34_en, data_in=>h34_out, data_out=>buff34_out, burst_r=>en_out(33), fifo_empty=> open, fifo_full=> open ); 
Buf35 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(34), enw=>h35_en, data_in=>h35_out, data_out=>buff35_out, burst_r=>en_out(34), fifo_empty=> open, fifo_full=> open ); 
Buf36 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(35), enw=>h36_en, data_in=>h36_out, data_out=>buff36_out, burst_r=>en_out(35), fifo_empty=> open, fifo_full=> open ); 
Buf37 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(36), enw=>h37_en, data_in=>h37_out, data_out=>buff37_out, burst_r=>en_out(36), fifo_empty=> open, fifo_full=> open ); 
Buf38 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(37), enw=>h38_en, data_in=>h38_out, data_out=>buff38_out, burst_r=>en_out(37), fifo_empty=> open, fifo_full=> open ); 
Buf39 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(38), enw=>h39_en, data_in=>h39_out, data_out=>buff39_out, burst_r=>en_out(38), fifo_empty=> open, fifo_full=> open ); 
Buf40 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(39), enw=>h40_en, data_in=>h40_out, data_out=>buff40_out, burst_r=>en_out(39), fifo_empty=> open, fifo_full=> open ); 
Buf41 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(40), enw=>h41_en, data_in=>h41_out, data_out=>buff41_out, burst_r=>en_out(40), fifo_empty=> open, fifo_full=> open ); 
Buf42 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(41), enw=>h42_en, data_in=>h42_out, data_out=>buff42_out, burst_r=>en_out(41), fifo_empty=> open, fifo_full=> open ); 
Buf43 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(42), enw=>h43_en, data_in=>h43_out, data_out=>buff43_out, burst_r=>en_out(42), fifo_empty=> open, fifo_full=> open ); 
Buf44 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(43), enw=>h44_en, data_in=>h44_out, data_out=>buff44_out, burst_r=>en_out(43), fifo_empty=> open, fifo_full=> open ); 
Buf45 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(44), enw=>h45_en, data_in=>h45_out, data_out=>buff45_out, burst_r=>en_out(44), fifo_empty=> open, fifo_full=> open ); 
Buf46 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(45), enw=>h46_en, data_in=>h46_out, data_out=>buff46_out, burst_r=>en_out(45), fifo_empty=> open, fifo_full=> open ); 
Buf47 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(46), enw=>h47_en, data_in=>h47_out, data_out=>buff47_out, burst_r=>en_out(46), fifo_empty=> open, fifo_full=> open ); 
Buf48 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(47), enw=>h48_en, data_in=>h48_out, data_out=>buff48_out, burst_r=>en_out(47), fifo_empty=> open, fifo_full=> open ); 
Buf49 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(48), enw=>h49_en, data_in=>h49_out, data_out=>buff49_out, burst_r=>en_out(48), fifo_empty=> open, fifo_full=> open ); 
Buf50 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(49), enw=>h50_en, data_in=>h50_out, data_out=>buff50_out, burst_r=>en_out(49), fifo_empty=> open, fifo_full=> open ); 
Buf51 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(50), enw=>h51_en, data_in=>h51_out, data_out=>buff51_out, burst_r=>en_out(50), fifo_empty=> open, fifo_full=> open ); 
Buf52 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(51), enw=>h52_en, data_in=>h52_out, data_out=>buff52_out, burst_r=>en_out(51), fifo_empty=> open, fifo_full=> open ); 
Buf53 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(52), enw=>h53_en, data_in=>h53_out, data_out=>buff53_out, burst_r=>en_out(52), fifo_empty=> open, fifo_full=> open ); 
Buf54 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(53), enw=>h54_en, data_in=>h54_out, data_out=>buff54_out, burst_r=>en_out(53), fifo_empty=> open, fifo_full=> open ); 
Buf55 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(54), enw=>h55_en, data_in=>h55_out, data_out=>buff55_out, burst_r=>en_out(54), fifo_empty=> open, fifo_full=> open ); 
Buf56 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(55), enw=>h56_en, data_in=>h56_out, data_out=>buff56_out, burst_r=>en_out(55), fifo_empty=> open, fifo_full=> open ); 
Buf57 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(56), enw=>h57_en, data_in=>h57_out, data_out=>buff57_out, burst_r=>en_out(56), fifo_empty=> open, fifo_full=> open ); 
Buf58 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(57), enw=>h58_en, data_in=>h58_out, data_out=>buff58_out, burst_r=>en_out(57), fifo_empty=> open, fifo_full=> open ); 
Buf59 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(58), enw=>h59_en, data_in=>h59_out, data_out=>buff59_out, burst_r=>en_out(58), fifo_empty=> open, fifo_full=> open ); 
Buf60 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(59), enw=>h60_en, data_in=>h60_out, data_out=>buff60_out, burst_r=>en_out(59), fifo_empty=> open, fifo_full=> open ); 
Buf61 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(60), enw=>h61_en, data_in=>h61_out, data_out=>buff61_out, burst_r=>en_out(60), fifo_empty=> open, fifo_full=> open ); 
Buf62 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(61), enw=>h62_en, data_in=>h62_out, data_out=>buff62_out, burst_r=>en_out(61), fifo_empty=> open, fifo_full=> open ); 
Buf63 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(62), enw=>h63_en, data_in=>h63_out, data_out=>buff63_out, burst_r=>en_out(62), fifo_empty=> open, fifo_full=> open ); 
Buf64 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(63), enw=>h64_en, data_in=>h64_out, data_out=>buff64_out, burst_r=>en_out(63), fifo_empty=> open, fifo_full=> open ); 

Buf65  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 64), enw=>h65_en , data_in=>h65_out , data_out=>buff65_out , burst_r=>en_out( 64), fifo_empty=> open, fifo_full=> open ); 
Buf66  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 65), enw=>h66_en , data_in=>h66_out , data_out=>buff66_out , burst_r=>en_out( 65), fifo_empty=> open, fifo_full=> open ); 
Buf67  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 66), enw=>h67_en , data_in=>h67_out , data_out=>buff67_out , burst_r=>en_out( 66), fifo_empty=> open, fifo_full=> open ); 
Buf68  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 67), enw=>h68_en , data_in=>h68_out , data_out=>buff68_out , burst_r=>en_out( 67), fifo_empty=> open, fifo_full=> open ); 
Buf69  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 68), enw=>h69_en , data_in=>h69_out , data_out=>buff69_out , burst_r=>en_out( 68), fifo_empty=> open, fifo_full=> open ); 
Buf70  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 69), enw=>h70_en , data_in=>h70_out , data_out=>buff70_out , burst_r=>en_out( 69), fifo_empty=> open, fifo_full=> open ); 
Buf71  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 70), enw=>h71_en , data_in=>h71_out , data_out=>buff71_out , burst_r=>en_out( 70), fifo_empty=> open, fifo_full=> open ); 
Buf72  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 71), enw=>h72_en , data_in=>h72_out , data_out=>buff72_out , burst_r=>en_out( 71), fifo_empty=> open, fifo_full=> open ); 
Buf73  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 72), enw=>h73_en , data_in=>h73_out , data_out=>buff73_out , burst_r=>en_out( 72), fifo_empty=> open, fifo_full=> open ); 
Buf74  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 73), enw=>h74_en , data_in=>h74_out , data_out=>buff74_out , burst_r=>en_out( 73), fifo_empty=> open, fifo_full=> open ); 
Buf75  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 74), enw=>h75_en , data_in=>h75_out , data_out=>buff75_out , burst_r=>en_out( 74), fifo_empty=> open, fifo_full=> open ); 
Buf76  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 75), enw=>h76_en , data_in=>h76_out , data_out=>buff76_out , burst_r=>en_out( 75), fifo_empty=> open, fifo_full=> open ); 
Buf77  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 76), enw=>h77_en , data_in=>h77_out , data_out=>buff77_out , burst_r=>en_out( 76), fifo_empty=> open, fifo_full=> open ); 
Buf78  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 77), enw=>h78_en , data_in=>h78_out , data_out=>buff78_out , burst_r=>en_out( 77), fifo_empty=> open, fifo_full=> open ); 
Buf79  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 78), enw=>h79_en , data_in=>h79_out , data_out=>buff79_out , burst_r=>en_out( 78), fifo_empty=> open, fifo_full=> open ); 
Buf80  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 79), enw=>h80_en , data_in=>h80_out , data_out=>buff80_out , burst_r=>en_out( 79), fifo_empty=> open, fifo_full=> open ); 
Buf81  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 80), enw=>h81_en , data_in=>h81_out , data_out=>buff81_out , burst_r=>en_out( 80), fifo_empty=> open, fifo_full=> open ); 
Buf82  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 81), enw=>h82_en , data_in=>h82_out , data_out=>buff82_out , burst_r=>en_out( 81), fifo_empty=> open, fifo_full=> open ); 
Buf83  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 82), enw=>h83_en , data_in=>h83_out , data_out=>buff83_out , burst_r=>en_out( 82), fifo_empty=> open, fifo_full=> open ); 
Buf84  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 83), enw=>h84_en , data_in=>h84_out , data_out=>buff84_out , burst_r=>en_out( 83), fifo_empty=> open, fifo_full=> open ); 
Buf85  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 84), enw=>h85_en , data_in=>h85_out , data_out=>buff85_out , burst_r=>en_out( 84), fifo_empty=> open, fifo_full=> open ); 
Buf86  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 85), enw=>h86_en , data_in=>h86_out , data_out=>buff86_out , burst_r=>en_out( 85), fifo_empty=> open, fifo_full=> open ); 
Buf87  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 86), enw=>h87_en , data_in=>h87_out , data_out=>buff87_out , burst_r=>en_out( 86), fifo_empty=> open, fifo_full=> open ); 
Buf88  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 87), enw=>h88_en , data_in=>h88_out , data_out=>buff88_out , burst_r=>en_out( 87), fifo_empty=> open, fifo_full=> open ); 
Buf89  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 88), enw=>h89_en , data_in=>h89_out , data_out=>buff89_out , burst_r=>en_out( 88), fifo_empty=> open, fifo_full=> open ); 
Buf90  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 89), enw=>h90_en , data_in=>h90_out , data_out=>buff90_out , burst_r=>en_out( 89), fifo_empty=> open, fifo_full=> open ); 
Buf91  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 90), enw=>h91_en , data_in=>h91_out , data_out=>buff91_out , burst_r=>en_out( 90), fifo_empty=> open, fifo_full=> open ); 
Buf92  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 91), enw=>h92_en , data_in=>h92_out , data_out=>buff92_out , burst_r=>en_out( 91), fifo_empty=> open, fifo_full=> open ); 
Buf93  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 92), enw=>h93_en , data_in=>h93_out , data_out=>buff93_out , burst_r=>en_out( 92), fifo_empty=> open, fifo_full=> open ); 
Buf94  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 93), enw=>h94_en , data_in=>h94_out , data_out=>buff94_out , burst_r=>en_out( 93), fifo_empty=> open, fifo_full=> open ); 
Buf95  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 94), enw=>h95_en , data_in=>h95_out , data_out=>buff95_out , burst_r=>en_out( 94), fifo_empty=> open, fifo_full=> open ); 
Buf96  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 95), enw=>h96_en , data_in=>h96_out , data_out=>buff96_out , burst_r=>en_out( 95), fifo_empty=> open, fifo_full=> open ); 
Buf97  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 96), enw=>h97_en , data_in=>h97_out , data_out=>buff97_out , burst_r=>en_out( 96), fifo_empty=> open, fifo_full=> open ); 
Buf98  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 97), enw=>h98_en , data_in=>h98_out , data_out=>buff98_out , burst_r=>en_out( 97), fifo_empty=> open, fifo_full=> open ); 
Buf99  : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 98), enw=>h99_en , data_in=>h99_out , data_out=>buff99_out , burst_r=>en_out( 98), fifo_empty=> open, fifo_full=> open ); 
Buf100 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd( 99), enw=>h100_en, data_in=>h100_out, data_out=>buff100_out, burst_r=>en_out( 99), fifo_empty=> open, fifo_full=> open ); 
Buf101 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(100), enw=>h101_en, data_in=>h101_out, data_out=>buff101_out, burst_r=>en_out(100), fifo_empty=> open, fifo_full=> open ); 
Buf102 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(101), enw=>h102_en, data_in=>h102_out, data_out=>buff102_out, burst_r=>en_out(101), fifo_empty=> open, fifo_full=> open ); 
Buf103 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(102), enw=>h103_en, data_in=>h103_out, data_out=>buff103_out, burst_r=>en_out(102), fifo_empty=> open, fifo_full=> open ); 
Buf104 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(103), enw=>h104_en, data_in=>h104_out, data_out=>buff104_out, burst_r=>en_out(103), fifo_empty=> open, fifo_full=> open ); 
Buf105 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(104), enw=>h105_en, data_in=>h105_out, data_out=>buff105_out, burst_r=>en_out(104), fifo_empty=> open, fifo_full=> open ); 
Buf106 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(105), enw=>h106_en, data_in=>h106_out, data_out=>buff106_out, burst_r=>en_out(105), fifo_empty=> open, fifo_full=> open ); 
Buf107 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(106), enw=>h107_en, data_in=>h107_out, data_out=>buff107_out, burst_r=>en_out(106), fifo_empty=> open, fifo_full=> open ); 
Buf108 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(107), enw=>h108_en, data_in=>h108_out, data_out=>buff108_out, burst_r=>en_out(107), fifo_empty=> open, fifo_full=> open ); 
Buf109 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(108), enw=>h109_en, data_in=>h109_out, data_out=>buff109_out, burst_r=>en_out(108), fifo_empty=> open, fifo_full=> open ); 
Buf110 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(109), enw=>h110_en, data_in=>h110_out, data_out=>buff110_out, burst_r=>en_out(109), fifo_empty=> open, fifo_full=> open ); 
Buf111 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(110), enw=>h111_en, data_in=>h111_out, data_out=>buff111_out, burst_r=>en_out(110), fifo_empty=> open, fifo_full=> open ); 
Buf112 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(111), enw=>h112_en, data_in=>h112_out, data_out=>buff112_out, burst_r=>en_out(111), fifo_empty=> open, fifo_full=> open ); 
Buf113 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(112), enw=>h113_en, data_in=>h113_out, data_out=>buff113_out, burst_r=>en_out(112), fifo_empty=> open, fifo_full=> open ); 
Buf114 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(113), enw=>h114_en, data_in=>h114_out, data_out=>buff114_out, burst_r=>en_out(113), fifo_empty=> open, fifo_full=> open ); 
Buf115 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(114), enw=>h115_en, data_in=>h115_out, data_out=>buff115_out, burst_r=>en_out(114), fifo_empty=> open, fifo_full=> open ); 
Buf116 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(115), enw=>h116_en, data_in=>h116_out, data_out=>buff116_out, burst_r=>en_out(115), fifo_empty=> open, fifo_full=> open ); 
Buf117 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(116), enw=>h117_en, data_in=>h117_out, data_out=>buff117_out, burst_r=>en_out(116), fifo_empty=> open, fifo_full=> open ); 
Buf118 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(117), enw=>h118_en, data_in=>h118_out, data_out=>buff118_out, burst_r=>en_out(117), fifo_empty=> open, fifo_full=> open ); 
Buf119 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(118), enw=>h119_en, data_in=>h119_out, data_out=>buff119_out, burst_r=>en_out(118), fifo_empty=> open, fifo_full=> open ); 
Buf120 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(119), enw=>h120_en, data_in=>h120_out, data_out=>buff120_out, burst_r=>en_out(119), fifo_empty=> open, fifo_full=> open ); 
Buf121 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(120), enw=>h121_en, data_in=>h121_out, data_out=>buff121_out, burst_r=>en_out(120), fifo_empty=> open, fifo_full=> open ); 
Buf122 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(121), enw=>h122_en, data_in=>h122_out, data_out=>buff122_out, burst_r=>en_out(121), fifo_empty=> open, fifo_full=> open ); 
Buf123 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(122), enw=>h123_en, data_in=>h123_out, data_out=>buff123_out, burst_r=>en_out(122), fifo_empty=> open, fifo_full=> open ); 
Buf124 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(123), enw=>h124_en, data_in=>h124_out, data_out=>buff124_out, burst_r=>en_out(123), fifo_empty=> open, fifo_full=> open ); 
Buf125 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(124), enw=>h125_en, data_in=>h125_out, data_out=>buff125_out, burst_r=>en_out(124), fifo_empty=> open, fifo_full=> open ); 
Buf126 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(125), enw=>h126_en, data_in=>h126_out, data_out=>buff126_out, burst_r=>en_out(125), fifo_empty=> open, fifo_full=> open ); 
Buf127 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(126), enw=>h127_en, data_in=>h127_out, data_out=>buff127_out, burst_r=>en_out(126), fifo_empty=> open, fifo_full=> open ); 
Buf128 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(127), enw=>h128_en, data_in=>h128_out, data_out=>buff128_out, burst_r=>en_out(127), fifo_empty=> open, fifo_full=> open ); 

Buf129 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(128), enw=>h129_en, data_in=>h129_out, data_out=>buff129_out, burst_r=>en_out(128), fifo_empty=> open, fifo_full=> open ); 
Buf130 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(129), enw=>h130_en, data_in=>h130_out, data_out=>buff130_out, burst_r=>en_out(129), fifo_empty=> open, fifo_full=> open ); 
Buf131 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(130), enw=>h131_en, data_in=>h131_out, data_out=>buff131_out, burst_r=>en_out(130), fifo_empty=> open, fifo_full=> open ); 
Buf132 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(131), enw=>h132_en, data_in=>h132_out, data_out=>buff132_out, burst_r=>en_out(131), fifo_empty=> open, fifo_full=> open ); 
Buf133 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(132), enw=>h133_en, data_in=>h133_out, data_out=>buff133_out, burst_r=>en_out(132), fifo_empty=> open, fifo_full=> open ); 
Buf134 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(133), enw=>h134_en, data_in=>h134_out, data_out=>buff134_out, burst_r=>en_out(133), fifo_empty=> open, fifo_full=> open ); 
Buf135 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(134), enw=>h135_en, data_in=>h135_out, data_out=>buff135_out, burst_r=>en_out(134), fifo_empty=> open, fifo_full=> open ); 
Buf136 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(135), enw=>h136_en, data_in=>h136_out, data_out=>buff136_out, burst_r=>en_out(135), fifo_empty=> open, fifo_full=> open ); 
Buf137 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(136), enw=>h137_en, data_in=>h137_out, data_out=>buff137_out, burst_r=>en_out(136), fifo_empty=> open, fifo_full=> open ); 
Buf138 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(137), enw=>h138_en, data_in=>h138_out, data_out=>buff138_out, burst_r=>en_out(137), fifo_empty=> open, fifo_full=> open ); 
Buf139 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(138), enw=>h139_en, data_in=>h139_out, data_out=>buff139_out, burst_r=>en_out(138), fifo_empty=> open, fifo_full=> open ); 
Buf140 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(139), enw=>h140_en, data_in=>h140_out, data_out=>buff140_out, burst_r=>en_out(139), fifo_empty=> open, fifo_full=> open ); 
Buf141 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(140), enw=>h141_en, data_in=>h141_out, data_out=>buff141_out, burst_r=>en_out(140), fifo_empty=> open, fifo_full=> open ); 
Buf142 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(141), enw=>h142_en, data_in=>h142_out, data_out=>buff142_out, burst_r=>en_out(141), fifo_empty=> open, fifo_full=> open ); 
Buf143 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(142), enw=>h143_en, data_in=>h143_out, data_out=>buff143_out, burst_r=>en_out(142), fifo_empty=> open, fifo_full=> open ); 
Buf144 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(143), enw=>h144_en, data_in=>h144_out, data_out=>buff144_out, burst_r=>en_out(143), fifo_empty=> open, fifo_full=> open ); 
Buf145 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(144), enw=>h145_en, data_in=>h145_out, data_out=>buff145_out, burst_r=>en_out(144), fifo_empty=> open, fifo_full=> open ); 
Buf146 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(145), enw=>h146_en, data_in=>h146_out, data_out=>buff146_out, burst_r=>en_out(145), fifo_empty=> open, fifo_full=> open ); 
Buf147 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(146), enw=>h147_en, data_in=>h147_out, data_out=>buff147_out, burst_r=>en_out(146), fifo_empty=> open, fifo_full=> open ); 
Buf148 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(147), enw=>h148_en, data_in=>h148_out, data_out=>buff148_out, burst_r=>en_out(147), fifo_empty=> open, fifo_full=> open ); 
Buf149 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(148), enw=>h149_en, data_in=>h149_out, data_out=>buff149_out, burst_r=>en_out(148), fifo_empty=> open, fifo_full=> open ); 
Buf150 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(149), enw=>h150_en, data_in=>h150_out, data_out=>buff150_out, burst_r=>en_out(149), fifo_empty=> open, fifo_full=> open ); 
Buf151 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(150), enw=>h151_en, data_in=>h151_out, data_out=>buff151_out, burst_r=>en_out(150), fifo_empty=> open, fifo_full=> open ); 
Buf152 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(151), enw=>h152_en, data_in=>h152_out, data_out=>buff152_out, burst_r=>en_out(151), fifo_empty=> open, fifo_full=> open ); 
Buf153 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(152), enw=>h153_en, data_in=>h153_out, data_out=>buff153_out, burst_r=>en_out(152), fifo_empty=> open, fifo_full=> open ); 
Buf154 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(153), enw=>h154_en, data_in=>h154_out, data_out=>buff154_out, burst_r=>en_out(153), fifo_empty=> open, fifo_full=> open ); 
Buf155 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(154), enw=>h155_en, data_in=>h155_out, data_out=>buff155_out, burst_r=>en_out(154), fifo_empty=> open, fifo_full=> open ); 
Buf156 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(155), enw=>h156_en, data_in=>h156_out, data_out=>buff156_out, burst_r=>en_out(155), fifo_empty=> open, fifo_full=> open ); 
Buf157 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(156), enw=>h157_en, data_in=>h157_out, data_out=>buff157_out, burst_r=>en_out(156), fifo_empty=> open, fifo_full=> open ); 
Buf158 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(157), enw=>h158_en, data_in=>h158_out, data_out=>buff158_out, burst_r=>en_out(157), fifo_empty=> open, fifo_full=> open ); 
Buf159 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(158), enw=>h159_en, data_in=>h159_out, data_out=>buff159_out, burst_r=>en_out(158), fifo_empty=> open, fifo_full=> open ); 
Buf160 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(159), enw=>h160_en, data_in=>h160_out, data_out=>buff160_out, burst_r=>en_out(159), fifo_empty=> open, fifo_full=> open ); 
Buf161 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(160), enw=>h161_en, data_in=>h161_out, data_out=>buff161_out, burst_r=>en_out(160), fifo_empty=> open, fifo_full=> open ); 
Buf162 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(161), enw=>h162_en, data_in=>h162_out, data_out=>buff162_out, burst_r=>en_out(161), fifo_empty=> open, fifo_full=> open ); 
Buf163 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(162), enw=>h163_en, data_in=>h163_out, data_out=>buff163_out, burst_r=>en_out(162), fifo_empty=> open, fifo_full=> open ); 
Buf164 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(163), enw=>h164_en, data_in=>h164_out, data_out=>buff164_out, burst_r=>en_out(163), fifo_empty=> open, fifo_full=> open ); 
Buf165 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(164), enw=>h165_en, data_in=>h165_out, data_out=>buff165_out, burst_r=>en_out(164), fifo_empty=> open, fifo_full=> open ); 
Buf166 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(165), enw=>h166_en, data_in=>h166_out, data_out=>buff166_out, burst_r=>en_out(165), fifo_empty=> open, fifo_full=> open ); 
Buf167 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(166), enw=>h167_en, data_in=>h167_out, data_out=>buff167_out, burst_r=>en_out(166), fifo_empty=> open, fifo_full=> open ); 
Buf168 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(167), enw=>h168_en, data_in=>h168_out, data_out=>buff168_out, burst_r=>en_out(167), fifo_empty=> open, fifo_full=> open ); 
Buf169 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(168), enw=>h169_en, data_in=>h169_out, data_out=>buff169_out, burst_r=>en_out(168), fifo_empty=> open, fifo_full=> open ); 
Buf170 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(169), enw=>h170_en, data_in=>h170_out, data_out=>buff170_out, burst_r=>en_out(169), fifo_empty=> open, fifo_full=> open ); 
Buf171 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(170), enw=>h171_en, data_in=>h171_out, data_out=>buff171_out, burst_r=>en_out(170), fifo_empty=> open, fifo_full=> open ); 
Buf172 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(171), enw=>h172_en, data_in=>h172_out, data_out=>buff172_out, burst_r=>en_out(171), fifo_empty=> open, fifo_full=> open ); 
Buf173 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(172), enw=>h173_en, data_in=>h173_out, data_out=>buff173_out, burst_r=>en_out(172), fifo_empty=> open, fifo_full=> open ); 
Buf174 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(173), enw=>h174_en, data_in=>h174_out, data_out=>buff174_out, burst_r=>en_out(173), fifo_empty=> open, fifo_full=> open ); 
Buf175 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(174), enw=>h175_en, data_in=>h175_out, data_out=>buff175_out, burst_r=>en_out(174), fifo_empty=> open, fifo_full=> open ); 
Buf176 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(175), enw=>h176_en, data_in=>h176_out, data_out=>buff176_out, burst_r=>en_out(175), fifo_empty=> open, fifo_full=> open ); 
Buf177 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(176), enw=>h177_en, data_in=>h177_out, data_out=>buff177_out, burst_r=>en_out(176), fifo_empty=> open, fifo_full=> open ); 
Buf178 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(177), enw=>h178_en, data_in=>h178_out, data_out=>buff178_out, burst_r=>en_out(177), fifo_empty=> open, fifo_full=> open ); 
Buf179 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(178), enw=>h179_en, data_in=>h179_out, data_out=>buff179_out, burst_r=>en_out(178), fifo_empty=> open, fifo_full=> open ); 
Buf180 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(179), enw=>h180_en, data_in=>h180_out, data_out=>buff180_out, burst_r=>en_out(179), fifo_empty=> open, fifo_full=> open ); 
Buf181 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(180), enw=>h181_en, data_in=>h181_out, data_out=>buff181_out, burst_r=>en_out(180), fifo_empty=> open, fifo_full=> open ); 
Buf182 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(181), enw=>h182_en, data_in=>h182_out, data_out=>buff182_out, burst_r=>en_out(181), fifo_empty=> open, fifo_full=> open ); 
Buf183 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(182), enw=>h183_en, data_in=>h183_out, data_out=>buff183_out, burst_r=>en_out(182), fifo_empty=> open, fifo_full=> open ); 
Buf184 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(183), enw=>h184_en, data_in=>h184_out, data_out=>buff184_out, burst_r=>en_out(183), fifo_empty=> open, fifo_full=> open ); 
Buf185 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(184), enw=>h185_en, data_in=>h185_out, data_out=>buff185_out, burst_r=>en_out(184), fifo_empty=> open, fifo_full=> open ); 
Buf186 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(185), enw=>h186_en, data_in=>h186_out, data_out=>buff186_out, burst_r=>en_out(185), fifo_empty=> open, fifo_full=> open ); 
Buf187 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(186), enw=>h187_en, data_in=>h187_out, data_out=>buff187_out, burst_r=>en_out(186), fifo_empty=> open, fifo_full=> open ); 
Buf188 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(187), enw=>h188_en, data_in=>h188_out, data_out=>buff188_out, burst_r=>en_out(187), fifo_empty=> open, fifo_full=> open ); 
Buf189 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(188), enw=>h189_en, data_in=>h189_out, data_out=>buff189_out, burst_r=>en_out(188), fifo_empty=> open, fifo_full=> open ); 
Buf190 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(189), enw=>h190_en, data_in=>h190_out, data_out=>buff190_out, burst_r=>en_out(189), fifo_empty=> open, fifo_full=> open ); 
Buf191 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(190), enw=>h191_en, data_in=>h191_out, data_out=>buff191_out, burst_r=>en_out(190), fifo_empty=> open, fifo_full=> open ); 
Buf192 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(191), enw=>h192_en, data_in=>h192_out, data_out=>buff192_out, burst_r=>en_out(191), fifo_empty=> open, fifo_full=> open ); 

Buf193 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(192), enw=>h193_en, data_in=>h193_out, data_out=>buff193_out, burst_r=>en_out(192), fifo_empty=> open, fifo_full=> open ); 
Buf194 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(193), enw=>h194_en, data_in=>h194_out, data_out=>buff194_out, burst_r=>en_out(193), fifo_empty=> open, fifo_full=> open ); 
Buf195 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(194), enw=>h195_en, data_in=>h195_out, data_out=>buff195_out, burst_r=>en_out(194), fifo_empty=> open, fifo_full=> open ); 
Buf196 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(195), enw=>h196_en, data_in=>h196_out, data_out=>buff196_out, burst_r=>en_out(195), fifo_empty=> open, fifo_full=> open ); 
Buf197 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(196), enw=>h197_en, data_in=>h197_out, data_out=>buff197_out, burst_r=>en_out(196), fifo_empty=> open, fifo_full=> open ); 
Buf198 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(197), enw=>h198_en, data_in=>h198_out, data_out=>buff198_out, burst_r=>en_out(197), fifo_empty=> open, fifo_full=> open ); 
Buf199 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(198), enw=>h199_en, data_in=>h199_out, data_out=>buff199_out, burst_r=>en_out(198), fifo_empty=> open, fifo_full=> open ); 
Buf200 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(199), enw=>h200_en, data_in=>h200_out, data_out=>buff200_out, burst_r=>en_out(199), fifo_empty=> open, fifo_full=> open ); 
Buf201 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(200), enw=>h201_en, data_in=>h201_out, data_out=>buff201_out, burst_r=>en_out(200), fifo_empty=> open, fifo_full=> open ); 
Buf202 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(201), enw=>h202_en, data_in=>h202_out, data_out=>buff202_out, burst_r=>en_out(201), fifo_empty=> open, fifo_full=> open ); 
Buf203 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(202), enw=>h203_en, data_in=>h203_out, data_out=>buff203_out, burst_r=>en_out(202), fifo_empty=> open, fifo_full=> open ); 
Buf204 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(203), enw=>h204_en, data_in=>h204_out, data_out=>buff204_out, burst_r=>en_out(203), fifo_empty=> open, fifo_full=> open ); 
Buf205 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(204), enw=>h205_en, data_in=>h205_out, data_out=>buff205_out, burst_r=>en_out(204), fifo_empty=> open, fifo_full=> open ); 
Buf206 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(205), enw=>h206_en, data_in=>h206_out, data_out=>buff206_out, burst_r=>en_out(205), fifo_empty=> open, fifo_full=> open ); 
Buf207 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(206), enw=>h207_en, data_in=>h207_out, data_out=>buff207_out, burst_r=>en_out(206), fifo_empty=> open, fifo_full=> open ); 
Buf208 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(207), enw=>h208_en, data_in=>h208_out, data_out=>buff208_out, burst_r=>en_out(207), fifo_empty=> open, fifo_full=> open ); 
Buf209 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(208), enw=>h209_en, data_in=>h209_out, data_out=>buff209_out, burst_r=>en_out(208), fifo_empty=> open, fifo_full=> open ); 
Buf210 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(209), enw=>h210_en, data_in=>h210_out, data_out=>buff210_out, burst_r=>en_out(209), fifo_empty=> open, fifo_full=> open ); 
Buf211 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(210), enw=>h211_en, data_in=>h211_out, data_out=>buff211_out, burst_r=>en_out(210), fifo_empty=> open, fifo_full=> open ); 
Buf212 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(211), enw=>h212_en, data_in=>h212_out, data_out=>buff212_out, burst_r=>en_out(211), fifo_empty=> open, fifo_full=> open ); 
Buf213 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(212), enw=>h213_en, data_in=>h213_out, data_out=>buff213_out, burst_r=>en_out(212), fifo_empty=> open, fifo_full=> open ); 
Buf214 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(213), enw=>h214_en, data_in=>h214_out, data_out=>buff214_out, burst_r=>en_out(213), fifo_empty=> open, fifo_full=> open ); 
Buf215 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(214), enw=>h215_en, data_in=>h215_out, data_out=>buff215_out, burst_r=>en_out(214), fifo_empty=> open, fifo_full=> open ); 
Buf216 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(215), enw=>h216_en, data_in=>h216_out, data_out=>buff216_out, burst_r=>en_out(215), fifo_empty=> open, fifo_full=> open ); 
Buf217 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(216), enw=>h217_en, data_in=>h217_out, data_out=>buff217_out, burst_r=>en_out(216), fifo_empty=> open, fifo_full=> open ); 
Buf218 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(217), enw=>h218_en, data_in=>h218_out, data_out=>buff218_out, burst_r=>en_out(217), fifo_empty=> open, fifo_full=> open ); 
Buf219 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(218), enw=>h219_en, data_in=>h219_out, data_out=>buff219_out, burst_r=>en_out(218), fifo_empty=> open, fifo_full=> open ); 
Buf220 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(219), enw=>h220_en, data_in=>h220_out, data_out=>buff220_out, burst_r=>en_out(219), fifo_empty=> open, fifo_full=> open ); 
Buf221 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(220), enw=>h221_en, data_in=>h221_out, data_out=>buff221_out, burst_r=>en_out(220), fifo_empty=> open, fifo_full=> open ); 
Buf222 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(221), enw=>h222_en, data_in=>h222_out, data_out=>buff222_out, burst_r=>en_out(221), fifo_empty=> open, fifo_full=> open ); 
Buf223 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(222), enw=>h223_en, data_in=>h223_out, data_out=>buff223_out, burst_r=>en_out(222), fifo_empty=> open, fifo_full=> open ); 
Buf224 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(223), enw=>h224_en, data_in=>h224_out, data_out=>buff224_out, burst_r=>en_out(223), fifo_empty=> open, fifo_full=> open ); 
Buf225 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(224), enw=>h225_en, data_in=>h225_out, data_out=>buff225_out, burst_r=>en_out(224), fifo_empty=> open, fifo_full=> open ); 
Buf226 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(225), enw=>h226_en, data_in=>h226_out, data_out=>buff226_out, burst_r=>en_out(225), fifo_empty=> open, fifo_full=> open ); 
Buf227 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(226), enw=>h227_en, data_in=>h227_out, data_out=>buff227_out, burst_r=>en_out(226), fifo_empty=> open, fifo_full=> open ); 
Buf228 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(227), enw=>h228_en, data_in=>h228_out, data_out=>buff228_out, burst_r=>en_out(227), fifo_empty=> open, fifo_full=> open ); 
Buf229 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(228), enw=>h229_en, data_in=>h229_out, data_out=>buff229_out, burst_r=>en_out(228), fifo_empty=> open, fifo_full=> open ); 
Buf230 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(229), enw=>h230_en, data_in=>h230_out, data_out=>buff230_out, burst_r=>en_out(229), fifo_empty=> open, fifo_full=> open ); 
Buf231 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(230), enw=>h231_en, data_in=>h231_out, data_out=>buff231_out, burst_r=>en_out(230), fifo_empty=> open, fifo_full=> open ); 
Buf232 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(231), enw=>h232_en, data_in=>h232_out, data_out=>buff232_out, burst_r=>en_out(231), fifo_empty=> open, fifo_full=> open ); 
Buf233 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(232), enw=>h233_en, data_in=>h233_out, data_out=>buff233_out, burst_r=>en_out(232), fifo_empty=> open, fifo_full=> open ); 
Buf234 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(233), enw=>h234_en, data_in=>h234_out, data_out=>buff234_out, burst_r=>en_out(233), fifo_empty=> open, fifo_full=> open ); 
Buf235 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(234), enw=>h235_en, data_in=>h235_out, data_out=>buff235_out, burst_r=>en_out(234), fifo_empty=> open, fifo_full=> open ); 
Buf236 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(235), enw=>h236_en, data_in=>h236_out, data_out=>buff236_out, burst_r=>en_out(235), fifo_empty=> open, fifo_full=> open ); 
Buf237 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(236), enw=>h237_en, data_in=>h237_out, data_out=>buff237_out, burst_r=>en_out(236), fifo_empty=> open, fifo_full=> open ); 
Buf238 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(237), enw=>h238_en, data_in=>h238_out, data_out=>buff238_out, burst_r=>en_out(237), fifo_empty=> open, fifo_full=> open ); 
Buf239 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(238), enw=>h239_en, data_in=>h239_out, data_out=>buff239_out, burst_r=>en_out(238), fifo_empty=> open, fifo_full=> open ); 
Buf240 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(239), enw=>h240_en, data_in=>h240_out, data_out=>buff240_out, burst_r=>en_out(239), fifo_empty=> open, fifo_full=> open ); 
Buf241 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(240), enw=>h241_en, data_in=>h241_out, data_out=>buff241_out, burst_r=>en_out(240), fifo_empty=> open, fifo_full=> open ); 
Buf242 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(241), enw=>h242_en, data_in=>h242_out, data_out=>buff242_out, burst_r=>en_out(241), fifo_empty=> open, fifo_full=> open ); 
Buf243 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(242), enw=>h243_en, data_in=>h243_out, data_out=>buff243_out, burst_r=>en_out(242), fifo_empty=> open, fifo_full=> open ); 
Buf244 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(243), enw=>h244_en, data_in=>h244_out, data_out=>buff244_out, burst_r=>en_out(243), fifo_empty=> open, fifo_full=> open ); 
Buf245 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(244), enw=>h245_en, data_in=>h245_out, data_out=>buff245_out, burst_r=>en_out(244), fifo_empty=> open, fifo_full=> open ); 
Buf246 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(245), enw=>h246_en, data_in=>h246_out, data_out=>buff246_out, burst_r=>en_out(245), fifo_empty=> open, fifo_full=> open ); 
Buf247 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(246), enw=>h247_en, data_in=>h247_out, data_out=>buff247_out, burst_r=>en_out(246), fifo_empty=> open, fifo_full=> open ); 
Buf248 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(247), enw=>h248_en, data_in=>h248_out, data_out=>buff248_out, burst_r=>en_out(247), fifo_empty=> open, fifo_full=> open ); 
Buf249 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(248), enw=>h249_en, data_in=>h249_out, data_out=>buff249_out, burst_r=>en_out(248), fifo_empty=> open, fifo_full=> open ); 
Buf250 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(249), enw=>h250_en, data_in=>h250_out, data_out=>buff250_out, burst_r=>en_out(249), fifo_empty=> open, fifo_full=> open ); 
Buf251 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(250), enw=>h251_en, data_in=>h251_out, data_out=>buff251_out, burst_r=>en_out(250), fifo_empty=> open, fifo_full=> open ); 
Buf252 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(251), enw=>h252_en, data_in=>h252_out, data_out=>buff252_out, burst_r=>en_out(251), fifo_empty=> open, fifo_full=> open ); 
Buf253 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(252), enw=>h253_en, data_in=>h253_out, data_out=>buff253_out, burst_r=>en_out(252), fifo_empty=> open, fifo_full=> open ); 
Buf254 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(253), enw=>h254_en, data_in=>h254_out, data_out=>buff254_out, burst_r=>en_out(253), fifo_empty=> open, fifo_full=> open ); 
Buf255 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(254), enw=>h255_en, data_in=>h255_out, data_out=>buff255_out, burst_r=>en_out(254), fifo_empty=> open, fifo_full=> open ); 
Buf256 : fifo generic map(depth=>depth, burst=>burst, Win=>Wh, Wout=>Wb) port map(clk =>clk, rst =>rst, enr =>b_rd(255), enw=>h256_en, data_in=>h256_out, data_out=>buff256_out, burst_r=>en_out(255), fifo_empty=> open, fifo_full=> open ); 
--b_rd <= x"0000000000000001"; -- one Huffman
--d_out <= buff01_out;         -- one Huffman
p_rd_ctr :     process (clk, rst)
begin
   if ( rst = '1') then
      b_rd <= conv_std_logic_vector(0, b_rd'length);
   elsif(rising_edge(clk)) then   
      if buf_rd = '1' then
         --case
         if conv_integer('0' & buf_num) =    0 then b_rd <= x"0000000000000000000000000000000000000000000000000000000000000001"; end if;
         if conv_integer('0' & buf_num) =    1 then b_rd <= x"0000000000000000000000000000000000000000000000000000000000000002"; end if;
         if conv_integer('0' & buf_num) =    2 then b_rd <= x"0000000000000000000000000000000000000000000000000000000000000004"; end if;
         if conv_integer('0' & buf_num) =    3 then b_rd <= x"0000000000000000000000000000000000000000000000000000000000000008"; end if;
         if conv_integer('0' & buf_num) =    4 then b_rd <= x"0000000000000000000000000000000000000000000000000000000000000010"; end if;
         if conv_integer('0' & buf_num) =    5 then b_rd <= x"0000000000000000000000000000000000000000000000000000000000000020"; end if;
         if conv_integer('0' & buf_num) =    6 then b_rd <= x"0000000000000000000000000000000000000000000000000000000000000040"; end if;
         if conv_integer('0' & buf_num) =    7 then b_rd <= x"0000000000000000000000000000000000000000000000000000000000000080"; end if;
         if conv_integer('0' & buf_num) =    8 then b_rd <= x"0000000000000000000000000000000000000000000000000000000000000100"; end if;
         if conv_integer('0' & buf_num) =    9 then b_rd <= x"0000000000000000000000000000000000000000000000000000000000000200"; end if;
         if conv_integer('0' & buf_num) =   10 then b_rd <= x"0000000000000000000000000000000000000000000000000000000000000400"; end if;
         if conv_integer('0' & buf_num) =   11 then b_rd <= x"0000000000000000000000000000000000000000000000000000000000000800"; end if;
         if conv_integer('0' & buf_num) =   12 then b_rd <= x"0000000000000000000000000000000000000000000000000000000000001000"; end if;
         if conv_integer('0' & buf_num) =   13 then b_rd <= x"0000000000000000000000000000000000000000000000000000000000002000"; end if;
         if conv_integer('0' & buf_num) =   14 then b_rd <= x"0000000000000000000000000000000000000000000000000000000000004000"; end if;
         if conv_integer('0' & buf_num) =   15 then b_rd <= x"0000000000000000000000000000000000000000000000000000000000008000"; end if;
         if conv_integer('0' & buf_num) =   16 then b_rd <= x"0000000000000000000000000000000000000000000000000000000000010000"; end if;
         if conv_integer('0' & buf_num) =   17 then b_rd <= x"0000000000000000000000000000000000000000000000000000000000020000"; end if;
         if conv_integer('0' & buf_num) =   18 then b_rd <= x"0000000000000000000000000000000000000000000000000000000000040000"; end if;
         if conv_integer('0' & buf_num) =   19 then b_rd <= x"0000000000000000000000000000000000000000000000000000000000080000"; end if;
         if conv_integer('0' & buf_num) =   20 then b_rd <= x"0000000000000000000000000000000000000000000000000000000000100000"; end if;
         if conv_integer('0' & buf_num) =   21 then b_rd <= x"0000000000000000000000000000000000000000000000000000000000200000"; end if;
         if conv_integer('0' & buf_num) =   22 then b_rd <= x"0000000000000000000000000000000000000000000000000000000000400000"; end if;
         if conv_integer('0' & buf_num) =   23 then b_rd <= x"0000000000000000000000000000000000000000000000000000000000800000"; end if;
         if conv_integer('0' & buf_num) =   24 then b_rd <= x"0000000000000000000000000000000000000000000000000000000001000000"; end if;
         if conv_integer('0' & buf_num) =   25 then b_rd <= x"0000000000000000000000000000000000000000000000000000000002000000"; end if;
         if conv_integer('0' & buf_num) =   26 then b_rd <= x"0000000000000000000000000000000000000000000000000000000004000000"; end if;
         if conv_integer('0' & buf_num) =   27 then b_rd <= x"0000000000000000000000000000000000000000000000000000000008000000"; end if;
         if conv_integer('0' & buf_num) =   28 then b_rd <= x"0000000000000000000000000000000000000000000000000000000010000000"; end if;
         if conv_integer('0' & buf_num) =   29 then b_rd <= x"0000000000000000000000000000000000000000000000000000000020000000"; end if;
         if conv_integer('0' & buf_num) =   30 then b_rd <= x"0000000000000000000000000000000000000000000000000000000040000000"; end if;
         if conv_integer('0' & buf_num) =   31 then b_rd <= x"0000000000000000000000000000000000000000000000000000000080000000"; end if;
         if conv_integer('0' & buf_num) =   32 then b_rd <= x"0000000000000000000000000000000000000000000000000000000100000000"; end if;
         if conv_integer('0' & buf_num) =   33 then b_rd <= x"0000000000000000000000000000000000000000000000000000000200000000"; end if;
         if conv_integer('0' & buf_num) =   34 then b_rd <= x"0000000000000000000000000000000000000000000000000000000400000000"; end if;
         if conv_integer('0' & buf_num) =   35 then b_rd <= x"0000000000000000000000000000000000000000000000000000000800000000"; end if;
         if conv_integer('0' & buf_num) =   36 then b_rd <= x"0000000000000000000000000000000000000000000000000000001000000000"; end if;
         if conv_integer('0' & buf_num) =   37 then b_rd <= x"0000000000000000000000000000000000000000000000000000002000000000"; end if;
         if conv_integer('0' & buf_num) =   38 then b_rd <= x"0000000000000000000000000000000000000000000000000000004000000000"; end if;
         if conv_integer('0' & buf_num) =   39 then b_rd <= x"0000000000000000000000000000000000000000000000000000008000000000"; end if;
         if conv_integer('0' & buf_num) =   40 then b_rd <= x"0000000000000000000000000000000000000000000000000000010000000000"; end if;
         if conv_integer('0' & buf_num) =   41 then b_rd <= x"0000000000000000000000000000000000000000000000000000020000000000"; end if;
         if conv_integer('0' & buf_num) =   42 then b_rd <= x"0000000000000000000000000000000000000000000000000000040000000000"; end if;
         if conv_integer('0' & buf_num) =   43 then b_rd <= x"0000000000000000000000000000000000000000000000000000080000000000"; end if;
         if conv_integer('0' & buf_num) =   44 then b_rd <= x"0000000000000000000000000000000000000000000000000000100000000000"; end if;
         if conv_integer('0' & buf_num) =   45 then b_rd <= x"0000000000000000000000000000000000000000000000000000200000000000"; end if;
         if conv_integer('0' & buf_num) =   46 then b_rd <= x"0000000000000000000000000000000000000000000000000000400000000000"; end if;
         if conv_integer('0' & buf_num) =   47 then b_rd <= x"0000000000000000000000000000000000000000000000000000800000000000"; end if;
         if conv_integer('0' & buf_num) =   48 then b_rd <= x"0000000000000000000000000000000000000000000000000001000000000000"; end if;
         if conv_integer('0' & buf_num) =   49 then b_rd <= x"0000000000000000000000000000000000000000000000000002000000000000"; end if;
         if conv_integer('0' & buf_num) =   50 then b_rd <= x"0000000000000000000000000000000000000000000000000004000000000000"; end if;
         if conv_integer('0' & buf_num) =   51 then b_rd <= x"0000000000000000000000000000000000000000000000000008000000000000"; end if;
         if conv_integer('0' & buf_num) =   52 then b_rd <= x"0000000000000000000000000000000000000000000000000010000000000000"; end if;
         if conv_integer('0' & buf_num) =   53 then b_rd <= x"0000000000000000000000000000000000000000000000000020000000000000"; end if;
         if conv_integer('0' & buf_num) =   54 then b_rd <= x"0000000000000000000000000000000000000000000000000040000000000000"; end if;
         if conv_integer('0' & buf_num) =   55 then b_rd <= x"0000000000000000000000000000000000000000000000000080000000000000"; end if;
         if conv_integer('0' & buf_num) =   56 then b_rd <= x"0000000000000000000000000000000000000000000000000100000000000000"; end if;
         if conv_integer('0' & buf_num) =   57 then b_rd <= x"0000000000000000000000000000000000000000000000000200000000000000"; end if;
         if conv_integer('0' & buf_num) =   58 then b_rd <= x"0000000000000000000000000000000000000000000000000400000000000000"; end if;
         if conv_integer('0' & buf_num) =   59 then b_rd <= x"0000000000000000000000000000000000000000000000000800000000000000"; end if;
         if conv_integer('0' & buf_num) =   60 then b_rd <= x"0000000000000000000000000000000000000000000000001000000000000000"; end if;
         if conv_integer('0' & buf_num) =   61 then b_rd <= x"0000000000000000000000000000000000000000000000002000000000000000"; end if;
         if conv_integer('0' & buf_num) =   62 then b_rd <= x"0000000000000000000000000000000000000000000000004000000000000000"; end if;
         if conv_integer('0' & buf_num) =   63 then b_rd <= x"0000000000000000000000000000000000000000000000008000000000000000"; end if;

         if conv_integer('0' & buf_num) =   64  then b_rd <= x"0000000000000000000000000000000000000000000000010000000000000000"; end if;
         if conv_integer('0' & buf_num) =   65  then b_rd <= x"0000000000000000000000000000000000000000000000020000000000000000"; end if;
         if conv_integer('0' & buf_num) =   66  then b_rd <= x"0000000000000000000000000000000000000000000000040000000000000000"; end if;
         if conv_integer('0' & buf_num) =   67  then b_rd <= x"0000000000000000000000000000000000000000000000080000000000000000"; end if;
         if conv_integer('0' & buf_num) =   68  then b_rd <= x"0000000000000000000000000000000000000000000000100000000000000000"; end if;
         if conv_integer('0' & buf_num) =   69  then b_rd <= x"0000000000000000000000000000000000000000000000200000000000000000"; end if;
         if conv_integer('0' & buf_num) =   70  then b_rd <= x"0000000000000000000000000000000000000000000000400000000000000000"; end if;
         if conv_integer('0' & buf_num) =   71  then b_rd <= x"0000000000000000000000000000000000000000000000800000000000000000"; end if;
         if conv_integer('0' & buf_num) =   72  then b_rd <= x"0000000000000000000000000000000000000000000001000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   73  then b_rd <= x"0000000000000000000000000000000000000000000002000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   74  then b_rd <= x"0000000000000000000000000000000000000000000004000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   75  then b_rd <= x"0000000000000000000000000000000000000000000008000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   76  then b_rd <= x"0000000000000000000000000000000000000000000010000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   77  then b_rd <= x"0000000000000000000000000000000000000000000020000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   78  then b_rd <= x"0000000000000000000000000000000000000000000040000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   79  then b_rd <= x"0000000000000000000000000000000000000000000080000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   80  then b_rd <= x"0000000000000000000000000000000000000000000100000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   81  then b_rd <= x"0000000000000000000000000000000000000000000200000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   82  then b_rd <= x"0000000000000000000000000000000000000000000400000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   83  then b_rd <= x"0000000000000000000000000000000000000000000800000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   84  then b_rd <= x"0000000000000000000000000000000000000000001000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   85  then b_rd <= x"0000000000000000000000000000000000000000002000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   86  then b_rd <= x"0000000000000000000000000000000000000000004000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   87  then b_rd <= x"0000000000000000000000000000000000000000008000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   88  then b_rd <= x"0000000000000000000000000000000000000000010000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   89  then b_rd <= x"0000000000000000000000000000000000000000020000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   90  then b_rd <= x"0000000000000000000000000000000000000000040000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   91  then b_rd <= x"0000000000000000000000000000000000000000080000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   92  then b_rd <= x"0000000000000000000000000000000000000000100000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   93  then b_rd <= x"0000000000000000000000000000000000000000200000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   94  then b_rd <= x"0000000000000000000000000000000000000000400000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   95  then b_rd <= x"0000000000000000000000000000000000000000800000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   96  then b_rd <= x"0000000000000000000000000000000000000001000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   97  then b_rd <= x"0000000000000000000000000000000000000002000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   98  then b_rd <= x"0000000000000000000000000000000000000004000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =   99  then b_rd <= x"0000000000000000000000000000000000000008000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  100  then b_rd <= x"0000000000000000000000000000000000000010000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  101  then b_rd <= x"0000000000000000000000000000000000000020000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  102  then b_rd <= x"0000000000000000000000000000000000000040000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  103  then b_rd <= x"0000000000000000000000000000000000000080000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  104  then b_rd <= x"0000000000000000000000000000000000000100000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  105  then b_rd <= x"0000000000000000000000000000000000000200000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  106  then b_rd <= x"0000000000000000000000000000000000000400000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  107  then b_rd <= x"0000000000000000000000000000000000000800000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  108  then b_rd <= x"0000000000000000000000000000000000001000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  109  then b_rd <= x"0000000000000000000000000000000000002000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  110  then b_rd <= x"0000000000000000000000000000000000004000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  111  then b_rd <= x"0000000000000000000000000000000000008000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  112  then b_rd <= x"0000000000000000000000000000000000010000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  113  then b_rd <= x"0000000000000000000000000000000000020000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  114  then b_rd <= x"0000000000000000000000000000000000040000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  115  then b_rd <= x"0000000000000000000000000000000000080000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  116  then b_rd <= x"0000000000000000000000000000000000100000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  117  then b_rd <= x"0000000000000000000000000000000000200000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  118  then b_rd <= x"0000000000000000000000000000000000400000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  119  then b_rd <= x"0000000000000000000000000000000000800000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  120  then b_rd <= x"0000000000000000000000000000000001000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  121  then b_rd <= x"0000000000000000000000000000000002000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  122  then b_rd <= x"0000000000000000000000000000000004000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  123  then b_rd <= x"0000000000000000000000000000000008000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  124  then b_rd <= x"0000000000000000000000000000000010000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  125  then b_rd <= x"0000000000000000000000000000000020000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  126  then b_rd <= x"0000000000000000000000000000000040000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  127  then b_rd <= x"0000000000000000000000000000000080000000000000000000000000000000"; end if;

         if conv_integer('0' & buf_num) =  128 then b_rd <= x"0000000000000000000000000000000100000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  129 then b_rd <= x"0000000000000000000000000000000200000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  130 then b_rd <= x"0000000000000000000000000000000400000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  131 then b_rd <= x"0000000000000000000000000000000800000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  132 then b_rd <= x"0000000000000000000000000000001000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  133 then b_rd <= x"0000000000000000000000000000002000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  134 then b_rd <= x"0000000000000000000000000000004000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  135 then b_rd <= x"0000000000000000000000000000008000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  136 then b_rd <= x"0000000000000000000000000000010000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  137 then b_rd <= x"0000000000000000000000000000020000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  138 then b_rd <= x"0000000000000000000000000000040000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  139 then b_rd <= x"0000000000000000000000000000080000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  140 then b_rd <= x"0000000000000000000000000000100000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  141 then b_rd <= x"0000000000000000000000000000200000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  142 then b_rd <= x"0000000000000000000000000000400000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  143 then b_rd <= x"0000000000000000000000000000800000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  144 then b_rd <= x"0000000000000000000000000001000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  145 then b_rd <= x"0000000000000000000000000002000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  146 then b_rd <= x"0000000000000000000000000004000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  147 then b_rd <= x"0000000000000000000000000008000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  148 then b_rd <= x"0000000000000000000000000010000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  149 then b_rd <= x"0000000000000000000000000020000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  150 then b_rd <= x"0000000000000000000000000040000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  151 then b_rd <= x"0000000000000000000000000080000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  152 then b_rd <= x"0000000000000000000000000100000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  153 then b_rd <= x"0000000000000000000000000200000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  154 then b_rd <= x"0000000000000000000000000400000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  155 then b_rd <= x"0000000000000000000000000800000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  156 then b_rd <= x"0000000000000000000000001000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  157 then b_rd <= x"0000000000000000000000002000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  158 then b_rd <= x"0000000000000000000000004000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  159 then b_rd <= x"0000000000000000000000008000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  160 then b_rd <= x"0000000000000000000000010000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  161 then b_rd <= x"0000000000000000000000020000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  162 then b_rd <= x"0000000000000000000000040000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  163 then b_rd <= x"0000000000000000000000080000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  164 then b_rd <= x"0000000000000000000000100000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  165 then b_rd <= x"0000000000000000000000200000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  166 then b_rd <= x"0000000000000000000000400000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  167 then b_rd <= x"0000000000000000000000800000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  168 then b_rd <= x"0000000000000000000001000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  169 then b_rd <= x"0000000000000000000002000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  170 then b_rd <= x"0000000000000000000004000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  171 then b_rd <= x"0000000000000000000008000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  172 then b_rd <= x"0000000000000000000010000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  173 then b_rd <= x"0000000000000000000020000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  174 then b_rd <= x"0000000000000000000040000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  175 then b_rd <= x"0000000000000000000080000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  176 then b_rd <= x"0000000000000000000100000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  177 then b_rd <= x"0000000000000000000200000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  178 then b_rd <= x"0000000000000000000400000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  179 then b_rd <= x"0000000000000000000800000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  180 then b_rd <= x"0000000000000000001000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  181 then b_rd <= x"0000000000000000002000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  182 then b_rd <= x"0000000000000000004000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  183 then b_rd <= x"0000000000000000008000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  184 then b_rd <= x"0000000000000000010000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  185 then b_rd <= x"0000000000000000020000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  186 then b_rd <= x"0000000000000000040000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  187 then b_rd <= x"0000000000000000080000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  188 then b_rd <= x"0000000000000000100000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  189 then b_rd <= x"0000000000000000200000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  190 then b_rd <= x"0000000000000000400000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  191 then b_rd <= x"0000000000000000800000000000000000000000000000000000000000000000"; end if;

         if conv_integer('0' & buf_num) =  192 then b_rd <= x"0000000000000001000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  193 then b_rd <= x"0000000000000002000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  194 then b_rd <= x"0000000000000004000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  195 then b_rd <= x"0000000000000008000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  196 then b_rd <= x"0000000000000010000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  197 then b_rd <= x"0000000000000020000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  198 then b_rd <= x"0000000000000040000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  199 then b_rd <= x"0000000000000080000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  200 then b_rd <= x"0000000000000100000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  201 then b_rd <= x"0000000000000200000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  202 then b_rd <= x"0000000000000400000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  203 then b_rd <= x"0000000000000800000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  204 then b_rd <= x"0000000000001000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  205 then b_rd <= x"0000000000002000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  206 then b_rd <= x"0000000000004000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  207 then b_rd <= x"0000000000008000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  208 then b_rd <= x"0000000000010000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  209 then b_rd <= x"0000000000020000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  210 then b_rd <= x"0000000000040000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  211 then b_rd <= x"0000000000080000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  212 then b_rd <= x"0000000000100000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  213 then b_rd <= x"0000000000200000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  214 then b_rd <= x"0000000000400000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  215 then b_rd <= x"0000000000800000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  216 then b_rd <= x"0000000001000000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  217 then b_rd <= x"0000000002000000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  218 then b_rd <= x"0000000004000000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  219 then b_rd <= x"0000000008000000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  220 then b_rd <= x"0000000010000000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  221 then b_rd <= x"0000000020000000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  222 then b_rd <= x"0000000040000000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  223 then b_rd <= x"0000000080000000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  224 then b_rd <= x"0000000100000000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  225 then b_rd <= x"0000000200000000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  226 then b_rd <= x"0000000400000000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  227 then b_rd <= x"0000000800000000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  228 then b_rd <= x"0000001000000000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  229 then b_rd <= x"0000002000000000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  230 then b_rd <= x"0000004000000000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  231 then b_rd <= x"0000008000000000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  232 then b_rd <= x"0000010000000000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  233 then b_rd <= x"0000020000000000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  234 then b_rd <= x"0000040000000000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  235 then b_rd <= x"0000080000000000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  236 then b_rd <= x"0000100000000000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  237 then b_rd <= x"0000200000000000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  238 then b_rd <= x"0000400000000000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  239 then b_rd <= x"0000800000000000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  240 then b_rd <= x"0001000000000000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  241 then b_rd <= x"0002000000000000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  242 then b_rd <= x"0004000000000000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  243 then b_rd <= x"0008000000000000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  244 then b_rd <= x"0010000000000000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  245 then b_rd <= x"0020000000000000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  246 then b_rd <= x"0040000000000000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  247 then b_rd <= x"0080000000000000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  248 then b_rd <= x"0100000000000000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  249 then b_rd <= x"0200000000000000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  250 then b_rd <= x"0400000000000000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  251 then b_rd <= x"0800000000000000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  252 then b_rd <= x"1000000000000000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  253 then b_rd <= x"2000000000000000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  254 then b_rd <= x"4000000000000000000000000000000000000000000000000000000000000000"; end if;
         if conv_integer('0' & buf_num) =  255 then b_rd <= x"8000000000000000000000000000000000000000000000000000000000000000"; end if;
            --for i in 0 to (2**C_INPUT_SIZE)-1 generate
            ----begin
            --    when (i = conv_integer(buf_num)) => b_rd <= conv_std_logic_vector((i*2), b_rd'length);        
            --end generate;
            --when others => b_rd <= conv_std_logic_vector(0, b_rd'length);
         --end case;
      end if;
      if conv_integer('0' & buf_num) =  0 then d_out <= buff01_out; end if;
      if conv_integer('0' & buf_num) =  1 then d_out <= buff02_out; end if;
      if conv_integer('0' & buf_num) =  2 then d_out <= buff03_out; end if;
      if conv_integer('0' & buf_num) =  3 then d_out <= buff04_out; end if;
      if conv_integer('0' & buf_num) =  4 then d_out <= buff05_out; end if;
      if conv_integer('0' & buf_num) =  5 then d_out <= buff06_out; end if;
      if conv_integer('0' & buf_num) =  6 then d_out <= buff07_out; end if;
      if conv_integer('0' & buf_num) =  7 then d_out <= buff08_out; end if;
      if conv_integer('0' & buf_num) =  8 then d_out <= buff09_out; end if;
      if conv_integer('0' & buf_num) =  9 then d_out <= buff10_out; end if;
      if conv_integer('0' & buf_num) = 10 then d_out <= buff11_out; end if;
      if conv_integer('0' & buf_num) = 11 then d_out <= buff12_out; end if;
      if conv_integer('0' & buf_num) = 12 then d_out <= buff13_out; end if;
      if conv_integer('0' & buf_num) = 13 then d_out <= buff14_out; end if;
      if conv_integer('0' & buf_num) = 14 then d_out <= buff15_out; end if;
      if conv_integer('0' & buf_num) = 15 then d_out <= buff16_out; end if;
      if conv_integer('0' & buf_num) = 16 then d_out <= buff17_out; end if;
      if conv_integer('0' & buf_num) = 17 then d_out <= buff18_out; end if;
      if conv_integer('0' & buf_num) = 18 then d_out <= buff19_out; end if;
      if conv_integer('0' & buf_num) = 19 then d_out <= buff20_out; end if;
      if conv_integer('0' & buf_num) = 20 then d_out <= buff21_out; end if;
      if conv_integer('0' & buf_num) = 21 then d_out <= buff22_out; end if;
      if conv_integer('0' & buf_num) = 22 then d_out <= buff23_out; end if;
      if conv_integer('0' & buf_num) = 23 then d_out <= buff24_out; end if;
      if conv_integer('0' & buf_num) = 24 then d_out <= buff25_out; end if;
      if conv_integer('0' & buf_num) = 25 then d_out <= buff26_out; end if;
      if conv_integer('0' & buf_num) = 26 then d_out <= buff27_out; end if;
      if conv_integer('0' & buf_num) = 27 then d_out <= buff28_out; end if;
      if conv_integer('0' & buf_num) = 28 then d_out <= buff29_out; end if;
      if conv_integer('0' & buf_num) = 29 then d_out <= buff30_out; end if;
      if conv_integer('0' & buf_num) = 30 then d_out <= buff31_out; end if;
      if conv_integer('0' & buf_num) = 31 then d_out <= buff32_out; end if;
      if conv_integer('0' & buf_num) = 32 then d_out <= buff33_out; end if;
      if conv_integer('0' & buf_num) = 33 then d_out <= buff34_out; end if;
      if conv_integer('0' & buf_num) = 34 then d_out <= buff35_out; end if;
      if conv_integer('0' & buf_num) = 35 then d_out <= buff36_out; end if;
      if conv_integer('0' & buf_num) = 36 then d_out <= buff37_out; end if;
      if conv_integer('0' & buf_num) = 37 then d_out <= buff38_out; end if;
      if conv_integer('0' & buf_num) = 38 then d_out <= buff39_out; end if;
      if conv_integer('0' & buf_num) = 39 then d_out <= buff40_out; end if;
      if conv_integer('0' & buf_num) = 40 then d_out <= buff41_out; end if;
      if conv_integer('0' & buf_num) = 41 then d_out <= buff42_out; end if;
      if conv_integer('0' & buf_num) = 42 then d_out <= buff43_out; end if;
      if conv_integer('0' & buf_num) = 43 then d_out <= buff44_out; end if;
      if conv_integer('0' & buf_num) = 44 then d_out <= buff45_out; end if;
      if conv_integer('0' & buf_num) = 45 then d_out <= buff46_out; end if;
      if conv_integer('0' & buf_num) = 46 then d_out <= buff47_out; end if;
      if conv_integer('0' & buf_num) = 47 then d_out <= buff48_out; end if;
      if conv_integer('0' & buf_num) = 48 then d_out <= buff49_out; end if;
      if conv_integer('0' & buf_num) = 49 then d_out <= buff50_out; end if;
      if conv_integer('0' & buf_num) = 50 then d_out <= buff51_out; end if;
      if conv_integer('0' & buf_num) = 51 then d_out <= buff52_out; end if;
      if conv_integer('0' & buf_num) = 52 then d_out <= buff53_out; end if;
      if conv_integer('0' & buf_num) = 53 then d_out <= buff54_out; end if;
      if conv_integer('0' & buf_num) = 54 then d_out <= buff55_out; end if;
      if conv_integer('0' & buf_num) = 55 then d_out <= buff56_out; end if;
      if conv_integer('0' & buf_num) = 56 then d_out <= buff57_out; end if;
      if conv_integer('0' & buf_num) = 57 then d_out <= buff58_out; end if;
      if conv_integer('0' & buf_num) = 58 then d_out <= buff59_out; end if;
      if conv_integer('0' & buf_num) = 59 then d_out <= buff60_out; end if;
      if conv_integer('0' & buf_num) = 60 then d_out <= buff61_out; end if;
      if conv_integer('0' & buf_num) = 61 then d_out <= buff62_out; end if;
      if conv_integer('0' & buf_num) = 62 then d_out <= buff63_out; end if;
      if conv_integer('0' & buf_num) = 63 then d_out <= buff64_out; end if;

      if conv_integer('0' & buf_num) = 64 then d_out <= buff65_out ; end if;
      if conv_integer('0' & buf_num) = 65  then d_out <= buff66_out ; end if;
      if conv_integer('0' & buf_num) = 66  then d_out <= buff67_out ; end if;
      if conv_integer('0' & buf_num) = 67  then d_out <= buff68_out ; end if;
      if conv_integer('0' & buf_num) = 68  then d_out <= buff69_out ; end if;
      if conv_integer('0' & buf_num) = 69  then d_out <= buff70_out ; end if;
      if conv_integer('0' & buf_num) = 70  then d_out <= buff71_out ; end if;
      if conv_integer('0' & buf_num) = 71  then d_out <= buff72_out ; end if;
      if conv_integer('0' & buf_num) = 72  then d_out <= buff73_out ; end if;
      if conv_integer('0' & buf_num) = 73  then d_out <= buff74_out ; end if;
      if conv_integer('0' & buf_num) = 74  then d_out <= buff75_out ; end if;
      if conv_integer('0' & buf_num) = 75  then d_out <= buff76_out ; end if;
      if conv_integer('0' & buf_num) = 76  then d_out <= buff77_out ; end if;
      if conv_integer('0' & buf_num) = 77  then d_out <= buff78_out ; end if;
      if conv_integer('0' & buf_num) = 78  then d_out <= buff79_out ; end if;
      if conv_integer('0' & buf_num) = 79  then d_out <= buff80_out ; end if;
      if conv_integer('0' & buf_num) = 80  then d_out <= buff81_out ; end if;
      if conv_integer('0' & buf_num) = 81  then d_out <= buff82_out ; end if;
      if conv_integer('0' & buf_num) = 82  then d_out <= buff83_out ; end if;
      if conv_integer('0' & buf_num) = 83  then d_out <= buff84_out ; end if;
      if conv_integer('0' & buf_num) = 84  then d_out <= buff85_out ; end if;
      if conv_integer('0' & buf_num) = 85  then d_out <= buff86_out ; end if;
      if conv_integer('0' & buf_num) = 86  then d_out <= buff87_out ; end if;
      if conv_integer('0' & buf_num) = 87  then d_out <= buff88_out ; end if;
      if conv_integer('0' & buf_num) = 88  then d_out <= buff89_out ; end if;
      if conv_integer('0' & buf_num) = 89  then d_out <= buff90_out ; end if;
      if conv_integer('0' & buf_num) = 90  then d_out <= buff91_out ; end if;
      if conv_integer('0' & buf_num) = 91  then d_out <= buff92_out ; end if;
      if conv_integer('0' & buf_num) = 92  then d_out <= buff93_out ; end if;
      if conv_integer('0' & buf_num) = 93  then d_out <= buff94_out ; end if;
      if conv_integer('0' & buf_num) = 94  then d_out <= buff95_out ; end if;
      if conv_integer('0' & buf_num) = 95  then d_out <= buff96_out ; end if;
      if conv_integer('0' & buf_num) = 96  then d_out <= buff97_out ; end if;
      if conv_integer('0' & buf_num) = 97  then d_out <= buff98_out ; end if;
      if conv_integer('0' & buf_num) = 98  then d_out <= buff99_out ; end if;
      if conv_integer('0' & buf_num) = 99  then d_out <= buff100_out; end if;
      if conv_integer('0' & buf_num) =100  then d_out <= buff101_out; end if;
      if conv_integer('0' & buf_num) =101  then d_out <= buff102_out; end if;
      if conv_integer('0' & buf_num) =102  then d_out <= buff103_out; end if;
      if conv_integer('0' & buf_num) =103  then d_out <= buff104_out; end if;
      if conv_integer('0' & buf_num) =104  then d_out <= buff105_out; end if;
      if conv_integer('0' & buf_num) =105  then d_out <= buff106_out; end if;
      if conv_integer('0' & buf_num) =106  then d_out <= buff107_out; end if;
      if conv_integer('0' & buf_num) =107  then d_out <= buff108_out; end if;
      if conv_integer('0' & buf_num) =108  then d_out <= buff109_out; end if;
      if conv_integer('0' & buf_num) =109  then d_out <= buff110_out; end if;
      if conv_integer('0' & buf_num) =110  then d_out <= buff111_out; end if;
      if conv_integer('0' & buf_num) =111  then d_out <= buff112_out; end if;
      if conv_integer('0' & buf_num) =112  then d_out <= buff113_out; end if;
      if conv_integer('0' & buf_num) =113  then d_out <= buff114_out; end if;
      if conv_integer('0' & buf_num) =114  then d_out <= buff115_out; end if;
      if conv_integer('0' & buf_num) =115  then d_out <= buff116_out; end if;
      if conv_integer('0' & buf_num) =116  then d_out <= buff117_out; end if;
      if conv_integer('0' & buf_num) =117  then d_out <= buff118_out; end if;
      if conv_integer('0' & buf_num) =118  then d_out <= buff119_out; end if;
      if conv_integer('0' & buf_num) =119  then d_out <= buff120_out; end if;
      if conv_integer('0' & buf_num) =120  then d_out <= buff121_out; end if;
      if conv_integer('0' & buf_num) =121  then d_out <= buff122_out; end if;
      if conv_integer('0' & buf_num) =122  then d_out <= buff123_out; end if;
      if conv_integer('0' & buf_num) =123  then d_out <= buff124_out; end if;
      if conv_integer('0' & buf_num) =124  then d_out <= buff125_out; end if;
      if conv_integer('0' & buf_num) =125  then d_out <= buff126_out; end if;
      if conv_integer('0' & buf_num) =126  then d_out <= buff127_out; end if;
      if conv_integer('0' & buf_num) =127  then d_out <= buff128_out; end if;

      if conv_integer('0' & buf_num) =128 then d_out <= buff129_out; end if;
      if conv_integer('0' & buf_num) =129 then d_out <= buff130_out; end if;
      if conv_integer('0' & buf_num) =130 then d_out <= buff131_out; end if;
      if conv_integer('0' & buf_num) =131 then d_out <= buff132_out; end if;
      if conv_integer('0' & buf_num) =132 then d_out <= buff133_out; end if;
      if conv_integer('0' & buf_num) =133 then d_out <= buff134_out; end if;
      if conv_integer('0' & buf_num) =134 then d_out <= buff135_out; end if;
      if conv_integer('0' & buf_num) =135 then d_out <= buff136_out; end if;
      if conv_integer('0' & buf_num) =136 then d_out <= buff137_out; end if;
      if conv_integer('0' & buf_num) =137 then d_out <= buff138_out; end if;
      if conv_integer('0' & buf_num) =138 then d_out <= buff139_out; end if;
      if conv_integer('0' & buf_num) =139 then d_out <= buff140_out; end if;
      if conv_integer('0' & buf_num) =140 then d_out <= buff141_out; end if;
      if conv_integer('0' & buf_num) =141 then d_out <= buff142_out; end if;
      if conv_integer('0' & buf_num) =142 then d_out <= buff143_out; end if;
      if conv_integer('0' & buf_num) =143 then d_out <= buff144_out; end if;
      if conv_integer('0' & buf_num) =144 then d_out <= buff145_out; end if;
      if conv_integer('0' & buf_num) =145 then d_out <= buff146_out; end if;
      if conv_integer('0' & buf_num) =146 then d_out <= buff147_out; end if;
      if conv_integer('0' & buf_num) =147 then d_out <= buff148_out; end if;
      if conv_integer('0' & buf_num) =148 then d_out <= buff149_out; end if;
      if conv_integer('0' & buf_num) =149 then d_out <= buff150_out; end if;
      if conv_integer('0' & buf_num) =150 then d_out <= buff151_out; end if;
      if conv_integer('0' & buf_num) =151 then d_out <= buff152_out; end if;
      if conv_integer('0' & buf_num) =152 then d_out <= buff153_out; end if;
      if conv_integer('0' & buf_num) =153 then d_out <= buff154_out; end if;
      if conv_integer('0' & buf_num) =154 then d_out <= buff155_out; end if;
      if conv_integer('0' & buf_num) =155 then d_out <= buff156_out; end if;
      if conv_integer('0' & buf_num) =156 then d_out <= buff157_out; end if;
      if conv_integer('0' & buf_num) =157 then d_out <= buff158_out; end if;
      if conv_integer('0' & buf_num) =158 then d_out <= buff159_out; end if;
      if conv_integer('0' & buf_num) =159 then d_out <= buff160_out; end if;
      if conv_integer('0' & buf_num) =160 then d_out <= buff161_out; end if;
      if conv_integer('0' & buf_num) =161 then d_out <= buff162_out; end if;
      if conv_integer('0' & buf_num) =162 then d_out <= buff163_out; end if;
      if conv_integer('0' & buf_num) =163 then d_out <= buff164_out; end if;
      if conv_integer('0' & buf_num) =164 then d_out <= buff165_out; end if;
      if conv_integer('0' & buf_num) =165 then d_out <= buff166_out; end if;
      if conv_integer('0' & buf_num) =166 then d_out <= buff167_out; end if;
      if conv_integer('0' & buf_num) =167 then d_out <= buff168_out; end if;
      if conv_integer('0' & buf_num) =168 then d_out <= buff169_out; end if;
      if conv_integer('0' & buf_num) =169 then d_out <= buff170_out; end if;
      if conv_integer('0' & buf_num) =170 then d_out <= buff171_out; end if;
      if conv_integer('0' & buf_num) =171 then d_out <= buff172_out; end if;
      if conv_integer('0' & buf_num) =172 then d_out <= buff173_out; end if;
      if conv_integer('0' & buf_num) =173 then d_out <= buff174_out; end if;
      if conv_integer('0' & buf_num) =174 then d_out <= buff175_out; end if;
      if conv_integer('0' & buf_num) =175 then d_out <= buff176_out; end if;
      if conv_integer('0' & buf_num) =176 then d_out <= buff177_out; end if;
      if conv_integer('0' & buf_num) =177 then d_out <= buff178_out; end if;
      if conv_integer('0' & buf_num) =178 then d_out <= buff179_out; end if;
      if conv_integer('0' & buf_num) =179 then d_out <= buff180_out; end if;
      if conv_integer('0' & buf_num) =180 then d_out <= buff181_out; end if;
      if conv_integer('0' & buf_num) =181 then d_out <= buff182_out; end if;
      if conv_integer('0' & buf_num) =182 then d_out <= buff183_out; end if;
      if conv_integer('0' & buf_num) =183 then d_out <= buff184_out; end if;
      if conv_integer('0' & buf_num) =184 then d_out <= buff185_out; end if;
      if conv_integer('0' & buf_num) =185 then d_out <= buff186_out; end if;
      if conv_integer('0' & buf_num) =186 then d_out <= buff187_out; end if;
      if conv_integer('0' & buf_num) =187 then d_out <= buff188_out; end if;
      if conv_integer('0' & buf_num) =188 then d_out <= buff189_out; end if;
      if conv_integer('0' & buf_num) =189 then d_out <= buff190_out; end if;
      if conv_integer('0' & buf_num) =190 then d_out <= buff191_out; end if;
      if conv_integer('0' & buf_num) =191 then d_out <= buff192_out; end if;

      if conv_integer('0' & buf_num) =192 then d_out <= buff01_out; end if;
      if conv_integer('0' & buf_num) =193 then d_out <= buff02_out; end if;
      if conv_integer('0' & buf_num) =194 then d_out <= buff03_out; end if;
      if conv_integer('0' & buf_num) =195 then d_out <= buff04_out; end if;
      if conv_integer('0' & buf_num) =196 then d_out <= buff05_out; end if;
      if conv_integer('0' & buf_num) =197 then d_out <= buff06_out; end if;
      if conv_integer('0' & buf_num) =198 then d_out <= buff07_out; end if;
      if conv_integer('0' & buf_num) =199 then d_out <= buff08_out; end if;
      if conv_integer('0' & buf_num) =200 then d_out <= buff09_out; end if;
      if conv_integer('0' & buf_num) =201 then d_out <= buff10_out; end if;
      if conv_integer('0' & buf_num) =202 then d_out <= buff11_out; end if;
      if conv_integer('0' & buf_num) =203 then d_out <= buff12_out; end if;
      if conv_integer('0' & buf_num) =204 then d_out <= buff13_out; end if;
      if conv_integer('0' & buf_num) =205 then d_out <= buff14_out; end if;
      if conv_integer('0' & buf_num) =206 then d_out <= buff15_out; end if;
      if conv_integer('0' & buf_num) =207 then d_out <= buff16_out; end if;
      if conv_integer('0' & buf_num) =208 then d_out <= buff17_out; end if;
      if conv_integer('0' & buf_num) =209 then d_out <= buff18_out; end if;
      if conv_integer('0' & buf_num) =210 then d_out <= buff19_out; end if;
      if conv_integer('0' & buf_num) =211 then d_out <= buff20_out; end if;
      if conv_integer('0' & buf_num) =212 then d_out <= buff21_out; end if;
      if conv_integer('0' & buf_num) =213 then d_out <= buff22_out; end if;
      if conv_integer('0' & buf_num) =214 then d_out <= buff23_out; end if;
      if conv_integer('0' & buf_num) =215 then d_out <= buff24_out; end if;
      if conv_integer('0' & buf_num) =216 then d_out <= buff25_out; end if;
      if conv_integer('0' & buf_num) =217 then d_out <= buff26_out; end if;
      if conv_integer('0' & buf_num) =218 then d_out <= buff27_out; end if;
      if conv_integer('0' & buf_num) =219 then d_out <= buff28_out; end if;
      if conv_integer('0' & buf_num) =220 then d_out <= buff29_out; end if;
      if conv_integer('0' & buf_num) =221 then d_out <= buff30_out; end if;
      if conv_integer('0' & buf_num) =222 then d_out <= buff31_out; end if;
      if conv_integer('0' & buf_num) =223 then d_out <= buff32_out; end if;
      if conv_integer('0' & buf_num) =224 then d_out <= buff33_out; end if;
      if conv_integer('0' & buf_num) =225 then d_out <= buff34_out; end if;
      if conv_integer('0' & buf_num) =226 then d_out <= buff35_out; end if;
      if conv_integer('0' & buf_num) =227 then d_out <= buff36_out; end if;
      if conv_integer('0' & buf_num) =228 then d_out <= buff37_out; end if;
      if conv_integer('0' & buf_num) =229 then d_out <= buff38_out; end if;
      if conv_integer('0' & buf_num) =230 then d_out <= buff39_out; end if;
      if conv_integer('0' & buf_num) =231 then d_out <= buff40_out; end if;
      if conv_integer('0' & buf_num) =232 then d_out <= buff41_out; end if;
      if conv_integer('0' & buf_num) =233 then d_out <= buff42_out; end if;
      if conv_integer('0' & buf_num) =234 then d_out <= buff43_out; end if;
      if conv_integer('0' & buf_num) =235 then d_out <= buff44_out; end if;
      if conv_integer('0' & buf_num) =236 then d_out <= buff45_out; end if;
      if conv_integer('0' & buf_num) =237 then d_out <= buff46_out; end if;
      if conv_integer('0' & buf_num) =238 then d_out <= buff47_out; end if;
      if conv_integer('0' & buf_num) =239 then d_out <= buff48_out; end if;
      if conv_integer('0' & buf_num) =240 then d_out <= buff49_out; end if;
      if conv_integer('0' & buf_num) =241 then d_out <= buff50_out; end if;
      if conv_integer('0' & buf_num) =242 then d_out <= buff51_out; end if;
      if conv_integer('0' & buf_num) =243 then d_out <= buff52_out; end if;
      if conv_integer('0' & buf_num) =244 then d_out <= buff53_out; end if;
      if conv_integer('0' & buf_num) =245 then d_out <= buff54_out; end if;
      if conv_integer('0' & buf_num) =246 then d_out <= buff55_out; end if;
      if conv_integer('0' & buf_num) =247 then d_out <= buff56_out; end if;
      if conv_integer('0' & buf_num) =248 then d_out <= buff57_out; end if;
      if conv_integer('0' & buf_num) =249 then d_out <= buff58_out; end if;
      if conv_integer('0' & buf_num) =250 then d_out <= buff59_out; end if;
      if conv_integer('0' & buf_num) =251 then d_out <= buff60_out; end if;
      if conv_integer('0' & buf_num) =252 then d_out <= buff61_out; end if;
      if conv_integer('0' & buf_num) =253 then d_out <= buff62_out; end if;
      if conv_integer('0' & buf_num) =254 then d_out <= buff63_out; end if;
      if conv_integer('0' & buf_num) =255 then d_out <= buff64_out; end if;
   end if;
end process p_rd_ctr;

end a;