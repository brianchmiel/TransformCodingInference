library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_SIGNED.ALL;

entity multROM is
  port    (
           clk           : in  std_logic;

           ROM_addr      : in  std_logic_vector(15 downto 0);
           ROM_data      : out std_logic_vector( 7 downto 0)
           );                        
end multROM;

architecture a of multROM is

    type ROM_Array is array (0 to (2**16-1)) 
  of std_logic_vector(7 downto 0);

    constant Content: ROM_Array := (
0 => conv_std_logic_vector(0, 8),
1 => conv_std_logic_vector(0, 8),
2 => conv_std_logic_vector(0, 8),
3 => conv_std_logic_vector(0, 8),
4 => conv_std_logic_vector(0, 8),
5 => conv_std_logic_vector(0, 8),
6 => conv_std_logic_vector(0, 8),
7 => conv_std_logic_vector(0, 8),
8 => conv_std_logic_vector(0, 8),
9 => conv_std_logic_vector(0, 8),
10 => conv_std_logic_vector(0, 8),
11 => conv_std_logic_vector(0, 8),
12 => conv_std_logic_vector(0, 8),
13 => conv_std_logic_vector(0, 8),
14 => conv_std_logic_vector(0, 8),
15 => conv_std_logic_vector(0, 8),
16 => conv_std_logic_vector(0, 8),
17 => conv_std_logic_vector(0, 8),
18 => conv_std_logic_vector(0, 8),
19 => conv_std_logic_vector(0, 8),
20 => conv_std_logic_vector(0, 8),
21 => conv_std_logic_vector(0, 8),
22 => conv_std_logic_vector(0, 8),
23 => conv_std_logic_vector(0, 8),
24 => conv_std_logic_vector(0, 8),
25 => conv_std_logic_vector(0, 8),
26 => conv_std_logic_vector(0, 8),
27 => conv_std_logic_vector(0, 8),
28 => conv_std_logic_vector(0, 8),
29 => conv_std_logic_vector(0, 8),
30 => conv_std_logic_vector(0, 8),
31 => conv_std_logic_vector(0, 8),
32 => conv_std_logic_vector(0, 8),
33 => conv_std_logic_vector(0, 8),
34 => conv_std_logic_vector(0, 8),
35 => conv_std_logic_vector(0, 8),
36 => conv_std_logic_vector(0, 8),
37 => conv_std_logic_vector(0, 8),
38 => conv_std_logic_vector(0, 8),
39 => conv_std_logic_vector(0, 8),
40 => conv_std_logic_vector(0, 8),
41 => conv_std_logic_vector(0, 8),
42 => conv_std_logic_vector(0, 8),
43 => conv_std_logic_vector(0, 8),
44 => conv_std_logic_vector(0, 8),
45 => conv_std_logic_vector(0, 8),
46 => conv_std_logic_vector(0, 8),
47 => conv_std_logic_vector(0, 8),
48 => conv_std_logic_vector(0, 8),
49 => conv_std_logic_vector(0, 8),
50 => conv_std_logic_vector(0, 8),
51 => conv_std_logic_vector(0, 8),
52 => conv_std_logic_vector(0, 8),
53 => conv_std_logic_vector(0, 8),
54 => conv_std_logic_vector(0, 8),
55 => conv_std_logic_vector(0, 8),
56 => conv_std_logic_vector(0, 8),
57 => conv_std_logic_vector(0, 8),
58 => conv_std_logic_vector(0, 8),
59 => conv_std_logic_vector(0, 8),
60 => conv_std_logic_vector(0, 8),
61 => conv_std_logic_vector(0, 8),
62 => conv_std_logic_vector(0, 8),
63 => conv_std_logic_vector(0, 8),
64 => conv_std_logic_vector(0, 8),
65 => conv_std_logic_vector(0, 8),
66 => conv_std_logic_vector(0, 8),
67 => conv_std_logic_vector(0, 8),
68 => conv_std_logic_vector(0, 8),
69 => conv_std_logic_vector(0, 8),
70 => conv_std_logic_vector(0, 8),
71 => conv_std_logic_vector(0, 8),
72 => conv_std_logic_vector(0, 8),
73 => conv_std_logic_vector(0, 8),
74 => conv_std_logic_vector(0, 8),
75 => conv_std_logic_vector(0, 8),
76 => conv_std_logic_vector(0, 8),
77 => conv_std_logic_vector(0, 8),
78 => conv_std_logic_vector(0, 8),
79 => conv_std_logic_vector(0, 8),
80 => conv_std_logic_vector(0, 8),
81 => conv_std_logic_vector(0, 8),
82 => conv_std_logic_vector(0, 8),
83 => conv_std_logic_vector(0, 8),
84 => conv_std_logic_vector(0, 8),
85 => conv_std_logic_vector(0, 8),
86 => conv_std_logic_vector(0, 8),
87 => conv_std_logic_vector(0, 8),
88 => conv_std_logic_vector(0, 8),
89 => conv_std_logic_vector(0, 8),
90 => conv_std_logic_vector(0, 8),
91 => conv_std_logic_vector(0, 8),
92 => conv_std_logic_vector(0, 8),
93 => conv_std_logic_vector(0, 8),
94 => conv_std_logic_vector(0, 8),
95 => conv_std_logic_vector(0, 8),
96 => conv_std_logic_vector(0, 8),
97 => conv_std_logic_vector(0, 8),
98 => conv_std_logic_vector(0, 8),
99 => conv_std_logic_vector(0, 8),
100 => conv_std_logic_vector(0, 8),
101 => conv_std_logic_vector(0, 8),
102 => conv_std_logic_vector(0, 8),
103 => conv_std_logic_vector(0, 8),
104 => conv_std_logic_vector(0, 8),
105 => conv_std_logic_vector(0, 8),
106 => conv_std_logic_vector(0, 8),
107 => conv_std_logic_vector(0, 8),
108 => conv_std_logic_vector(0, 8),
109 => conv_std_logic_vector(0, 8),
110 => conv_std_logic_vector(0, 8),
111 => conv_std_logic_vector(0, 8),
112 => conv_std_logic_vector(0, 8),
113 => conv_std_logic_vector(0, 8),
114 => conv_std_logic_vector(0, 8),
115 => conv_std_logic_vector(0, 8),
116 => conv_std_logic_vector(0, 8),
117 => conv_std_logic_vector(0, 8),
118 => conv_std_logic_vector(0, 8),
119 => conv_std_logic_vector(0, 8),
120 => conv_std_logic_vector(0, 8),
121 => conv_std_logic_vector(0, 8),
122 => conv_std_logic_vector(0, 8),
123 => conv_std_logic_vector(0, 8),
124 => conv_std_logic_vector(0, 8),
125 => conv_std_logic_vector(0, 8),
126 => conv_std_logic_vector(0, 8),
127 => conv_std_logic_vector(0, 8),
128 => conv_std_logic_vector(0, 8),
129 => conv_std_logic_vector(0, 8),
130 => conv_std_logic_vector(0, 8),
131 => conv_std_logic_vector(0, 8),
132 => conv_std_logic_vector(0, 8),
133 => conv_std_logic_vector(0, 8),
134 => conv_std_logic_vector(0, 8),
135 => conv_std_logic_vector(0, 8),
136 => conv_std_logic_vector(0, 8),
137 => conv_std_logic_vector(0, 8),
138 => conv_std_logic_vector(0, 8),
139 => conv_std_logic_vector(0, 8),
140 => conv_std_logic_vector(0, 8),
141 => conv_std_logic_vector(0, 8),
142 => conv_std_logic_vector(0, 8),
143 => conv_std_logic_vector(0, 8),
144 => conv_std_logic_vector(0, 8),
145 => conv_std_logic_vector(0, 8),
146 => conv_std_logic_vector(0, 8),
147 => conv_std_logic_vector(0, 8),
148 => conv_std_logic_vector(0, 8),
149 => conv_std_logic_vector(0, 8),
150 => conv_std_logic_vector(0, 8),
151 => conv_std_logic_vector(0, 8),
152 => conv_std_logic_vector(0, 8),
153 => conv_std_logic_vector(0, 8),
154 => conv_std_logic_vector(0, 8),
155 => conv_std_logic_vector(0, 8),
156 => conv_std_logic_vector(0, 8),
157 => conv_std_logic_vector(0, 8),
158 => conv_std_logic_vector(0, 8),
159 => conv_std_logic_vector(0, 8),
160 => conv_std_logic_vector(0, 8),
161 => conv_std_logic_vector(0, 8),
162 => conv_std_logic_vector(0, 8),
163 => conv_std_logic_vector(0, 8),
164 => conv_std_logic_vector(0, 8),
165 => conv_std_logic_vector(0, 8),
166 => conv_std_logic_vector(0, 8),
167 => conv_std_logic_vector(0, 8),
168 => conv_std_logic_vector(0, 8),
169 => conv_std_logic_vector(0, 8),
170 => conv_std_logic_vector(0, 8),
171 => conv_std_logic_vector(0, 8),
172 => conv_std_logic_vector(0, 8),
173 => conv_std_logic_vector(0, 8),
174 => conv_std_logic_vector(0, 8),
175 => conv_std_logic_vector(0, 8),
176 => conv_std_logic_vector(0, 8),
177 => conv_std_logic_vector(0, 8),
178 => conv_std_logic_vector(0, 8),
179 => conv_std_logic_vector(0, 8),
180 => conv_std_logic_vector(0, 8),
181 => conv_std_logic_vector(0, 8),
182 => conv_std_logic_vector(0, 8),
183 => conv_std_logic_vector(0, 8),
184 => conv_std_logic_vector(0, 8),
185 => conv_std_logic_vector(0, 8),
186 => conv_std_logic_vector(0, 8),
187 => conv_std_logic_vector(0, 8),
188 => conv_std_logic_vector(0, 8),
189 => conv_std_logic_vector(0, 8),
190 => conv_std_logic_vector(0, 8),
191 => conv_std_logic_vector(0, 8),
192 => conv_std_logic_vector(0, 8),
193 => conv_std_logic_vector(0, 8),
194 => conv_std_logic_vector(0, 8),
195 => conv_std_logic_vector(0, 8),
196 => conv_std_logic_vector(0, 8),
197 => conv_std_logic_vector(0, 8),
198 => conv_std_logic_vector(0, 8),
199 => conv_std_logic_vector(0, 8),
200 => conv_std_logic_vector(0, 8),
201 => conv_std_logic_vector(0, 8),
202 => conv_std_logic_vector(0, 8),
203 => conv_std_logic_vector(0, 8),
204 => conv_std_logic_vector(0, 8),
205 => conv_std_logic_vector(0, 8),
206 => conv_std_logic_vector(0, 8),
207 => conv_std_logic_vector(0, 8),
208 => conv_std_logic_vector(0, 8),
209 => conv_std_logic_vector(0, 8),
210 => conv_std_logic_vector(0, 8),
211 => conv_std_logic_vector(0, 8),
212 => conv_std_logic_vector(0, 8),
213 => conv_std_logic_vector(0, 8),
214 => conv_std_logic_vector(0, 8),
215 => conv_std_logic_vector(0, 8),
216 => conv_std_logic_vector(0, 8),
217 => conv_std_logic_vector(0, 8),
218 => conv_std_logic_vector(0, 8),
219 => conv_std_logic_vector(0, 8),
220 => conv_std_logic_vector(0, 8),
221 => conv_std_logic_vector(0, 8),
222 => conv_std_logic_vector(0, 8),
223 => conv_std_logic_vector(0, 8),
224 => conv_std_logic_vector(0, 8),
225 => conv_std_logic_vector(0, 8),
226 => conv_std_logic_vector(0, 8),
227 => conv_std_logic_vector(0, 8),
228 => conv_std_logic_vector(0, 8),
229 => conv_std_logic_vector(0, 8),
230 => conv_std_logic_vector(0, 8),
231 => conv_std_logic_vector(0, 8),
232 => conv_std_logic_vector(0, 8),
233 => conv_std_logic_vector(0, 8),
234 => conv_std_logic_vector(0, 8),
235 => conv_std_logic_vector(0, 8),
236 => conv_std_logic_vector(0, 8),
237 => conv_std_logic_vector(0, 8),
238 => conv_std_logic_vector(0, 8),
239 => conv_std_logic_vector(0, 8),
240 => conv_std_logic_vector(0, 8),
241 => conv_std_logic_vector(0, 8),
242 => conv_std_logic_vector(0, 8),
243 => conv_std_logic_vector(0, 8),
244 => conv_std_logic_vector(0, 8),
245 => conv_std_logic_vector(0, 8),
246 => conv_std_logic_vector(0, 8),
247 => conv_std_logic_vector(0, 8),
248 => conv_std_logic_vector(0, 8),
249 => conv_std_logic_vector(0, 8),
250 => conv_std_logic_vector(0, 8),
251 => conv_std_logic_vector(0, 8),
252 => conv_std_logic_vector(0, 8),
253 => conv_std_logic_vector(0, 8),
254 => conv_std_logic_vector(0, 8),
255 => conv_std_logic_vector(0, 8),
256 => conv_std_logic_vector(0, 8),
257 => conv_std_logic_vector(0, 8),
258 => conv_std_logic_vector(0, 8),
259 => conv_std_logic_vector(0, 8),
260 => conv_std_logic_vector(0, 8),
261 => conv_std_logic_vector(0, 8),
262 => conv_std_logic_vector(0, 8),
263 => conv_std_logic_vector(0, 8),
264 => conv_std_logic_vector(0, 8),
265 => conv_std_logic_vector(0, 8),
266 => conv_std_logic_vector(0, 8),
267 => conv_std_logic_vector(0, 8),
268 => conv_std_logic_vector(0, 8),
269 => conv_std_logic_vector(0, 8),
270 => conv_std_logic_vector(0, 8),
271 => conv_std_logic_vector(0, 8),
272 => conv_std_logic_vector(0, 8),
273 => conv_std_logic_vector(0, 8),
274 => conv_std_logic_vector(0, 8),
275 => conv_std_logic_vector(0, 8),
276 => conv_std_logic_vector(0, 8),
277 => conv_std_logic_vector(0, 8),
278 => conv_std_logic_vector(0, 8),
279 => conv_std_logic_vector(0, 8),
280 => conv_std_logic_vector(0, 8),
281 => conv_std_logic_vector(0, 8),
282 => conv_std_logic_vector(0, 8),
283 => conv_std_logic_vector(0, 8),
284 => conv_std_logic_vector(0, 8),
285 => conv_std_logic_vector(0, 8),
286 => conv_std_logic_vector(0, 8),
287 => conv_std_logic_vector(0, 8),
288 => conv_std_logic_vector(0, 8),
289 => conv_std_logic_vector(0, 8),
290 => conv_std_logic_vector(0, 8),
291 => conv_std_logic_vector(0, 8),
292 => conv_std_logic_vector(0, 8),
293 => conv_std_logic_vector(0, 8),
294 => conv_std_logic_vector(0, 8),
295 => conv_std_logic_vector(0, 8),
296 => conv_std_logic_vector(0, 8),
297 => conv_std_logic_vector(0, 8),
298 => conv_std_logic_vector(0, 8),
299 => conv_std_logic_vector(0, 8),
300 => conv_std_logic_vector(0, 8),
301 => conv_std_logic_vector(0, 8),
302 => conv_std_logic_vector(0, 8),
303 => conv_std_logic_vector(0, 8),
304 => conv_std_logic_vector(0, 8),
305 => conv_std_logic_vector(0, 8),
306 => conv_std_logic_vector(0, 8),
307 => conv_std_logic_vector(0, 8),
308 => conv_std_logic_vector(0, 8),
309 => conv_std_logic_vector(0, 8),
310 => conv_std_logic_vector(0, 8),
311 => conv_std_logic_vector(0, 8),
312 => conv_std_logic_vector(0, 8),
313 => conv_std_logic_vector(0, 8),
314 => conv_std_logic_vector(0, 8),
315 => conv_std_logic_vector(0, 8),
316 => conv_std_logic_vector(0, 8),
317 => conv_std_logic_vector(0, 8),
318 => conv_std_logic_vector(0, 8),
319 => conv_std_logic_vector(0, 8),
320 => conv_std_logic_vector(0, 8),
321 => conv_std_logic_vector(0, 8),
322 => conv_std_logic_vector(0, 8),
323 => conv_std_logic_vector(0, 8),
324 => conv_std_logic_vector(0, 8),
325 => conv_std_logic_vector(0, 8),
326 => conv_std_logic_vector(0, 8),
327 => conv_std_logic_vector(0, 8),
328 => conv_std_logic_vector(0, 8),
329 => conv_std_logic_vector(0, 8),
330 => conv_std_logic_vector(0, 8),
331 => conv_std_logic_vector(0, 8),
332 => conv_std_logic_vector(0, 8),
333 => conv_std_logic_vector(0, 8),
334 => conv_std_logic_vector(0, 8),
335 => conv_std_logic_vector(0, 8),
336 => conv_std_logic_vector(0, 8),
337 => conv_std_logic_vector(0, 8),
338 => conv_std_logic_vector(0, 8),
339 => conv_std_logic_vector(0, 8),
340 => conv_std_logic_vector(0, 8),
341 => conv_std_logic_vector(0, 8),
342 => conv_std_logic_vector(0, 8),
343 => conv_std_logic_vector(0, 8),
344 => conv_std_logic_vector(0, 8),
345 => conv_std_logic_vector(0, 8),
346 => conv_std_logic_vector(0, 8),
347 => conv_std_logic_vector(0, 8),
348 => conv_std_logic_vector(0, 8),
349 => conv_std_logic_vector(0, 8),
350 => conv_std_logic_vector(0, 8),
351 => conv_std_logic_vector(0, 8),
352 => conv_std_logic_vector(0, 8),
353 => conv_std_logic_vector(0, 8),
354 => conv_std_logic_vector(0, 8),
355 => conv_std_logic_vector(0, 8),
356 => conv_std_logic_vector(0, 8),
357 => conv_std_logic_vector(0, 8),
358 => conv_std_logic_vector(0, 8),
359 => conv_std_logic_vector(0, 8),
360 => conv_std_logic_vector(0, 8),
361 => conv_std_logic_vector(0, 8),
362 => conv_std_logic_vector(0, 8),
363 => conv_std_logic_vector(0, 8),
364 => conv_std_logic_vector(0, 8),
365 => conv_std_logic_vector(0, 8),
366 => conv_std_logic_vector(0, 8),
367 => conv_std_logic_vector(0, 8),
368 => conv_std_logic_vector(0, 8),
369 => conv_std_logic_vector(0, 8),
370 => conv_std_logic_vector(0, 8),
371 => conv_std_logic_vector(0, 8),
372 => conv_std_logic_vector(0, 8),
373 => conv_std_logic_vector(0, 8),
374 => conv_std_logic_vector(0, 8),
375 => conv_std_logic_vector(0, 8),
376 => conv_std_logic_vector(0, 8),
377 => conv_std_logic_vector(0, 8),
378 => conv_std_logic_vector(0, 8),
379 => conv_std_logic_vector(0, 8),
380 => conv_std_logic_vector(0, 8),
381 => conv_std_logic_vector(0, 8),
382 => conv_std_logic_vector(0, 8),
383 => conv_std_logic_vector(0, 8),
384 => conv_std_logic_vector(0, 8),
385 => conv_std_logic_vector(0, 8),
386 => conv_std_logic_vector(0, 8),
387 => conv_std_logic_vector(0, 8),
388 => conv_std_logic_vector(0, 8),
389 => conv_std_logic_vector(0, 8),
390 => conv_std_logic_vector(0, 8),
391 => conv_std_logic_vector(0, 8),
392 => conv_std_logic_vector(0, 8),
393 => conv_std_logic_vector(0, 8),
394 => conv_std_logic_vector(0, 8),
395 => conv_std_logic_vector(0, 8),
396 => conv_std_logic_vector(0, 8),
397 => conv_std_logic_vector(0, 8),
398 => conv_std_logic_vector(0, 8),
399 => conv_std_logic_vector(0, 8),
400 => conv_std_logic_vector(0, 8),
401 => conv_std_logic_vector(0, 8),
402 => conv_std_logic_vector(0, 8),
403 => conv_std_logic_vector(0, 8),
404 => conv_std_logic_vector(0, 8),
405 => conv_std_logic_vector(0, 8),
406 => conv_std_logic_vector(0, 8),
407 => conv_std_logic_vector(0, 8),
408 => conv_std_logic_vector(0, 8),
409 => conv_std_logic_vector(0, 8),
410 => conv_std_logic_vector(0, 8),
411 => conv_std_logic_vector(0, 8),
412 => conv_std_logic_vector(0, 8),
413 => conv_std_logic_vector(0, 8),
414 => conv_std_logic_vector(0, 8),
415 => conv_std_logic_vector(0, 8),
416 => conv_std_logic_vector(0, 8),
417 => conv_std_logic_vector(0, 8),
418 => conv_std_logic_vector(0, 8),
419 => conv_std_logic_vector(0, 8),
420 => conv_std_logic_vector(0, 8),
421 => conv_std_logic_vector(0, 8),
422 => conv_std_logic_vector(0, 8),
423 => conv_std_logic_vector(0, 8),
424 => conv_std_logic_vector(0, 8),
425 => conv_std_logic_vector(0, 8),
426 => conv_std_logic_vector(0, 8),
427 => conv_std_logic_vector(0, 8),
428 => conv_std_logic_vector(0, 8),
429 => conv_std_logic_vector(0, 8),
430 => conv_std_logic_vector(0, 8),
431 => conv_std_logic_vector(0, 8),
432 => conv_std_logic_vector(0, 8),
433 => conv_std_logic_vector(0, 8),
434 => conv_std_logic_vector(0, 8),
435 => conv_std_logic_vector(0, 8),
436 => conv_std_logic_vector(0, 8),
437 => conv_std_logic_vector(0, 8),
438 => conv_std_logic_vector(0, 8),
439 => conv_std_logic_vector(0, 8),
440 => conv_std_logic_vector(0, 8),
441 => conv_std_logic_vector(0, 8),
442 => conv_std_logic_vector(0, 8),
443 => conv_std_logic_vector(0, 8),
444 => conv_std_logic_vector(0, 8),
445 => conv_std_logic_vector(0, 8),
446 => conv_std_logic_vector(0, 8),
447 => conv_std_logic_vector(0, 8),
448 => conv_std_logic_vector(0, 8),
449 => conv_std_logic_vector(0, 8),
450 => conv_std_logic_vector(0, 8),
451 => conv_std_logic_vector(0, 8),
452 => conv_std_logic_vector(0, 8),
453 => conv_std_logic_vector(0, 8),
454 => conv_std_logic_vector(0, 8),
455 => conv_std_logic_vector(0, 8),
456 => conv_std_logic_vector(0, 8),
457 => conv_std_logic_vector(0, 8),
458 => conv_std_logic_vector(0, 8),
459 => conv_std_logic_vector(0, 8),
460 => conv_std_logic_vector(0, 8),
461 => conv_std_logic_vector(0, 8),
462 => conv_std_logic_vector(0, 8),
463 => conv_std_logic_vector(0, 8),
464 => conv_std_logic_vector(0, 8),
465 => conv_std_logic_vector(0, 8),
466 => conv_std_logic_vector(0, 8),
467 => conv_std_logic_vector(0, 8),
468 => conv_std_logic_vector(0, 8),
469 => conv_std_logic_vector(0, 8),
470 => conv_std_logic_vector(0, 8),
471 => conv_std_logic_vector(0, 8),
472 => conv_std_logic_vector(0, 8),
473 => conv_std_logic_vector(0, 8),
474 => conv_std_logic_vector(0, 8),
475 => conv_std_logic_vector(0, 8),
476 => conv_std_logic_vector(0, 8),
477 => conv_std_logic_vector(0, 8),
478 => conv_std_logic_vector(0, 8),
479 => conv_std_logic_vector(0, 8),
480 => conv_std_logic_vector(0, 8),
481 => conv_std_logic_vector(0, 8),
482 => conv_std_logic_vector(0, 8),
483 => conv_std_logic_vector(0, 8),
484 => conv_std_logic_vector(0, 8),
485 => conv_std_logic_vector(0, 8),
486 => conv_std_logic_vector(0, 8),
487 => conv_std_logic_vector(0, 8),
488 => conv_std_logic_vector(0, 8),
489 => conv_std_logic_vector(0, 8),
490 => conv_std_logic_vector(0, 8),
491 => conv_std_logic_vector(0, 8),
492 => conv_std_logic_vector(0, 8),
493 => conv_std_logic_vector(0, 8),
494 => conv_std_logic_vector(0, 8),
495 => conv_std_logic_vector(0, 8),
496 => conv_std_logic_vector(0, 8),
497 => conv_std_logic_vector(0, 8),
498 => conv_std_logic_vector(0, 8),
499 => conv_std_logic_vector(0, 8),
500 => conv_std_logic_vector(0, 8),
501 => conv_std_logic_vector(0, 8),
502 => conv_std_logic_vector(0, 8),
503 => conv_std_logic_vector(0, 8),
504 => conv_std_logic_vector(0, 8),
505 => conv_std_logic_vector(0, 8),
506 => conv_std_logic_vector(0, 8),
507 => conv_std_logic_vector(0, 8),
508 => conv_std_logic_vector(0, 8),
509 => conv_std_logic_vector(0, 8),
510 => conv_std_logic_vector(0, 8),
511 => conv_std_logic_vector(0, 8),
512 => conv_std_logic_vector(0, 8),
513 => conv_std_logic_vector(0, 8),
514 => conv_std_logic_vector(0, 8),
515 => conv_std_logic_vector(0, 8),
516 => conv_std_logic_vector(0, 8),
517 => conv_std_logic_vector(0, 8),
518 => conv_std_logic_vector(0, 8),
519 => conv_std_logic_vector(0, 8),
520 => conv_std_logic_vector(0, 8),
521 => conv_std_logic_vector(0, 8),
522 => conv_std_logic_vector(0, 8),
523 => conv_std_logic_vector(0, 8),
524 => conv_std_logic_vector(0, 8),
525 => conv_std_logic_vector(0, 8),
526 => conv_std_logic_vector(0, 8),
527 => conv_std_logic_vector(0, 8),
528 => conv_std_logic_vector(0, 8),
529 => conv_std_logic_vector(0, 8),
530 => conv_std_logic_vector(0, 8),
531 => conv_std_logic_vector(0, 8),
532 => conv_std_logic_vector(0, 8),
533 => conv_std_logic_vector(0, 8),
534 => conv_std_logic_vector(0, 8),
535 => conv_std_logic_vector(0, 8),
536 => conv_std_logic_vector(0, 8),
537 => conv_std_logic_vector(0, 8),
538 => conv_std_logic_vector(0, 8),
539 => conv_std_logic_vector(0, 8),
540 => conv_std_logic_vector(0, 8),
541 => conv_std_logic_vector(0, 8),
542 => conv_std_logic_vector(0, 8),
543 => conv_std_logic_vector(0, 8),
544 => conv_std_logic_vector(0, 8),
545 => conv_std_logic_vector(0, 8),
546 => conv_std_logic_vector(0, 8),
547 => conv_std_logic_vector(0, 8),
548 => conv_std_logic_vector(0, 8),
549 => conv_std_logic_vector(0, 8),
550 => conv_std_logic_vector(0, 8),
551 => conv_std_logic_vector(0, 8),
552 => conv_std_logic_vector(0, 8),
553 => conv_std_logic_vector(0, 8),
554 => conv_std_logic_vector(0, 8),
555 => conv_std_logic_vector(0, 8),
556 => conv_std_logic_vector(0, 8),
557 => conv_std_logic_vector(0, 8),
558 => conv_std_logic_vector(0, 8),
559 => conv_std_logic_vector(0, 8),
560 => conv_std_logic_vector(0, 8),
561 => conv_std_logic_vector(0, 8),
562 => conv_std_logic_vector(0, 8),
563 => conv_std_logic_vector(0, 8),
564 => conv_std_logic_vector(0, 8),
565 => conv_std_logic_vector(0, 8),
566 => conv_std_logic_vector(0, 8),
567 => conv_std_logic_vector(0, 8),
568 => conv_std_logic_vector(0, 8),
569 => conv_std_logic_vector(0, 8),
570 => conv_std_logic_vector(0, 8),
571 => conv_std_logic_vector(0, 8),
572 => conv_std_logic_vector(0, 8),
573 => conv_std_logic_vector(0, 8),
574 => conv_std_logic_vector(0, 8),
575 => conv_std_logic_vector(0, 8),
576 => conv_std_logic_vector(0, 8),
577 => conv_std_logic_vector(0, 8),
578 => conv_std_logic_vector(0, 8),
579 => conv_std_logic_vector(0, 8),
580 => conv_std_logic_vector(0, 8),
581 => conv_std_logic_vector(0, 8),
582 => conv_std_logic_vector(0, 8),
583 => conv_std_logic_vector(0, 8),
584 => conv_std_logic_vector(0, 8),
585 => conv_std_logic_vector(0, 8),
586 => conv_std_logic_vector(0, 8),
587 => conv_std_logic_vector(0, 8),
588 => conv_std_logic_vector(0, 8),
589 => conv_std_logic_vector(0, 8),
590 => conv_std_logic_vector(0, 8),
591 => conv_std_logic_vector(0, 8),
592 => conv_std_logic_vector(0, 8),
593 => conv_std_logic_vector(0, 8),
594 => conv_std_logic_vector(0, 8),
595 => conv_std_logic_vector(0, 8),
596 => conv_std_logic_vector(0, 8),
597 => conv_std_logic_vector(0, 8),
598 => conv_std_logic_vector(0, 8),
599 => conv_std_logic_vector(0, 8),
600 => conv_std_logic_vector(0, 8),
601 => conv_std_logic_vector(0, 8),
602 => conv_std_logic_vector(0, 8),
603 => conv_std_logic_vector(0, 8),
604 => conv_std_logic_vector(0, 8),
605 => conv_std_logic_vector(0, 8),
606 => conv_std_logic_vector(0, 8),
607 => conv_std_logic_vector(0, 8),
608 => conv_std_logic_vector(0, 8),
609 => conv_std_logic_vector(0, 8),
610 => conv_std_logic_vector(0, 8),
611 => conv_std_logic_vector(0, 8),
612 => conv_std_logic_vector(0, 8),
613 => conv_std_logic_vector(0, 8),
614 => conv_std_logic_vector(0, 8),
615 => conv_std_logic_vector(0, 8),
616 => conv_std_logic_vector(0, 8),
617 => conv_std_logic_vector(0, 8),
618 => conv_std_logic_vector(0, 8),
619 => conv_std_logic_vector(0, 8),
620 => conv_std_logic_vector(0, 8),
621 => conv_std_logic_vector(0, 8),
622 => conv_std_logic_vector(0, 8),
623 => conv_std_logic_vector(0, 8),
624 => conv_std_logic_vector(0, 8),
625 => conv_std_logic_vector(0, 8),
626 => conv_std_logic_vector(0, 8),
627 => conv_std_logic_vector(0, 8),
628 => conv_std_logic_vector(0, 8),
629 => conv_std_logic_vector(0, 8),
630 => conv_std_logic_vector(0, 8),
631 => conv_std_logic_vector(0, 8),
632 => conv_std_logic_vector(0, 8),
633 => conv_std_logic_vector(0, 8),
634 => conv_std_logic_vector(0, 8),
635 => conv_std_logic_vector(0, 8),
636 => conv_std_logic_vector(0, 8),
637 => conv_std_logic_vector(0, 8),
638 => conv_std_logic_vector(0, 8),
639 => conv_std_logic_vector(0, 8),
640 => conv_std_logic_vector(1, 8),
641 => conv_std_logic_vector(1, 8),
642 => conv_std_logic_vector(1, 8),
643 => conv_std_logic_vector(1, 8),
644 => conv_std_logic_vector(1, 8),
645 => conv_std_logic_vector(1, 8),
646 => conv_std_logic_vector(1, 8),
647 => conv_std_logic_vector(1, 8),
648 => conv_std_logic_vector(1, 8),
649 => conv_std_logic_vector(1, 8),
650 => conv_std_logic_vector(1, 8),
651 => conv_std_logic_vector(1, 8),
652 => conv_std_logic_vector(1, 8),
653 => conv_std_logic_vector(1, 8),
654 => conv_std_logic_vector(1, 8),
655 => conv_std_logic_vector(1, 8),
656 => conv_std_logic_vector(1, 8),
657 => conv_std_logic_vector(1, 8),
658 => conv_std_logic_vector(1, 8),
659 => conv_std_logic_vector(1, 8),
660 => conv_std_logic_vector(1, 8),
661 => conv_std_logic_vector(1, 8),
662 => conv_std_logic_vector(1, 8),
663 => conv_std_logic_vector(1, 8),
664 => conv_std_logic_vector(1, 8),
665 => conv_std_logic_vector(1, 8),
666 => conv_std_logic_vector(1, 8),
667 => conv_std_logic_vector(1, 8),
668 => conv_std_logic_vector(1, 8),
669 => conv_std_logic_vector(1, 8),
670 => conv_std_logic_vector(1, 8),
671 => conv_std_logic_vector(1, 8),
672 => conv_std_logic_vector(1, 8),
673 => conv_std_logic_vector(1, 8),
674 => conv_std_logic_vector(1, 8),
675 => conv_std_logic_vector(1, 8),
676 => conv_std_logic_vector(1, 8),
677 => conv_std_logic_vector(1, 8),
678 => conv_std_logic_vector(1, 8),
679 => conv_std_logic_vector(1, 8),
680 => conv_std_logic_vector(1, 8),
681 => conv_std_logic_vector(1, 8),
682 => conv_std_logic_vector(1, 8),
683 => conv_std_logic_vector(1, 8),
684 => conv_std_logic_vector(1, 8),
685 => conv_std_logic_vector(1, 8),
686 => conv_std_logic_vector(1, 8),
687 => conv_std_logic_vector(1, 8),
688 => conv_std_logic_vector(1, 8),
689 => conv_std_logic_vector(1, 8),
690 => conv_std_logic_vector(1, 8),
691 => conv_std_logic_vector(1, 8),
692 => conv_std_logic_vector(1, 8),
693 => conv_std_logic_vector(1, 8),
694 => conv_std_logic_vector(1, 8),
695 => conv_std_logic_vector(1, 8),
696 => conv_std_logic_vector(1, 8),
697 => conv_std_logic_vector(1, 8),
698 => conv_std_logic_vector(1, 8),
699 => conv_std_logic_vector(1, 8),
700 => conv_std_logic_vector(1, 8),
701 => conv_std_logic_vector(1, 8),
702 => conv_std_logic_vector(1, 8),
703 => conv_std_logic_vector(1, 8),
704 => conv_std_logic_vector(1, 8),
705 => conv_std_logic_vector(1, 8),
706 => conv_std_logic_vector(1, 8),
707 => conv_std_logic_vector(1, 8),
708 => conv_std_logic_vector(1, 8),
709 => conv_std_logic_vector(1, 8),
710 => conv_std_logic_vector(1, 8),
711 => conv_std_logic_vector(1, 8),
712 => conv_std_logic_vector(1, 8),
713 => conv_std_logic_vector(1, 8),
714 => conv_std_logic_vector(1, 8),
715 => conv_std_logic_vector(1, 8),
716 => conv_std_logic_vector(1, 8),
717 => conv_std_logic_vector(1, 8),
718 => conv_std_logic_vector(1, 8),
719 => conv_std_logic_vector(1, 8),
720 => conv_std_logic_vector(1, 8),
721 => conv_std_logic_vector(1, 8),
722 => conv_std_logic_vector(1, 8),
723 => conv_std_logic_vector(1, 8),
724 => conv_std_logic_vector(1, 8),
725 => conv_std_logic_vector(1, 8),
726 => conv_std_logic_vector(1, 8),
727 => conv_std_logic_vector(1, 8),
728 => conv_std_logic_vector(1, 8),
729 => conv_std_logic_vector(1, 8),
730 => conv_std_logic_vector(1, 8),
731 => conv_std_logic_vector(1, 8),
732 => conv_std_logic_vector(1, 8),
733 => conv_std_logic_vector(1, 8),
734 => conv_std_logic_vector(1, 8),
735 => conv_std_logic_vector(1, 8),
736 => conv_std_logic_vector(1, 8),
737 => conv_std_logic_vector(1, 8),
738 => conv_std_logic_vector(1, 8),
739 => conv_std_logic_vector(1, 8),
740 => conv_std_logic_vector(1, 8),
741 => conv_std_logic_vector(1, 8),
742 => conv_std_logic_vector(1, 8),
743 => conv_std_logic_vector(1, 8),
744 => conv_std_logic_vector(1, 8),
745 => conv_std_logic_vector(1, 8),
746 => conv_std_logic_vector(1, 8),
747 => conv_std_logic_vector(1, 8),
748 => conv_std_logic_vector(1, 8),
749 => conv_std_logic_vector(1, 8),
750 => conv_std_logic_vector(1, 8),
751 => conv_std_logic_vector(1, 8),
752 => conv_std_logic_vector(1, 8),
753 => conv_std_logic_vector(1, 8),
754 => conv_std_logic_vector(1, 8),
755 => conv_std_logic_vector(1, 8),
756 => conv_std_logic_vector(1, 8),
757 => conv_std_logic_vector(1, 8),
758 => conv_std_logic_vector(1, 8),
759 => conv_std_logic_vector(1, 8),
760 => conv_std_logic_vector(1, 8),
761 => conv_std_logic_vector(1, 8),
762 => conv_std_logic_vector(1, 8),
763 => conv_std_logic_vector(1, 8),
764 => conv_std_logic_vector(1, 8),
765 => conv_std_logic_vector(1, 8),
766 => conv_std_logic_vector(1, 8),
767 => conv_std_logic_vector(1, 8),
768 => conv_std_logic_vector(0, 8),
769 => conv_std_logic_vector(0, 8),
770 => conv_std_logic_vector(0, 8),
771 => conv_std_logic_vector(0, 8),
772 => conv_std_logic_vector(0, 8),
773 => conv_std_logic_vector(0, 8),
774 => conv_std_logic_vector(0, 8),
775 => conv_std_logic_vector(0, 8),
776 => conv_std_logic_vector(0, 8),
777 => conv_std_logic_vector(0, 8),
778 => conv_std_logic_vector(0, 8),
779 => conv_std_logic_vector(0, 8),
780 => conv_std_logic_vector(0, 8),
781 => conv_std_logic_vector(0, 8),
782 => conv_std_logic_vector(0, 8),
783 => conv_std_logic_vector(0, 8),
784 => conv_std_logic_vector(0, 8),
785 => conv_std_logic_vector(0, 8),
786 => conv_std_logic_vector(0, 8),
787 => conv_std_logic_vector(0, 8),
788 => conv_std_logic_vector(0, 8),
789 => conv_std_logic_vector(0, 8),
790 => conv_std_logic_vector(0, 8),
791 => conv_std_logic_vector(0, 8),
792 => conv_std_logic_vector(0, 8),
793 => conv_std_logic_vector(0, 8),
794 => conv_std_logic_vector(0, 8),
795 => conv_std_logic_vector(0, 8),
796 => conv_std_logic_vector(0, 8),
797 => conv_std_logic_vector(0, 8),
798 => conv_std_logic_vector(0, 8),
799 => conv_std_logic_vector(0, 8),
800 => conv_std_logic_vector(0, 8),
801 => conv_std_logic_vector(0, 8),
802 => conv_std_logic_vector(0, 8),
803 => conv_std_logic_vector(0, 8),
804 => conv_std_logic_vector(0, 8),
805 => conv_std_logic_vector(0, 8),
806 => conv_std_logic_vector(0, 8),
807 => conv_std_logic_vector(0, 8),
808 => conv_std_logic_vector(0, 8),
809 => conv_std_logic_vector(0, 8),
810 => conv_std_logic_vector(0, 8),
811 => conv_std_logic_vector(0, 8),
812 => conv_std_logic_vector(0, 8),
813 => conv_std_logic_vector(0, 8),
814 => conv_std_logic_vector(0, 8),
815 => conv_std_logic_vector(0, 8),
816 => conv_std_logic_vector(0, 8),
817 => conv_std_logic_vector(0, 8),
818 => conv_std_logic_vector(0, 8),
819 => conv_std_logic_vector(0, 8),
820 => conv_std_logic_vector(0, 8),
821 => conv_std_logic_vector(0, 8),
822 => conv_std_logic_vector(0, 8),
823 => conv_std_logic_vector(0, 8),
824 => conv_std_logic_vector(0, 8),
825 => conv_std_logic_vector(0, 8),
826 => conv_std_logic_vector(0, 8),
827 => conv_std_logic_vector(0, 8),
828 => conv_std_logic_vector(0, 8),
829 => conv_std_logic_vector(0, 8),
830 => conv_std_logic_vector(0, 8),
831 => conv_std_logic_vector(0, 8),
832 => conv_std_logic_vector(0, 8),
833 => conv_std_logic_vector(0, 8),
834 => conv_std_logic_vector(0, 8),
835 => conv_std_logic_vector(0, 8),
836 => conv_std_logic_vector(0, 8),
837 => conv_std_logic_vector(0, 8),
838 => conv_std_logic_vector(0, 8),
839 => conv_std_logic_vector(0, 8),
840 => conv_std_logic_vector(0, 8),
841 => conv_std_logic_vector(0, 8),
842 => conv_std_logic_vector(0, 8),
843 => conv_std_logic_vector(0, 8),
844 => conv_std_logic_vector(0, 8),
845 => conv_std_logic_vector(0, 8),
846 => conv_std_logic_vector(0, 8),
847 => conv_std_logic_vector(0, 8),
848 => conv_std_logic_vector(0, 8),
849 => conv_std_logic_vector(0, 8),
850 => conv_std_logic_vector(0, 8),
851 => conv_std_logic_vector(0, 8),
852 => conv_std_logic_vector(0, 8),
853 => conv_std_logic_vector(0, 8),
854 => conv_std_logic_vector(1, 8),
855 => conv_std_logic_vector(1, 8),
856 => conv_std_logic_vector(1, 8),
857 => conv_std_logic_vector(1, 8),
858 => conv_std_logic_vector(1, 8),
859 => conv_std_logic_vector(1, 8),
860 => conv_std_logic_vector(1, 8),
861 => conv_std_logic_vector(1, 8),
862 => conv_std_logic_vector(1, 8),
863 => conv_std_logic_vector(1, 8),
864 => conv_std_logic_vector(1, 8),
865 => conv_std_logic_vector(1, 8),
866 => conv_std_logic_vector(1, 8),
867 => conv_std_logic_vector(1, 8),
868 => conv_std_logic_vector(1, 8),
869 => conv_std_logic_vector(1, 8),
870 => conv_std_logic_vector(1, 8),
871 => conv_std_logic_vector(1, 8),
872 => conv_std_logic_vector(1, 8),
873 => conv_std_logic_vector(1, 8),
874 => conv_std_logic_vector(1, 8),
875 => conv_std_logic_vector(1, 8),
876 => conv_std_logic_vector(1, 8),
877 => conv_std_logic_vector(1, 8),
878 => conv_std_logic_vector(1, 8),
879 => conv_std_logic_vector(1, 8),
880 => conv_std_logic_vector(1, 8),
881 => conv_std_logic_vector(1, 8),
882 => conv_std_logic_vector(1, 8),
883 => conv_std_logic_vector(1, 8),
884 => conv_std_logic_vector(1, 8),
885 => conv_std_logic_vector(1, 8),
886 => conv_std_logic_vector(1, 8),
887 => conv_std_logic_vector(1, 8),
888 => conv_std_logic_vector(1, 8),
889 => conv_std_logic_vector(1, 8),
890 => conv_std_logic_vector(1, 8),
891 => conv_std_logic_vector(1, 8),
892 => conv_std_logic_vector(1, 8),
893 => conv_std_logic_vector(1, 8),
894 => conv_std_logic_vector(1, 8),
895 => conv_std_logic_vector(1, 8),
896 => conv_std_logic_vector(1, 8),
897 => conv_std_logic_vector(1, 8),
898 => conv_std_logic_vector(1, 8),
899 => conv_std_logic_vector(1, 8),
900 => conv_std_logic_vector(1, 8),
901 => conv_std_logic_vector(1, 8),
902 => conv_std_logic_vector(1, 8),
903 => conv_std_logic_vector(1, 8),
904 => conv_std_logic_vector(1, 8),
905 => conv_std_logic_vector(1, 8),
906 => conv_std_logic_vector(1, 8),
907 => conv_std_logic_vector(1, 8),
908 => conv_std_logic_vector(1, 8),
909 => conv_std_logic_vector(1, 8),
910 => conv_std_logic_vector(1, 8),
911 => conv_std_logic_vector(1, 8),
912 => conv_std_logic_vector(1, 8),
913 => conv_std_logic_vector(1, 8),
914 => conv_std_logic_vector(1, 8),
915 => conv_std_logic_vector(1, 8),
916 => conv_std_logic_vector(1, 8),
917 => conv_std_logic_vector(1, 8),
918 => conv_std_logic_vector(1, 8),
919 => conv_std_logic_vector(1, 8),
920 => conv_std_logic_vector(1, 8),
921 => conv_std_logic_vector(1, 8),
922 => conv_std_logic_vector(1, 8),
923 => conv_std_logic_vector(1, 8),
924 => conv_std_logic_vector(1, 8),
925 => conv_std_logic_vector(1, 8),
926 => conv_std_logic_vector(1, 8),
927 => conv_std_logic_vector(1, 8),
928 => conv_std_logic_vector(1, 8),
929 => conv_std_logic_vector(1, 8),
930 => conv_std_logic_vector(1, 8),
931 => conv_std_logic_vector(1, 8),
932 => conv_std_logic_vector(1, 8),
933 => conv_std_logic_vector(1, 8),
934 => conv_std_logic_vector(1, 8),
935 => conv_std_logic_vector(1, 8),
936 => conv_std_logic_vector(1, 8),
937 => conv_std_logic_vector(1, 8),
938 => conv_std_logic_vector(1, 8),
939 => conv_std_logic_vector(2, 8),
940 => conv_std_logic_vector(2, 8),
941 => conv_std_logic_vector(2, 8),
942 => conv_std_logic_vector(2, 8),
943 => conv_std_logic_vector(2, 8),
944 => conv_std_logic_vector(2, 8),
945 => conv_std_logic_vector(2, 8),
946 => conv_std_logic_vector(2, 8),
947 => conv_std_logic_vector(2, 8),
948 => conv_std_logic_vector(2, 8),
949 => conv_std_logic_vector(2, 8),
950 => conv_std_logic_vector(2, 8),
951 => conv_std_logic_vector(2, 8),
952 => conv_std_logic_vector(2, 8),
953 => conv_std_logic_vector(2, 8),
954 => conv_std_logic_vector(2, 8),
955 => conv_std_logic_vector(2, 8),
956 => conv_std_logic_vector(2, 8),
957 => conv_std_logic_vector(2, 8),
958 => conv_std_logic_vector(2, 8),
959 => conv_std_logic_vector(2, 8),
960 => conv_std_logic_vector(2, 8),
961 => conv_std_logic_vector(2, 8),
962 => conv_std_logic_vector(2, 8),
963 => conv_std_logic_vector(2, 8),
964 => conv_std_logic_vector(2, 8),
965 => conv_std_logic_vector(2, 8),
966 => conv_std_logic_vector(2, 8),
967 => conv_std_logic_vector(2, 8),
968 => conv_std_logic_vector(2, 8),
969 => conv_std_logic_vector(2, 8),
970 => conv_std_logic_vector(2, 8),
971 => conv_std_logic_vector(2, 8),
972 => conv_std_logic_vector(2, 8),
973 => conv_std_logic_vector(2, 8),
974 => conv_std_logic_vector(2, 8),
975 => conv_std_logic_vector(2, 8),
976 => conv_std_logic_vector(2, 8),
977 => conv_std_logic_vector(2, 8),
978 => conv_std_logic_vector(2, 8),
979 => conv_std_logic_vector(2, 8),
980 => conv_std_logic_vector(2, 8),
981 => conv_std_logic_vector(2, 8),
982 => conv_std_logic_vector(2, 8),
983 => conv_std_logic_vector(2, 8),
984 => conv_std_logic_vector(2, 8),
985 => conv_std_logic_vector(2, 8),
986 => conv_std_logic_vector(2, 8),
987 => conv_std_logic_vector(2, 8),
988 => conv_std_logic_vector(2, 8),
989 => conv_std_logic_vector(2, 8),
990 => conv_std_logic_vector(2, 8),
991 => conv_std_logic_vector(2, 8),
992 => conv_std_logic_vector(2, 8),
993 => conv_std_logic_vector(2, 8),
994 => conv_std_logic_vector(2, 8),
995 => conv_std_logic_vector(2, 8),
996 => conv_std_logic_vector(2, 8),
997 => conv_std_logic_vector(2, 8),
998 => conv_std_logic_vector(2, 8),
999 => conv_std_logic_vector(2, 8),
1000 => conv_std_logic_vector(2, 8),
1001 => conv_std_logic_vector(2, 8),
1002 => conv_std_logic_vector(2, 8),
1003 => conv_std_logic_vector(2, 8),
1004 => conv_std_logic_vector(2, 8),
1005 => conv_std_logic_vector(2, 8),
1006 => conv_std_logic_vector(2, 8),
1007 => conv_std_logic_vector(2, 8),
1008 => conv_std_logic_vector(2, 8),
1009 => conv_std_logic_vector(2, 8),
1010 => conv_std_logic_vector(2, 8),
1011 => conv_std_logic_vector(2, 8),
1012 => conv_std_logic_vector(2, 8),
1013 => conv_std_logic_vector(2, 8),
1014 => conv_std_logic_vector(2, 8),
1015 => conv_std_logic_vector(2, 8),
1016 => conv_std_logic_vector(2, 8),
1017 => conv_std_logic_vector(2, 8),
1018 => conv_std_logic_vector(2, 8),
1019 => conv_std_logic_vector(2, 8),
1020 => conv_std_logic_vector(2, 8),
1021 => conv_std_logic_vector(2, 8),
1022 => conv_std_logic_vector(2, 8),
1023 => conv_std_logic_vector(2, 8),
1024 => conv_std_logic_vector(0, 8),
1025 => conv_std_logic_vector(0, 8),
1026 => conv_std_logic_vector(0, 8),
1027 => conv_std_logic_vector(0, 8),
1028 => conv_std_logic_vector(0, 8),
1029 => conv_std_logic_vector(0, 8),
1030 => conv_std_logic_vector(0, 8),
1031 => conv_std_logic_vector(0, 8),
1032 => conv_std_logic_vector(0, 8),
1033 => conv_std_logic_vector(0, 8),
1034 => conv_std_logic_vector(0, 8),
1035 => conv_std_logic_vector(0, 8),
1036 => conv_std_logic_vector(0, 8),
1037 => conv_std_logic_vector(0, 8),
1038 => conv_std_logic_vector(0, 8),
1039 => conv_std_logic_vector(0, 8),
1040 => conv_std_logic_vector(0, 8),
1041 => conv_std_logic_vector(0, 8),
1042 => conv_std_logic_vector(0, 8),
1043 => conv_std_logic_vector(0, 8),
1044 => conv_std_logic_vector(0, 8),
1045 => conv_std_logic_vector(0, 8),
1046 => conv_std_logic_vector(0, 8),
1047 => conv_std_logic_vector(0, 8),
1048 => conv_std_logic_vector(0, 8),
1049 => conv_std_logic_vector(0, 8),
1050 => conv_std_logic_vector(0, 8),
1051 => conv_std_logic_vector(0, 8),
1052 => conv_std_logic_vector(0, 8),
1053 => conv_std_logic_vector(0, 8),
1054 => conv_std_logic_vector(0, 8),
1055 => conv_std_logic_vector(0, 8),
1056 => conv_std_logic_vector(0, 8),
1057 => conv_std_logic_vector(0, 8),
1058 => conv_std_logic_vector(0, 8),
1059 => conv_std_logic_vector(0, 8),
1060 => conv_std_logic_vector(0, 8),
1061 => conv_std_logic_vector(0, 8),
1062 => conv_std_logic_vector(0, 8),
1063 => conv_std_logic_vector(0, 8),
1064 => conv_std_logic_vector(0, 8),
1065 => conv_std_logic_vector(0, 8),
1066 => conv_std_logic_vector(0, 8),
1067 => conv_std_logic_vector(0, 8),
1068 => conv_std_logic_vector(0, 8),
1069 => conv_std_logic_vector(0, 8),
1070 => conv_std_logic_vector(0, 8),
1071 => conv_std_logic_vector(0, 8),
1072 => conv_std_logic_vector(0, 8),
1073 => conv_std_logic_vector(0, 8),
1074 => conv_std_logic_vector(0, 8),
1075 => conv_std_logic_vector(0, 8),
1076 => conv_std_logic_vector(0, 8),
1077 => conv_std_logic_vector(0, 8),
1078 => conv_std_logic_vector(0, 8),
1079 => conv_std_logic_vector(0, 8),
1080 => conv_std_logic_vector(0, 8),
1081 => conv_std_logic_vector(0, 8),
1082 => conv_std_logic_vector(0, 8),
1083 => conv_std_logic_vector(0, 8),
1084 => conv_std_logic_vector(0, 8),
1085 => conv_std_logic_vector(0, 8),
1086 => conv_std_logic_vector(0, 8),
1087 => conv_std_logic_vector(0, 8),
1088 => conv_std_logic_vector(1, 8),
1089 => conv_std_logic_vector(1, 8),
1090 => conv_std_logic_vector(1, 8),
1091 => conv_std_logic_vector(1, 8),
1092 => conv_std_logic_vector(1, 8),
1093 => conv_std_logic_vector(1, 8),
1094 => conv_std_logic_vector(1, 8),
1095 => conv_std_logic_vector(1, 8),
1096 => conv_std_logic_vector(1, 8),
1097 => conv_std_logic_vector(1, 8),
1098 => conv_std_logic_vector(1, 8),
1099 => conv_std_logic_vector(1, 8),
1100 => conv_std_logic_vector(1, 8),
1101 => conv_std_logic_vector(1, 8),
1102 => conv_std_logic_vector(1, 8),
1103 => conv_std_logic_vector(1, 8),
1104 => conv_std_logic_vector(1, 8),
1105 => conv_std_logic_vector(1, 8),
1106 => conv_std_logic_vector(1, 8),
1107 => conv_std_logic_vector(1, 8),
1108 => conv_std_logic_vector(1, 8),
1109 => conv_std_logic_vector(1, 8),
1110 => conv_std_logic_vector(1, 8),
1111 => conv_std_logic_vector(1, 8),
1112 => conv_std_logic_vector(1, 8),
1113 => conv_std_logic_vector(1, 8),
1114 => conv_std_logic_vector(1, 8),
1115 => conv_std_logic_vector(1, 8),
1116 => conv_std_logic_vector(1, 8),
1117 => conv_std_logic_vector(1, 8),
1118 => conv_std_logic_vector(1, 8),
1119 => conv_std_logic_vector(1, 8),
1120 => conv_std_logic_vector(1, 8),
1121 => conv_std_logic_vector(1, 8),
1122 => conv_std_logic_vector(1, 8),
1123 => conv_std_logic_vector(1, 8),
1124 => conv_std_logic_vector(1, 8),
1125 => conv_std_logic_vector(1, 8),
1126 => conv_std_logic_vector(1, 8),
1127 => conv_std_logic_vector(1, 8),
1128 => conv_std_logic_vector(1, 8),
1129 => conv_std_logic_vector(1, 8),
1130 => conv_std_logic_vector(1, 8),
1131 => conv_std_logic_vector(1, 8),
1132 => conv_std_logic_vector(1, 8),
1133 => conv_std_logic_vector(1, 8),
1134 => conv_std_logic_vector(1, 8),
1135 => conv_std_logic_vector(1, 8),
1136 => conv_std_logic_vector(1, 8),
1137 => conv_std_logic_vector(1, 8),
1138 => conv_std_logic_vector(1, 8),
1139 => conv_std_logic_vector(1, 8),
1140 => conv_std_logic_vector(1, 8),
1141 => conv_std_logic_vector(1, 8),
1142 => conv_std_logic_vector(1, 8),
1143 => conv_std_logic_vector(1, 8),
1144 => conv_std_logic_vector(1, 8),
1145 => conv_std_logic_vector(1, 8),
1146 => conv_std_logic_vector(1, 8),
1147 => conv_std_logic_vector(1, 8),
1148 => conv_std_logic_vector(1, 8),
1149 => conv_std_logic_vector(1, 8),
1150 => conv_std_logic_vector(1, 8),
1151 => conv_std_logic_vector(1, 8),
1152 => conv_std_logic_vector(2, 8),
1153 => conv_std_logic_vector(2, 8),
1154 => conv_std_logic_vector(2, 8),
1155 => conv_std_logic_vector(2, 8),
1156 => conv_std_logic_vector(2, 8),
1157 => conv_std_logic_vector(2, 8),
1158 => conv_std_logic_vector(2, 8),
1159 => conv_std_logic_vector(2, 8),
1160 => conv_std_logic_vector(2, 8),
1161 => conv_std_logic_vector(2, 8),
1162 => conv_std_logic_vector(2, 8),
1163 => conv_std_logic_vector(2, 8),
1164 => conv_std_logic_vector(2, 8),
1165 => conv_std_logic_vector(2, 8),
1166 => conv_std_logic_vector(2, 8),
1167 => conv_std_logic_vector(2, 8),
1168 => conv_std_logic_vector(2, 8),
1169 => conv_std_logic_vector(2, 8),
1170 => conv_std_logic_vector(2, 8),
1171 => conv_std_logic_vector(2, 8),
1172 => conv_std_logic_vector(2, 8),
1173 => conv_std_logic_vector(2, 8),
1174 => conv_std_logic_vector(2, 8),
1175 => conv_std_logic_vector(2, 8),
1176 => conv_std_logic_vector(2, 8),
1177 => conv_std_logic_vector(2, 8),
1178 => conv_std_logic_vector(2, 8),
1179 => conv_std_logic_vector(2, 8),
1180 => conv_std_logic_vector(2, 8),
1181 => conv_std_logic_vector(2, 8),
1182 => conv_std_logic_vector(2, 8),
1183 => conv_std_logic_vector(2, 8),
1184 => conv_std_logic_vector(2, 8),
1185 => conv_std_logic_vector(2, 8),
1186 => conv_std_logic_vector(2, 8),
1187 => conv_std_logic_vector(2, 8),
1188 => conv_std_logic_vector(2, 8),
1189 => conv_std_logic_vector(2, 8),
1190 => conv_std_logic_vector(2, 8),
1191 => conv_std_logic_vector(2, 8),
1192 => conv_std_logic_vector(2, 8),
1193 => conv_std_logic_vector(2, 8),
1194 => conv_std_logic_vector(2, 8),
1195 => conv_std_logic_vector(2, 8),
1196 => conv_std_logic_vector(2, 8),
1197 => conv_std_logic_vector(2, 8),
1198 => conv_std_logic_vector(2, 8),
1199 => conv_std_logic_vector(2, 8),
1200 => conv_std_logic_vector(2, 8),
1201 => conv_std_logic_vector(2, 8),
1202 => conv_std_logic_vector(2, 8),
1203 => conv_std_logic_vector(2, 8),
1204 => conv_std_logic_vector(2, 8),
1205 => conv_std_logic_vector(2, 8),
1206 => conv_std_logic_vector(2, 8),
1207 => conv_std_logic_vector(2, 8),
1208 => conv_std_logic_vector(2, 8),
1209 => conv_std_logic_vector(2, 8),
1210 => conv_std_logic_vector(2, 8),
1211 => conv_std_logic_vector(2, 8),
1212 => conv_std_logic_vector(2, 8),
1213 => conv_std_logic_vector(2, 8),
1214 => conv_std_logic_vector(2, 8),
1215 => conv_std_logic_vector(2, 8),
1216 => conv_std_logic_vector(3, 8),
1217 => conv_std_logic_vector(3, 8),
1218 => conv_std_logic_vector(3, 8),
1219 => conv_std_logic_vector(3, 8),
1220 => conv_std_logic_vector(3, 8),
1221 => conv_std_logic_vector(3, 8),
1222 => conv_std_logic_vector(3, 8),
1223 => conv_std_logic_vector(3, 8),
1224 => conv_std_logic_vector(3, 8),
1225 => conv_std_logic_vector(3, 8),
1226 => conv_std_logic_vector(3, 8),
1227 => conv_std_logic_vector(3, 8),
1228 => conv_std_logic_vector(3, 8),
1229 => conv_std_logic_vector(3, 8),
1230 => conv_std_logic_vector(3, 8),
1231 => conv_std_logic_vector(3, 8),
1232 => conv_std_logic_vector(3, 8),
1233 => conv_std_logic_vector(3, 8),
1234 => conv_std_logic_vector(3, 8),
1235 => conv_std_logic_vector(3, 8),
1236 => conv_std_logic_vector(3, 8),
1237 => conv_std_logic_vector(3, 8),
1238 => conv_std_logic_vector(3, 8),
1239 => conv_std_logic_vector(3, 8),
1240 => conv_std_logic_vector(3, 8),
1241 => conv_std_logic_vector(3, 8),
1242 => conv_std_logic_vector(3, 8),
1243 => conv_std_logic_vector(3, 8),
1244 => conv_std_logic_vector(3, 8),
1245 => conv_std_logic_vector(3, 8),
1246 => conv_std_logic_vector(3, 8),
1247 => conv_std_logic_vector(3, 8),
1248 => conv_std_logic_vector(3, 8),
1249 => conv_std_logic_vector(3, 8),
1250 => conv_std_logic_vector(3, 8),
1251 => conv_std_logic_vector(3, 8),
1252 => conv_std_logic_vector(3, 8),
1253 => conv_std_logic_vector(3, 8),
1254 => conv_std_logic_vector(3, 8),
1255 => conv_std_logic_vector(3, 8),
1256 => conv_std_logic_vector(3, 8),
1257 => conv_std_logic_vector(3, 8),
1258 => conv_std_logic_vector(3, 8),
1259 => conv_std_logic_vector(3, 8),
1260 => conv_std_logic_vector(3, 8),
1261 => conv_std_logic_vector(3, 8),
1262 => conv_std_logic_vector(3, 8),
1263 => conv_std_logic_vector(3, 8),
1264 => conv_std_logic_vector(3, 8),
1265 => conv_std_logic_vector(3, 8),
1266 => conv_std_logic_vector(3, 8),
1267 => conv_std_logic_vector(3, 8),
1268 => conv_std_logic_vector(3, 8),
1269 => conv_std_logic_vector(3, 8),
1270 => conv_std_logic_vector(3, 8),
1271 => conv_std_logic_vector(3, 8),
1272 => conv_std_logic_vector(3, 8),
1273 => conv_std_logic_vector(3, 8),
1274 => conv_std_logic_vector(3, 8),
1275 => conv_std_logic_vector(3, 8),
1276 => conv_std_logic_vector(3, 8),
1277 => conv_std_logic_vector(3, 8),
1278 => conv_std_logic_vector(3, 8),
1279 => conv_std_logic_vector(3, 8),
1280 => conv_std_logic_vector(0, 8),
1281 => conv_std_logic_vector(0, 8),
1282 => conv_std_logic_vector(0, 8),
1283 => conv_std_logic_vector(0, 8),
1284 => conv_std_logic_vector(0, 8),
1285 => conv_std_logic_vector(0, 8),
1286 => conv_std_logic_vector(0, 8),
1287 => conv_std_logic_vector(0, 8),
1288 => conv_std_logic_vector(0, 8),
1289 => conv_std_logic_vector(0, 8),
1290 => conv_std_logic_vector(0, 8),
1291 => conv_std_logic_vector(0, 8),
1292 => conv_std_logic_vector(0, 8),
1293 => conv_std_logic_vector(0, 8),
1294 => conv_std_logic_vector(0, 8),
1295 => conv_std_logic_vector(0, 8),
1296 => conv_std_logic_vector(0, 8),
1297 => conv_std_logic_vector(0, 8),
1298 => conv_std_logic_vector(0, 8),
1299 => conv_std_logic_vector(0, 8),
1300 => conv_std_logic_vector(0, 8),
1301 => conv_std_logic_vector(0, 8),
1302 => conv_std_logic_vector(0, 8),
1303 => conv_std_logic_vector(0, 8),
1304 => conv_std_logic_vector(0, 8),
1305 => conv_std_logic_vector(0, 8),
1306 => conv_std_logic_vector(0, 8),
1307 => conv_std_logic_vector(0, 8),
1308 => conv_std_logic_vector(0, 8),
1309 => conv_std_logic_vector(0, 8),
1310 => conv_std_logic_vector(0, 8),
1311 => conv_std_logic_vector(0, 8),
1312 => conv_std_logic_vector(0, 8),
1313 => conv_std_logic_vector(0, 8),
1314 => conv_std_logic_vector(0, 8),
1315 => conv_std_logic_vector(0, 8),
1316 => conv_std_logic_vector(0, 8),
1317 => conv_std_logic_vector(0, 8),
1318 => conv_std_logic_vector(0, 8),
1319 => conv_std_logic_vector(0, 8),
1320 => conv_std_logic_vector(0, 8),
1321 => conv_std_logic_vector(0, 8),
1322 => conv_std_logic_vector(0, 8),
1323 => conv_std_logic_vector(0, 8),
1324 => conv_std_logic_vector(0, 8),
1325 => conv_std_logic_vector(0, 8),
1326 => conv_std_logic_vector(0, 8),
1327 => conv_std_logic_vector(0, 8),
1328 => conv_std_logic_vector(0, 8),
1329 => conv_std_logic_vector(0, 8),
1330 => conv_std_logic_vector(0, 8),
1331 => conv_std_logic_vector(0, 8),
1332 => conv_std_logic_vector(1, 8),
1333 => conv_std_logic_vector(1, 8),
1334 => conv_std_logic_vector(1, 8),
1335 => conv_std_logic_vector(1, 8),
1336 => conv_std_logic_vector(1, 8),
1337 => conv_std_logic_vector(1, 8),
1338 => conv_std_logic_vector(1, 8),
1339 => conv_std_logic_vector(1, 8),
1340 => conv_std_logic_vector(1, 8),
1341 => conv_std_logic_vector(1, 8),
1342 => conv_std_logic_vector(1, 8),
1343 => conv_std_logic_vector(1, 8),
1344 => conv_std_logic_vector(1, 8),
1345 => conv_std_logic_vector(1, 8),
1346 => conv_std_logic_vector(1, 8),
1347 => conv_std_logic_vector(1, 8),
1348 => conv_std_logic_vector(1, 8),
1349 => conv_std_logic_vector(1, 8),
1350 => conv_std_logic_vector(1, 8),
1351 => conv_std_logic_vector(1, 8),
1352 => conv_std_logic_vector(1, 8),
1353 => conv_std_logic_vector(1, 8),
1354 => conv_std_logic_vector(1, 8),
1355 => conv_std_logic_vector(1, 8),
1356 => conv_std_logic_vector(1, 8),
1357 => conv_std_logic_vector(1, 8),
1358 => conv_std_logic_vector(1, 8),
1359 => conv_std_logic_vector(1, 8),
1360 => conv_std_logic_vector(1, 8),
1361 => conv_std_logic_vector(1, 8),
1362 => conv_std_logic_vector(1, 8),
1363 => conv_std_logic_vector(1, 8),
1364 => conv_std_logic_vector(1, 8),
1365 => conv_std_logic_vector(1, 8),
1366 => conv_std_logic_vector(1, 8),
1367 => conv_std_logic_vector(1, 8),
1368 => conv_std_logic_vector(1, 8),
1369 => conv_std_logic_vector(1, 8),
1370 => conv_std_logic_vector(1, 8),
1371 => conv_std_logic_vector(1, 8),
1372 => conv_std_logic_vector(1, 8),
1373 => conv_std_logic_vector(1, 8),
1374 => conv_std_logic_vector(1, 8),
1375 => conv_std_logic_vector(1, 8),
1376 => conv_std_logic_vector(1, 8),
1377 => conv_std_logic_vector(1, 8),
1378 => conv_std_logic_vector(1, 8),
1379 => conv_std_logic_vector(1, 8),
1380 => conv_std_logic_vector(1, 8),
1381 => conv_std_logic_vector(1, 8),
1382 => conv_std_logic_vector(1, 8),
1383 => conv_std_logic_vector(2, 8),
1384 => conv_std_logic_vector(2, 8),
1385 => conv_std_logic_vector(2, 8),
1386 => conv_std_logic_vector(2, 8),
1387 => conv_std_logic_vector(2, 8),
1388 => conv_std_logic_vector(2, 8),
1389 => conv_std_logic_vector(2, 8),
1390 => conv_std_logic_vector(2, 8),
1391 => conv_std_logic_vector(2, 8),
1392 => conv_std_logic_vector(2, 8),
1393 => conv_std_logic_vector(2, 8),
1394 => conv_std_logic_vector(2, 8),
1395 => conv_std_logic_vector(2, 8),
1396 => conv_std_logic_vector(2, 8),
1397 => conv_std_logic_vector(2, 8),
1398 => conv_std_logic_vector(2, 8),
1399 => conv_std_logic_vector(2, 8),
1400 => conv_std_logic_vector(2, 8),
1401 => conv_std_logic_vector(2, 8),
1402 => conv_std_logic_vector(2, 8),
1403 => conv_std_logic_vector(2, 8),
1404 => conv_std_logic_vector(2, 8),
1405 => conv_std_logic_vector(2, 8),
1406 => conv_std_logic_vector(2, 8),
1407 => conv_std_logic_vector(2, 8),
1408 => conv_std_logic_vector(2, 8),
1409 => conv_std_logic_vector(2, 8),
1410 => conv_std_logic_vector(2, 8),
1411 => conv_std_logic_vector(2, 8),
1412 => conv_std_logic_vector(2, 8),
1413 => conv_std_logic_vector(2, 8),
1414 => conv_std_logic_vector(2, 8),
1415 => conv_std_logic_vector(2, 8),
1416 => conv_std_logic_vector(2, 8),
1417 => conv_std_logic_vector(2, 8),
1418 => conv_std_logic_vector(2, 8),
1419 => conv_std_logic_vector(2, 8),
1420 => conv_std_logic_vector(2, 8),
1421 => conv_std_logic_vector(2, 8),
1422 => conv_std_logic_vector(2, 8),
1423 => conv_std_logic_vector(2, 8),
1424 => conv_std_logic_vector(2, 8),
1425 => conv_std_logic_vector(2, 8),
1426 => conv_std_logic_vector(2, 8),
1427 => conv_std_logic_vector(2, 8),
1428 => conv_std_logic_vector(2, 8),
1429 => conv_std_logic_vector(2, 8),
1430 => conv_std_logic_vector(2, 8),
1431 => conv_std_logic_vector(2, 8),
1432 => conv_std_logic_vector(2, 8),
1433 => conv_std_logic_vector(2, 8),
1434 => conv_std_logic_vector(3, 8),
1435 => conv_std_logic_vector(3, 8),
1436 => conv_std_logic_vector(3, 8),
1437 => conv_std_logic_vector(3, 8),
1438 => conv_std_logic_vector(3, 8),
1439 => conv_std_logic_vector(3, 8),
1440 => conv_std_logic_vector(3, 8),
1441 => conv_std_logic_vector(3, 8),
1442 => conv_std_logic_vector(3, 8),
1443 => conv_std_logic_vector(3, 8),
1444 => conv_std_logic_vector(3, 8),
1445 => conv_std_logic_vector(3, 8),
1446 => conv_std_logic_vector(3, 8),
1447 => conv_std_logic_vector(3, 8),
1448 => conv_std_logic_vector(3, 8),
1449 => conv_std_logic_vector(3, 8),
1450 => conv_std_logic_vector(3, 8),
1451 => conv_std_logic_vector(3, 8),
1452 => conv_std_logic_vector(3, 8),
1453 => conv_std_logic_vector(3, 8),
1454 => conv_std_logic_vector(3, 8),
1455 => conv_std_logic_vector(3, 8),
1456 => conv_std_logic_vector(3, 8),
1457 => conv_std_logic_vector(3, 8),
1458 => conv_std_logic_vector(3, 8),
1459 => conv_std_logic_vector(3, 8),
1460 => conv_std_logic_vector(3, 8),
1461 => conv_std_logic_vector(3, 8),
1462 => conv_std_logic_vector(3, 8),
1463 => conv_std_logic_vector(3, 8),
1464 => conv_std_logic_vector(3, 8),
1465 => conv_std_logic_vector(3, 8),
1466 => conv_std_logic_vector(3, 8),
1467 => conv_std_logic_vector(3, 8),
1468 => conv_std_logic_vector(3, 8),
1469 => conv_std_logic_vector(3, 8),
1470 => conv_std_logic_vector(3, 8),
1471 => conv_std_logic_vector(3, 8),
1472 => conv_std_logic_vector(3, 8),
1473 => conv_std_logic_vector(3, 8),
1474 => conv_std_logic_vector(3, 8),
1475 => conv_std_logic_vector(3, 8),
1476 => conv_std_logic_vector(3, 8),
1477 => conv_std_logic_vector(3, 8),
1478 => conv_std_logic_vector(3, 8),
1479 => conv_std_logic_vector(3, 8),
1480 => conv_std_logic_vector(3, 8),
1481 => conv_std_logic_vector(3, 8),
1482 => conv_std_logic_vector(3, 8),
1483 => conv_std_logic_vector(3, 8),
1484 => conv_std_logic_vector(3, 8),
1485 => conv_std_logic_vector(4, 8),
1486 => conv_std_logic_vector(4, 8),
1487 => conv_std_logic_vector(4, 8),
1488 => conv_std_logic_vector(4, 8),
1489 => conv_std_logic_vector(4, 8),
1490 => conv_std_logic_vector(4, 8),
1491 => conv_std_logic_vector(4, 8),
1492 => conv_std_logic_vector(4, 8),
1493 => conv_std_logic_vector(4, 8),
1494 => conv_std_logic_vector(4, 8),
1495 => conv_std_logic_vector(4, 8),
1496 => conv_std_logic_vector(4, 8),
1497 => conv_std_logic_vector(4, 8),
1498 => conv_std_logic_vector(4, 8),
1499 => conv_std_logic_vector(4, 8),
1500 => conv_std_logic_vector(4, 8),
1501 => conv_std_logic_vector(4, 8),
1502 => conv_std_logic_vector(4, 8),
1503 => conv_std_logic_vector(4, 8),
1504 => conv_std_logic_vector(4, 8),
1505 => conv_std_logic_vector(4, 8),
1506 => conv_std_logic_vector(4, 8),
1507 => conv_std_logic_vector(4, 8),
1508 => conv_std_logic_vector(4, 8),
1509 => conv_std_logic_vector(4, 8),
1510 => conv_std_logic_vector(4, 8),
1511 => conv_std_logic_vector(4, 8),
1512 => conv_std_logic_vector(4, 8),
1513 => conv_std_logic_vector(4, 8),
1514 => conv_std_logic_vector(4, 8),
1515 => conv_std_logic_vector(4, 8),
1516 => conv_std_logic_vector(4, 8),
1517 => conv_std_logic_vector(4, 8),
1518 => conv_std_logic_vector(4, 8),
1519 => conv_std_logic_vector(4, 8),
1520 => conv_std_logic_vector(4, 8),
1521 => conv_std_logic_vector(4, 8),
1522 => conv_std_logic_vector(4, 8),
1523 => conv_std_logic_vector(4, 8),
1524 => conv_std_logic_vector(4, 8),
1525 => conv_std_logic_vector(4, 8),
1526 => conv_std_logic_vector(4, 8),
1527 => conv_std_logic_vector(4, 8),
1528 => conv_std_logic_vector(4, 8),
1529 => conv_std_logic_vector(4, 8),
1530 => conv_std_logic_vector(4, 8),
1531 => conv_std_logic_vector(4, 8),
1532 => conv_std_logic_vector(4, 8),
1533 => conv_std_logic_vector(4, 8),
1534 => conv_std_logic_vector(4, 8),
1535 => conv_std_logic_vector(4, 8),
1536 => conv_std_logic_vector(0, 8),
1537 => conv_std_logic_vector(0, 8),
1538 => conv_std_logic_vector(0, 8),
1539 => conv_std_logic_vector(0, 8),
1540 => conv_std_logic_vector(0, 8),
1541 => conv_std_logic_vector(0, 8),
1542 => conv_std_logic_vector(0, 8),
1543 => conv_std_logic_vector(0, 8),
1544 => conv_std_logic_vector(0, 8),
1545 => conv_std_logic_vector(0, 8),
1546 => conv_std_logic_vector(0, 8),
1547 => conv_std_logic_vector(0, 8),
1548 => conv_std_logic_vector(0, 8),
1549 => conv_std_logic_vector(0, 8),
1550 => conv_std_logic_vector(0, 8),
1551 => conv_std_logic_vector(0, 8),
1552 => conv_std_logic_vector(0, 8),
1553 => conv_std_logic_vector(0, 8),
1554 => conv_std_logic_vector(0, 8),
1555 => conv_std_logic_vector(0, 8),
1556 => conv_std_logic_vector(0, 8),
1557 => conv_std_logic_vector(0, 8),
1558 => conv_std_logic_vector(0, 8),
1559 => conv_std_logic_vector(0, 8),
1560 => conv_std_logic_vector(0, 8),
1561 => conv_std_logic_vector(0, 8),
1562 => conv_std_logic_vector(0, 8),
1563 => conv_std_logic_vector(0, 8),
1564 => conv_std_logic_vector(0, 8),
1565 => conv_std_logic_vector(0, 8),
1566 => conv_std_logic_vector(0, 8),
1567 => conv_std_logic_vector(0, 8),
1568 => conv_std_logic_vector(0, 8),
1569 => conv_std_logic_vector(0, 8),
1570 => conv_std_logic_vector(0, 8),
1571 => conv_std_logic_vector(0, 8),
1572 => conv_std_logic_vector(0, 8),
1573 => conv_std_logic_vector(0, 8),
1574 => conv_std_logic_vector(0, 8),
1575 => conv_std_logic_vector(0, 8),
1576 => conv_std_logic_vector(0, 8),
1577 => conv_std_logic_vector(0, 8),
1578 => conv_std_logic_vector(0, 8),
1579 => conv_std_logic_vector(1, 8),
1580 => conv_std_logic_vector(1, 8),
1581 => conv_std_logic_vector(1, 8),
1582 => conv_std_logic_vector(1, 8),
1583 => conv_std_logic_vector(1, 8),
1584 => conv_std_logic_vector(1, 8),
1585 => conv_std_logic_vector(1, 8),
1586 => conv_std_logic_vector(1, 8),
1587 => conv_std_logic_vector(1, 8),
1588 => conv_std_logic_vector(1, 8),
1589 => conv_std_logic_vector(1, 8),
1590 => conv_std_logic_vector(1, 8),
1591 => conv_std_logic_vector(1, 8),
1592 => conv_std_logic_vector(1, 8),
1593 => conv_std_logic_vector(1, 8),
1594 => conv_std_logic_vector(1, 8),
1595 => conv_std_logic_vector(1, 8),
1596 => conv_std_logic_vector(1, 8),
1597 => conv_std_logic_vector(1, 8),
1598 => conv_std_logic_vector(1, 8),
1599 => conv_std_logic_vector(1, 8),
1600 => conv_std_logic_vector(1, 8),
1601 => conv_std_logic_vector(1, 8),
1602 => conv_std_logic_vector(1, 8),
1603 => conv_std_logic_vector(1, 8),
1604 => conv_std_logic_vector(1, 8),
1605 => conv_std_logic_vector(1, 8),
1606 => conv_std_logic_vector(1, 8),
1607 => conv_std_logic_vector(1, 8),
1608 => conv_std_logic_vector(1, 8),
1609 => conv_std_logic_vector(1, 8),
1610 => conv_std_logic_vector(1, 8),
1611 => conv_std_logic_vector(1, 8),
1612 => conv_std_logic_vector(1, 8),
1613 => conv_std_logic_vector(1, 8),
1614 => conv_std_logic_vector(1, 8),
1615 => conv_std_logic_vector(1, 8),
1616 => conv_std_logic_vector(1, 8),
1617 => conv_std_logic_vector(1, 8),
1618 => conv_std_logic_vector(1, 8),
1619 => conv_std_logic_vector(1, 8),
1620 => conv_std_logic_vector(1, 8),
1621 => conv_std_logic_vector(1, 8),
1622 => conv_std_logic_vector(2, 8),
1623 => conv_std_logic_vector(2, 8),
1624 => conv_std_logic_vector(2, 8),
1625 => conv_std_logic_vector(2, 8),
1626 => conv_std_logic_vector(2, 8),
1627 => conv_std_logic_vector(2, 8),
1628 => conv_std_logic_vector(2, 8),
1629 => conv_std_logic_vector(2, 8),
1630 => conv_std_logic_vector(2, 8),
1631 => conv_std_logic_vector(2, 8),
1632 => conv_std_logic_vector(2, 8),
1633 => conv_std_logic_vector(2, 8),
1634 => conv_std_logic_vector(2, 8),
1635 => conv_std_logic_vector(2, 8),
1636 => conv_std_logic_vector(2, 8),
1637 => conv_std_logic_vector(2, 8),
1638 => conv_std_logic_vector(2, 8),
1639 => conv_std_logic_vector(2, 8),
1640 => conv_std_logic_vector(2, 8),
1641 => conv_std_logic_vector(2, 8),
1642 => conv_std_logic_vector(2, 8),
1643 => conv_std_logic_vector(2, 8),
1644 => conv_std_logic_vector(2, 8),
1645 => conv_std_logic_vector(2, 8),
1646 => conv_std_logic_vector(2, 8),
1647 => conv_std_logic_vector(2, 8),
1648 => conv_std_logic_vector(2, 8),
1649 => conv_std_logic_vector(2, 8),
1650 => conv_std_logic_vector(2, 8),
1651 => conv_std_logic_vector(2, 8),
1652 => conv_std_logic_vector(2, 8),
1653 => conv_std_logic_vector(2, 8),
1654 => conv_std_logic_vector(2, 8),
1655 => conv_std_logic_vector(2, 8),
1656 => conv_std_logic_vector(2, 8),
1657 => conv_std_logic_vector(2, 8),
1658 => conv_std_logic_vector(2, 8),
1659 => conv_std_logic_vector(2, 8),
1660 => conv_std_logic_vector(2, 8),
1661 => conv_std_logic_vector(2, 8),
1662 => conv_std_logic_vector(2, 8),
1663 => conv_std_logic_vector(2, 8),
1664 => conv_std_logic_vector(3, 8),
1665 => conv_std_logic_vector(3, 8),
1666 => conv_std_logic_vector(3, 8),
1667 => conv_std_logic_vector(3, 8),
1668 => conv_std_logic_vector(3, 8),
1669 => conv_std_logic_vector(3, 8),
1670 => conv_std_logic_vector(3, 8),
1671 => conv_std_logic_vector(3, 8),
1672 => conv_std_logic_vector(3, 8),
1673 => conv_std_logic_vector(3, 8),
1674 => conv_std_logic_vector(3, 8),
1675 => conv_std_logic_vector(3, 8),
1676 => conv_std_logic_vector(3, 8),
1677 => conv_std_logic_vector(3, 8),
1678 => conv_std_logic_vector(3, 8),
1679 => conv_std_logic_vector(3, 8),
1680 => conv_std_logic_vector(3, 8),
1681 => conv_std_logic_vector(3, 8),
1682 => conv_std_logic_vector(3, 8),
1683 => conv_std_logic_vector(3, 8),
1684 => conv_std_logic_vector(3, 8),
1685 => conv_std_logic_vector(3, 8),
1686 => conv_std_logic_vector(3, 8),
1687 => conv_std_logic_vector(3, 8),
1688 => conv_std_logic_vector(3, 8),
1689 => conv_std_logic_vector(3, 8),
1690 => conv_std_logic_vector(3, 8),
1691 => conv_std_logic_vector(3, 8),
1692 => conv_std_logic_vector(3, 8),
1693 => conv_std_logic_vector(3, 8),
1694 => conv_std_logic_vector(3, 8),
1695 => conv_std_logic_vector(3, 8),
1696 => conv_std_logic_vector(3, 8),
1697 => conv_std_logic_vector(3, 8),
1698 => conv_std_logic_vector(3, 8),
1699 => conv_std_logic_vector(3, 8),
1700 => conv_std_logic_vector(3, 8),
1701 => conv_std_logic_vector(3, 8),
1702 => conv_std_logic_vector(3, 8),
1703 => conv_std_logic_vector(3, 8),
1704 => conv_std_logic_vector(3, 8),
1705 => conv_std_logic_vector(3, 8),
1706 => conv_std_logic_vector(3, 8),
1707 => conv_std_logic_vector(4, 8),
1708 => conv_std_logic_vector(4, 8),
1709 => conv_std_logic_vector(4, 8),
1710 => conv_std_logic_vector(4, 8),
1711 => conv_std_logic_vector(4, 8),
1712 => conv_std_logic_vector(4, 8),
1713 => conv_std_logic_vector(4, 8),
1714 => conv_std_logic_vector(4, 8),
1715 => conv_std_logic_vector(4, 8),
1716 => conv_std_logic_vector(4, 8),
1717 => conv_std_logic_vector(4, 8),
1718 => conv_std_logic_vector(4, 8),
1719 => conv_std_logic_vector(4, 8),
1720 => conv_std_logic_vector(4, 8),
1721 => conv_std_logic_vector(4, 8),
1722 => conv_std_logic_vector(4, 8),
1723 => conv_std_logic_vector(4, 8),
1724 => conv_std_logic_vector(4, 8),
1725 => conv_std_logic_vector(4, 8),
1726 => conv_std_logic_vector(4, 8),
1727 => conv_std_logic_vector(4, 8),
1728 => conv_std_logic_vector(4, 8),
1729 => conv_std_logic_vector(4, 8),
1730 => conv_std_logic_vector(4, 8),
1731 => conv_std_logic_vector(4, 8),
1732 => conv_std_logic_vector(4, 8),
1733 => conv_std_logic_vector(4, 8),
1734 => conv_std_logic_vector(4, 8),
1735 => conv_std_logic_vector(4, 8),
1736 => conv_std_logic_vector(4, 8),
1737 => conv_std_logic_vector(4, 8),
1738 => conv_std_logic_vector(4, 8),
1739 => conv_std_logic_vector(4, 8),
1740 => conv_std_logic_vector(4, 8),
1741 => conv_std_logic_vector(4, 8),
1742 => conv_std_logic_vector(4, 8),
1743 => conv_std_logic_vector(4, 8),
1744 => conv_std_logic_vector(4, 8),
1745 => conv_std_logic_vector(4, 8),
1746 => conv_std_logic_vector(4, 8),
1747 => conv_std_logic_vector(4, 8),
1748 => conv_std_logic_vector(4, 8),
1749 => conv_std_logic_vector(4, 8),
1750 => conv_std_logic_vector(5, 8),
1751 => conv_std_logic_vector(5, 8),
1752 => conv_std_logic_vector(5, 8),
1753 => conv_std_logic_vector(5, 8),
1754 => conv_std_logic_vector(5, 8),
1755 => conv_std_logic_vector(5, 8),
1756 => conv_std_logic_vector(5, 8),
1757 => conv_std_logic_vector(5, 8),
1758 => conv_std_logic_vector(5, 8),
1759 => conv_std_logic_vector(5, 8),
1760 => conv_std_logic_vector(5, 8),
1761 => conv_std_logic_vector(5, 8),
1762 => conv_std_logic_vector(5, 8),
1763 => conv_std_logic_vector(5, 8),
1764 => conv_std_logic_vector(5, 8),
1765 => conv_std_logic_vector(5, 8),
1766 => conv_std_logic_vector(5, 8),
1767 => conv_std_logic_vector(5, 8),
1768 => conv_std_logic_vector(5, 8),
1769 => conv_std_logic_vector(5, 8),
1770 => conv_std_logic_vector(5, 8),
1771 => conv_std_logic_vector(5, 8),
1772 => conv_std_logic_vector(5, 8),
1773 => conv_std_logic_vector(5, 8),
1774 => conv_std_logic_vector(5, 8),
1775 => conv_std_logic_vector(5, 8),
1776 => conv_std_logic_vector(5, 8),
1777 => conv_std_logic_vector(5, 8),
1778 => conv_std_logic_vector(5, 8),
1779 => conv_std_logic_vector(5, 8),
1780 => conv_std_logic_vector(5, 8),
1781 => conv_std_logic_vector(5, 8),
1782 => conv_std_logic_vector(5, 8),
1783 => conv_std_logic_vector(5, 8),
1784 => conv_std_logic_vector(5, 8),
1785 => conv_std_logic_vector(5, 8),
1786 => conv_std_logic_vector(5, 8),
1787 => conv_std_logic_vector(5, 8),
1788 => conv_std_logic_vector(5, 8),
1789 => conv_std_logic_vector(5, 8),
1790 => conv_std_logic_vector(5, 8),
1791 => conv_std_logic_vector(5, 8),
1792 => conv_std_logic_vector(0, 8),
1793 => conv_std_logic_vector(0, 8),
1794 => conv_std_logic_vector(0, 8),
1795 => conv_std_logic_vector(0, 8),
1796 => conv_std_logic_vector(0, 8),
1797 => conv_std_logic_vector(0, 8),
1798 => conv_std_logic_vector(0, 8),
1799 => conv_std_logic_vector(0, 8),
1800 => conv_std_logic_vector(0, 8),
1801 => conv_std_logic_vector(0, 8),
1802 => conv_std_logic_vector(0, 8),
1803 => conv_std_logic_vector(0, 8),
1804 => conv_std_logic_vector(0, 8),
1805 => conv_std_logic_vector(0, 8),
1806 => conv_std_logic_vector(0, 8),
1807 => conv_std_logic_vector(0, 8),
1808 => conv_std_logic_vector(0, 8),
1809 => conv_std_logic_vector(0, 8),
1810 => conv_std_logic_vector(0, 8),
1811 => conv_std_logic_vector(0, 8),
1812 => conv_std_logic_vector(0, 8),
1813 => conv_std_logic_vector(0, 8),
1814 => conv_std_logic_vector(0, 8),
1815 => conv_std_logic_vector(0, 8),
1816 => conv_std_logic_vector(0, 8),
1817 => conv_std_logic_vector(0, 8),
1818 => conv_std_logic_vector(0, 8),
1819 => conv_std_logic_vector(0, 8),
1820 => conv_std_logic_vector(0, 8),
1821 => conv_std_logic_vector(0, 8),
1822 => conv_std_logic_vector(0, 8),
1823 => conv_std_logic_vector(0, 8),
1824 => conv_std_logic_vector(0, 8),
1825 => conv_std_logic_vector(0, 8),
1826 => conv_std_logic_vector(0, 8),
1827 => conv_std_logic_vector(0, 8),
1828 => conv_std_logic_vector(0, 8),
1829 => conv_std_logic_vector(1, 8),
1830 => conv_std_logic_vector(1, 8),
1831 => conv_std_logic_vector(1, 8),
1832 => conv_std_logic_vector(1, 8),
1833 => conv_std_logic_vector(1, 8),
1834 => conv_std_logic_vector(1, 8),
1835 => conv_std_logic_vector(1, 8),
1836 => conv_std_logic_vector(1, 8),
1837 => conv_std_logic_vector(1, 8),
1838 => conv_std_logic_vector(1, 8),
1839 => conv_std_logic_vector(1, 8),
1840 => conv_std_logic_vector(1, 8),
1841 => conv_std_logic_vector(1, 8),
1842 => conv_std_logic_vector(1, 8),
1843 => conv_std_logic_vector(1, 8),
1844 => conv_std_logic_vector(1, 8),
1845 => conv_std_logic_vector(1, 8),
1846 => conv_std_logic_vector(1, 8),
1847 => conv_std_logic_vector(1, 8),
1848 => conv_std_logic_vector(1, 8),
1849 => conv_std_logic_vector(1, 8),
1850 => conv_std_logic_vector(1, 8),
1851 => conv_std_logic_vector(1, 8),
1852 => conv_std_logic_vector(1, 8),
1853 => conv_std_logic_vector(1, 8),
1854 => conv_std_logic_vector(1, 8),
1855 => conv_std_logic_vector(1, 8),
1856 => conv_std_logic_vector(1, 8),
1857 => conv_std_logic_vector(1, 8),
1858 => conv_std_logic_vector(1, 8),
1859 => conv_std_logic_vector(1, 8),
1860 => conv_std_logic_vector(1, 8),
1861 => conv_std_logic_vector(1, 8),
1862 => conv_std_logic_vector(1, 8),
1863 => conv_std_logic_vector(1, 8),
1864 => conv_std_logic_vector(1, 8),
1865 => conv_std_logic_vector(1, 8),
1866 => conv_std_logic_vector(2, 8),
1867 => conv_std_logic_vector(2, 8),
1868 => conv_std_logic_vector(2, 8),
1869 => conv_std_logic_vector(2, 8),
1870 => conv_std_logic_vector(2, 8),
1871 => conv_std_logic_vector(2, 8),
1872 => conv_std_logic_vector(2, 8),
1873 => conv_std_logic_vector(2, 8),
1874 => conv_std_logic_vector(2, 8),
1875 => conv_std_logic_vector(2, 8),
1876 => conv_std_logic_vector(2, 8),
1877 => conv_std_logic_vector(2, 8),
1878 => conv_std_logic_vector(2, 8),
1879 => conv_std_logic_vector(2, 8),
1880 => conv_std_logic_vector(2, 8),
1881 => conv_std_logic_vector(2, 8),
1882 => conv_std_logic_vector(2, 8),
1883 => conv_std_logic_vector(2, 8),
1884 => conv_std_logic_vector(2, 8),
1885 => conv_std_logic_vector(2, 8),
1886 => conv_std_logic_vector(2, 8),
1887 => conv_std_logic_vector(2, 8),
1888 => conv_std_logic_vector(2, 8),
1889 => conv_std_logic_vector(2, 8),
1890 => conv_std_logic_vector(2, 8),
1891 => conv_std_logic_vector(2, 8),
1892 => conv_std_logic_vector(2, 8),
1893 => conv_std_logic_vector(2, 8),
1894 => conv_std_logic_vector(2, 8),
1895 => conv_std_logic_vector(2, 8),
1896 => conv_std_logic_vector(2, 8),
1897 => conv_std_logic_vector(2, 8),
1898 => conv_std_logic_vector(2, 8),
1899 => conv_std_logic_vector(2, 8),
1900 => conv_std_logic_vector(2, 8),
1901 => conv_std_logic_vector(2, 8),
1902 => conv_std_logic_vector(3, 8),
1903 => conv_std_logic_vector(3, 8),
1904 => conv_std_logic_vector(3, 8),
1905 => conv_std_logic_vector(3, 8),
1906 => conv_std_logic_vector(3, 8),
1907 => conv_std_logic_vector(3, 8),
1908 => conv_std_logic_vector(3, 8),
1909 => conv_std_logic_vector(3, 8),
1910 => conv_std_logic_vector(3, 8),
1911 => conv_std_logic_vector(3, 8),
1912 => conv_std_logic_vector(3, 8),
1913 => conv_std_logic_vector(3, 8),
1914 => conv_std_logic_vector(3, 8),
1915 => conv_std_logic_vector(3, 8),
1916 => conv_std_logic_vector(3, 8),
1917 => conv_std_logic_vector(3, 8),
1918 => conv_std_logic_vector(3, 8),
1919 => conv_std_logic_vector(3, 8),
1920 => conv_std_logic_vector(3, 8),
1921 => conv_std_logic_vector(3, 8),
1922 => conv_std_logic_vector(3, 8),
1923 => conv_std_logic_vector(3, 8),
1924 => conv_std_logic_vector(3, 8),
1925 => conv_std_logic_vector(3, 8),
1926 => conv_std_logic_vector(3, 8),
1927 => conv_std_logic_vector(3, 8),
1928 => conv_std_logic_vector(3, 8),
1929 => conv_std_logic_vector(3, 8),
1930 => conv_std_logic_vector(3, 8),
1931 => conv_std_logic_vector(3, 8),
1932 => conv_std_logic_vector(3, 8),
1933 => conv_std_logic_vector(3, 8),
1934 => conv_std_logic_vector(3, 8),
1935 => conv_std_logic_vector(3, 8),
1936 => conv_std_logic_vector(3, 8),
1937 => conv_std_logic_vector(3, 8),
1938 => conv_std_logic_vector(3, 8),
1939 => conv_std_logic_vector(4, 8),
1940 => conv_std_logic_vector(4, 8),
1941 => conv_std_logic_vector(4, 8),
1942 => conv_std_logic_vector(4, 8),
1943 => conv_std_logic_vector(4, 8),
1944 => conv_std_logic_vector(4, 8),
1945 => conv_std_logic_vector(4, 8),
1946 => conv_std_logic_vector(4, 8),
1947 => conv_std_logic_vector(4, 8),
1948 => conv_std_logic_vector(4, 8),
1949 => conv_std_logic_vector(4, 8),
1950 => conv_std_logic_vector(4, 8),
1951 => conv_std_logic_vector(4, 8),
1952 => conv_std_logic_vector(4, 8),
1953 => conv_std_logic_vector(4, 8),
1954 => conv_std_logic_vector(4, 8),
1955 => conv_std_logic_vector(4, 8),
1956 => conv_std_logic_vector(4, 8),
1957 => conv_std_logic_vector(4, 8),
1958 => conv_std_logic_vector(4, 8),
1959 => conv_std_logic_vector(4, 8),
1960 => conv_std_logic_vector(4, 8),
1961 => conv_std_logic_vector(4, 8),
1962 => conv_std_logic_vector(4, 8),
1963 => conv_std_logic_vector(4, 8),
1964 => conv_std_logic_vector(4, 8),
1965 => conv_std_logic_vector(4, 8),
1966 => conv_std_logic_vector(4, 8),
1967 => conv_std_logic_vector(4, 8),
1968 => conv_std_logic_vector(4, 8),
1969 => conv_std_logic_vector(4, 8),
1970 => conv_std_logic_vector(4, 8),
1971 => conv_std_logic_vector(4, 8),
1972 => conv_std_logic_vector(4, 8),
1973 => conv_std_logic_vector(4, 8),
1974 => conv_std_logic_vector(4, 8),
1975 => conv_std_logic_vector(5, 8),
1976 => conv_std_logic_vector(5, 8),
1977 => conv_std_logic_vector(5, 8),
1978 => conv_std_logic_vector(5, 8),
1979 => conv_std_logic_vector(5, 8),
1980 => conv_std_logic_vector(5, 8),
1981 => conv_std_logic_vector(5, 8),
1982 => conv_std_logic_vector(5, 8),
1983 => conv_std_logic_vector(5, 8),
1984 => conv_std_logic_vector(5, 8),
1985 => conv_std_logic_vector(5, 8),
1986 => conv_std_logic_vector(5, 8),
1987 => conv_std_logic_vector(5, 8),
1988 => conv_std_logic_vector(5, 8),
1989 => conv_std_logic_vector(5, 8),
1990 => conv_std_logic_vector(5, 8),
1991 => conv_std_logic_vector(5, 8),
1992 => conv_std_logic_vector(5, 8),
1993 => conv_std_logic_vector(5, 8),
1994 => conv_std_logic_vector(5, 8),
1995 => conv_std_logic_vector(5, 8),
1996 => conv_std_logic_vector(5, 8),
1997 => conv_std_logic_vector(5, 8),
1998 => conv_std_logic_vector(5, 8),
1999 => conv_std_logic_vector(5, 8),
2000 => conv_std_logic_vector(5, 8),
2001 => conv_std_logic_vector(5, 8),
2002 => conv_std_logic_vector(5, 8),
2003 => conv_std_logic_vector(5, 8),
2004 => conv_std_logic_vector(5, 8),
2005 => conv_std_logic_vector(5, 8),
2006 => conv_std_logic_vector(5, 8),
2007 => conv_std_logic_vector(5, 8),
2008 => conv_std_logic_vector(5, 8),
2009 => conv_std_logic_vector(5, 8),
2010 => conv_std_logic_vector(5, 8),
2011 => conv_std_logic_vector(5, 8),
2012 => conv_std_logic_vector(6, 8),
2013 => conv_std_logic_vector(6, 8),
2014 => conv_std_logic_vector(6, 8),
2015 => conv_std_logic_vector(6, 8),
2016 => conv_std_logic_vector(6, 8),
2017 => conv_std_logic_vector(6, 8),
2018 => conv_std_logic_vector(6, 8),
2019 => conv_std_logic_vector(6, 8),
2020 => conv_std_logic_vector(6, 8),
2021 => conv_std_logic_vector(6, 8),
2022 => conv_std_logic_vector(6, 8),
2023 => conv_std_logic_vector(6, 8),
2024 => conv_std_logic_vector(6, 8),
2025 => conv_std_logic_vector(6, 8),
2026 => conv_std_logic_vector(6, 8),
2027 => conv_std_logic_vector(6, 8),
2028 => conv_std_logic_vector(6, 8),
2029 => conv_std_logic_vector(6, 8),
2030 => conv_std_logic_vector(6, 8),
2031 => conv_std_logic_vector(6, 8),
2032 => conv_std_logic_vector(6, 8),
2033 => conv_std_logic_vector(6, 8),
2034 => conv_std_logic_vector(6, 8),
2035 => conv_std_logic_vector(6, 8),
2036 => conv_std_logic_vector(6, 8),
2037 => conv_std_logic_vector(6, 8),
2038 => conv_std_logic_vector(6, 8),
2039 => conv_std_logic_vector(6, 8),
2040 => conv_std_logic_vector(6, 8),
2041 => conv_std_logic_vector(6, 8),
2042 => conv_std_logic_vector(6, 8),
2043 => conv_std_logic_vector(6, 8),
2044 => conv_std_logic_vector(6, 8),
2045 => conv_std_logic_vector(6, 8),
2046 => conv_std_logic_vector(6, 8),
2047 => conv_std_logic_vector(6, 8),
2048 => conv_std_logic_vector(0, 8),
2049 => conv_std_logic_vector(0, 8),
2050 => conv_std_logic_vector(0, 8),
2051 => conv_std_logic_vector(0, 8),
2052 => conv_std_logic_vector(0, 8),
2053 => conv_std_logic_vector(0, 8),
2054 => conv_std_logic_vector(0, 8),
2055 => conv_std_logic_vector(0, 8),
2056 => conv_std_logic_vector(0, 8),
2057 => conv_std_logic_vector(0, 8),
2058 => conv_std_logic_vector(0, 8),
2059 => conv_std_logic_vector(0, 8),
2060 => conv_std_logic_vector(0, 8),
2061 => conv_std_logic_vector(0, 8),
2062 => conv_std_logic_vector(0, 8),
2063 => conv_std_logic_vector(0, 8),
2064 => conv_std_logic_vector(0, 8),
2065 => conv_std_logic_vector(0, 8),
2066 => conv_std_logic_vector(0, 8),
2067 => conv_std_logic_vector(0, 8),
2068 => conv_std_logic_vector(0, 8),
2069 => conv_std_logic_vector(0, 8),
2070 => conv_std_logic_vector(0, 8),
2071 => conv_std_logic_vector(0, 8),
2072 => conv_std_logic_vector(0, 8),
2073 => conv_std_logic_vector(0, 8),
2074 => conv_std_logic_vector(0, 8),
2075 => conv_std_logic_vector(0, 8),
2076 => conv_std_logic_vector(0, 8),
2077 => conv_std_logic_vector(0, 8),
2078 => conv_std_logic_vector(0, 8),
2079 => conv_std_logic_vector(0, 8),
2080 => conv_std_logic_vector(1, 8),
2081 => conv_std_logic_vector(1, 8),
2082 => conv_std_logic_vector(1, 8),
2083 => conv_std_logic_vector(1, 8),
2084 => conv_std_logic_vector(1, 8),
2085 => conv_std_logic_vector(1, 8),
2086 => conv_std_logic_vector(1, 8),
2087 => conv_std_logic_vector(1, 8),
2088 => conv_std_logic_vector(1, 8),
2089 => conv_std_logic_vector(1, 8),
2090 => conv_std_logic_vector(1, 8),
2091 => conv_std_logic_vector(1, 8),
2092 => conv_std_logic_vector(1, 8),
2093 => conv_std_logic_vector(1, 8),
2094 => conv_std_logic_vector(1, 8),
2095 => conv_std_logic_vector(1, 8),
2096 => conv_std_logic_vector(1, 8),
2097 => conv_std_logic_vector(1, 8),
2098 => conv_std_logic_vector(1, 8),
2099 => conv_std_logic_vector(1, 8),
2100 => conv_std_logic_vector(1, 8),
2101 => conv_std_logic_vector(1, 8),
2102 => conv_std_logic_vector(1, 8),
2103 => conv_std_logic_vector(1, 8),
2104 => conv_std_logic_vector(1, 8),
2105 => conv_std_logic_vector(1, 8),
2106 => conv_std_logic_vector(1, 8),
2107 => conv_std_logic_vector(1, 8),
2108 => conv_std_logic_vector(1, 8),
2109 => conv_std_logic_vector(1, 8),
2110 => conv_std_logic_vector(1, 8),
2111 => conv_std_logic_vector(1, 8),
2112 => conv_std_logic_vector(2, 8),
2113 => conv_std_logic_vector(2, 8),
2114 => conv_std_logic_vector(2, 8),
2115 => conv_std_logic_vector(2, 8),
2116 => conv_std_logic_vector(2, 8),
2117 => conv_std_logic_vector(2, 8),
2118 => conv_std_logic_vector(2, 8),
2119 => conv_std_logic_vector(2, 8),
2120 => conv_std_logic_vector(2, 8),
2121 => conv_std_logic_vector(2, 8),
2122 => conv_std_logic_vector(2, 8),
2123 => conv_std_logic_vector(2, 8),
2124 => conv_std_logic_vector(2, 8),
2125 => conv_std_logic_vector(2, 8),
2126 => conv_std_logic_vector(2, 8),
2127 => conv_std_logic_vector(2, 8),
2128 => conv_std_logic_vector(2, 8),
2129 => conv_std_logic_vector(2, 8),
2130 => conv_std_logic_vector(2, 8),
2131 => conv_std_logic_vector(2, 8),
2132 => conv_std_logic_vector(2, 8),
2133 => conv_std_logic_vector(2, 8),
2134 => conv_std_logic_vector(2, 8),
2135 => conv_std_logic_vector(2, 8),
2136 => conv_std_logic_vector(2, 8),
2137 => conv_std_logic_vector(2, 8),
2138 => conv_std_logic_vector(2, 8),
2139 => conv_std_logic_vector(2, 8),
2140 => conv_std_logic_vector(2, 8),
2141 => conv_std_logic_vector(2, 8),
2142 => conv_std_logic_vector(2, 8),
2143 => conv_std_logic_vector(2, 8),
2144 => conv_std_logic_vector(3, 8),
2145 => conv_std_logic_vector(3, 8),
2146 => conv_std_logic_vector(3, 8),
2147 => conv_std_logic_vector(3, 8),
2148 => conv_std_logic_vector(3, 8),
2149 => conv_std_logic_vector(3, 8),
2150 => conv_std_logic_vector(3, 8),
2151 => conv_std_logic_vector(3, 8),
2152 => conv_std_logic_vector(3, 8),
2153 => conv_std_logic_vector(3, 8),
2154 => conv_std_logic_vector(3, 8),
2155 => conv_std_logic_vector(3, 8),
2156 => conv_std_logic_vector(3, 8),
2157 => conv_std_logic_vector(3, 8),
2158 => conv_std_logic_vector(3, 8),
2159 => conv_std_logic_vector(3, 8),
2160 => conv_std_logic_vector(3, 8),
2161 => conv_std_logic_vector(3, 8),
2162 => conv_std_logic_vector(3, 8),
2163 => conv_std_logic_vector(3, 8),
2164 => conv_std_logic_vector(3, 8),
2165 => conv_std_logic_vector(3, 8),
2166 => conv_std_logic_vector(3, 8),
2167 => conv_std_logic_vector(3, 8),
2168 => conv_std_logic_vector(3, 8),
2169 => conv_std_logic_vector(3, 8),
2170 => conv_std_logic_vector(3, 8),
2171 => conv_std_logic_vector(3, 8),
2172 => conv_std_logic_vector(3, 8),
2173 => conv_std_logic_vector(3, 8),
2174 => conv_std_logic_vector(3, 8),
2175 => conv_std_logic_vector(3, 8),
2176 => conv_std_logic_vector(4, 8),
2177 => conv_std_logic_vector(4, 8),
2178 => conv_std_logic_vector(4, 8),
2179 => conv_std_logic_vector(4, 8),
2180 => conv_std_logic_vector(4, 8),
2181 => conv_std_logic_vector(4, 8),
2182 => conv_std_logic_vector(4, 8),
2183 => conv_std_logic_vector(4, 8),
2184 => conv_std_logic_vector(4, 8),
2185 => conv_std_logic_vector(4, 8),
2186 => conv_std_logic_vector(4, 8),
2187 => conv_std_logic_vector(4, 8),
2188 => conv_std_logic_vector(4, 8),
2189 => conv_std_logic_vector(4, 8),
2190 => conv_std_logic_vector(4, 8),
2191 => conv_std_logic_vector(4, 8),
2192 => conv_std_logic_vector(4, 8),
2193 => conv_std_logic_vector(4, 8),
2194 => conv_std_logic_vector(4, 8),
2195 => conv_std_logic_vector(4, 8),
2196 => conv_std_logic_vector(4, 8),
2197 => conv_std_logic_vector(4, 8),
2198 => conv_std_logic_vector(4, 8),
2199 => conv_std_logic_vector(4, 8),
2200 => conv_std_logic_vector(4, 8),
2201 => conv_std_logic_vector(4, 8),
2202 => conv_std_logic_vector(4, 8),
2203 => conv_std_logic_vector(4, 8),
2204 => conv_std_logic_vector(4, 8),
2205 => conv_std_logic_vector(4, 8),
2206 => conv_std_logic_vector(4, 8),
2207 => conv_std_logic_vector(4, 8),
2208 => conv_std_logic_vector(5, 8),
2209 => conv_std_logic_vector(5, 8),
2210 => conv_std_logic_vector(5, 8),
2211 => conv_std_logic_vector(5, 8),
2212 => conv_std_logic_vector(5, 8),
2213 => conv_std_logic_vector(5, 8),
2214 => conv_std_logic_vector(5, 8),
2215 => conv_std_logic_vector(5, 8),
2216 => conv_std_logic_vector(5, 8),
2217 => conv_std_logic_vector(5, 8),
2218 => conv_std_logic_vector(5, 8),
2219 => conv_std_logic_vector(5, 8),
2220 => conv_std_logic_vector(5, 8),
2221 => conv_std_logic_vector(5, 8),
2222 => conv_std_logic_vector(5, 8),
2223 => conv_std_logic_vector(5, 8),
2224 => conv_std_logic_vector(5, 8),
2225 => conv_std_logic_vector(5, 8),
2226 => conv_std_logic_vector(5, 8),
2227 => conv_std_logic_vector(5, 8),
2228 => conv_std_logic_vector(5, 8),
2229 => conv_std_logic_vector(5, 8),
2230 => conv_std_logic_vector(5, 8),
2231 => conv_std_logic_vector(5, 8),
2232 => conv_std_logic_vector(5, 8),
2233 => conv_std_logic_vector(5, 8),
2234 => conv_std_logic_vector(5, 8),
2235 => conv_std_logic_vector(5, 8),
2236 => conv_std_logic_vector(5, 8),
2237 => conv_std_logic_vector(5, 8),
2238 => conv_std_logic_vector(5, 8),
2239 => conv_std_logic_vector(5, 8),
2240 => conv_std_logic_vector(6, 8),
2241 => conv_std_logic_vector(6, 8),
2242 => conv_std_logic_vector(6, 8),
2243 => conv_std_logic_vector(6, 8),
2244 => conv_std_logic_vector(6, 8),
2245 => conv_std_logic_vector(6, 8),
2246 => conv_std_logic_vector(6, 8),
2247 => conv_std_logic_vector(6, 8),
2248 => conv_std_logic_vector(6, 8),
2249 => conv_std_logic_vector(6, 8),
2250 => conv_std_logic_vector(6, 8),
2251 => conv_std_logic_vector(6, 8),
2252 => conv_std_logic_vector(6, 8),
2253 => conv_std_logic_vector(6, 8),
2254 => conv_std_logic_vector(6, 8),
2255 => conv_std_logic_vector(6, 8),
2256 => conv_std_logic_vector(6, 8),
2257 => conv_std_logic_vector(6, 8),
2258 => conv_std_logic_vector(6, 8),
2259 => conv_std_logic_vector(6, 8),
2260 => conv_std_logic_vector(6, 8),
2261 => conv_std_logic_vector(6, 8),
2262 => conv_std_logic_vector(6, 8),
2263 => conv_std_logic_vector(6, 8),
2264 => conv_std_logic_vector(6, 8),
2265 => conv_std_logic_vector(6, 8),
2266 => conv_std_logic_vector(6, 8),
2267 => conv_std_logic_vector(6, 8),
2268 => conv_std_logic_vector(6, 8),
2269 => conv_std_logic_vector(6, 8),
2270 => conv_std_logic_vector(6, 8),
2271 => conv_std_logic_vector(6, 8),
2272 => conv_std_logic_vector(7, 8),
2273 => conv_std_logic_vector(7, 8),
2274 => conv_std_logic_vector(7, 8),
2275 => conv_std_logic_vector(7, 8),
2276 => conv_std_logic_vector(7, 8),
2277 => conv_std_logic_vector(7, 8),
2278 => conv_std_logic_vector(7, 8),
2279 => conv_std_logic_vector(7, 8),
2280 => conv_std_logic_vector(7, 8),
2281 => conv_std_logic_vector(7, 8),
2282 => conv_std_logic_vector(7, 8),
2283 => conv_std_logic_vector(7, 8),
2284 => conv_std_logic_vector(7, 8),
2285 => conv_std_logic_vector(7, 8),
2286 => conv_std_logic_vector(7, 8),
2287 => conv_std_logic_vector(7, 8),
2288 => conv_std_logic_vector(7, 8),
2289 => conv_std_logic_vector(7, 8),
2290 => conv_std_logic_vector(7, 8),
2291 => conv_std_logic_vector(7, 8),
2292 => conv_std_logic_vector(7, 8),
2293 => conv_std_logic_vector(7, 8),
2294 => conv_std_logic_vector(7, 8),
2295 => conv_std_logic_vector(7, 8),
2296 => conv_std_logic_vector(7, 8),
2297 => conv_std_logic_vector(7, 8),
2298 => conv_std_logic_vector(7, 8),
2299 => conv_std_logic_vector(7, 8),
2300 => conv_std_logic_vector(7, 8),
2301 => conv_std_logic_vector(7, 8),
2302 => conv_std_logic_vector(7, 8),
2303 => conv_std_logic_vector(7, 8),
2304 => conv_std_logic_vector(0, 8),
2305 => conv_std_logic_vector(0, 8),
2306 => conv_std_logic_vector(0, 8),
2307 => conv_std_logic_vector(0, 8),
2308 => conv_std_logic_vector(0, 8),
2309 => conv_std_logic_vector(0, 8),
2310 => conv_std_logic_vector(0, 8),
2311 => conv_std_logic_vector(0, 8),
2312 => conv_std_logic_vector(0, 8),
2313 => conv_std_logic_vector(0, 8),
2314 => conv_std_logic_vector(0, 8),
2315 => conv_std_logic_vector(0, 8),
2316 => conv_std_logic_vector(0, 8),
2317 => conv_std_logic_vector(0, 8),
2318 => conv_std_logic_vector(0, 8),
2319 => conv_std_logic_vector(0, 8),
2320 => conv_std_logic_vector(0, 8),
2321 => conv_std_logic_vector(0, 8),
2322 => conv_std_logic_vector(0, 8),
2323 => conv_std_logic_vector(0, 8),
2324 => conv_std_logic_vector(0, 8),
2325 => conv_std_logic_vector(0, 8),
2326 => conv_std_logic_vector(0, 8),
2327 => conv_std_logic_vector(0, 8),
2328 => conv_std_logic_vector(0, 8),
2329 => conv_std_logic_vector(0, 8),
2330 => conv_std_logic_vector(0, 8),
2331 => conv_std_logic_vector(0, 8),
2332 => conv_std_logic_vector(0, 8),
2333 => conv_std_logic_vector(1, 8),
2334 => conv_std_logic_vector(1, 8),
2335 => conv_std_logic_vector(1, 8),
2336 => conv_std_logic_vector(1, 8),
2337 => conv_std_logic_vector(1, 8),
2338 => conv_std_logic_vector(1, 8),
2339 => conv_std_logic_vector(1, 8),
2340 => conv_std_logic_vector(1, 8),
2341 => conv_std_logic_vector(1, 8),
2342 => conv_std_logic_vector(1, 8),
2343 => conv_std_logic_vector(1, 8),
2344 => conv_std_logic_vector(1, 8),
2345 => conv_std_logic_vector(1, 8),
2346 => conv_std_logic_vector(1, 8),
2347 => conv_std_logic_vector(1, 8),
2348 => conv_std_logic_vector(1, 8),
2349 => conv_std_logic_vector(1, 8),
2350 => conv_std_logic_vector(1, 8),
2351 => conv_std_logic_vector(1, 8),
2352 => conv_std_logic_vector(1, 8),
2353 => conv_std_logic_vector(1, 8),
2354 => conv_std_logic_vector(1, 8),
2355 => conv_std_logic_vector(1, 8),
2356 => conv_std_logic_vector(1, 8),
2357 => conv_std_logic_vector(1, 8),
2358 => conv_std_logic_vector(1, 8),
2359 => conv_std_logic_vector(1, 8),
2360 => conv_std_logic_vector(1, 8),
2361 => conv_std_logic_vector(2, 8),
2362 => conv_std_logic_vector(2, 8),
2363 => conv_std_logic_vector(2, 8),
2364 => conv_std_logic_vector(2, 8),
2365 => conv_std_logic_vector(2, 8),
2366 => conv_std_logic_vector(2, 8),
2367 => conv_std_logic_vector(2, 8),
2368 => conv_std_logic_vector(2, 8),
2369 => conv_std_logic_vector(2, 8),
2370 => conv_std_logic_vector(2, 8),
2371 => conv_std_logic_vector(2, 8),
2372 => conv_std_logic_vector(2, 8),
2373 => conv_std_logic_vector(2, 8),
2374 => conv_std_logic_vector(2, 8),
2375 => conv_std_logic_vector(2, 8),
2376 => conv_std_logic_vector(2, 8),
2377 => conv_std_logic_vector(2, 8),
2378 => conv_std_logic_vector(2, 8),
2379 => conv_std_logic_vector(2, 8),
2380 => conv_std_logic_vector(2, 8),
2381 => conv_std_logic_vector(2, 8),
2382 => conv_std_logic_vector(2, 8),
2383 => conv_std_logic_vector(2, 8),
2384 => conv_std_logic_vector(2, 8),
2385 => conv_std_logic_vector(2, 8),
2386 => conv_std_logic_vector(2, 8),
2387 => conv_std_logic_vector(2, 8),
2388 => conv_std_logic_vector(2, 8),
2389 => conv_std_logic_vector(2, 8),
2390 => conv_std_logic_vector(3, 8),
2391 => conv_std_logic_vector(3, 8),
2392 => conv_std_logic_vector(3, 8),
2393 => conv_std_logic_vector(3, 8),
2394 => conv_std_logic_vector(3, 8),
2395 => conv_std_logic_vector(3, 8),
2396 => conv_std_logic_vector(3, 8),
2397 => conv_std_logic_vector(3, 8),
2398 => conv_std_logic_vector(3, 8),
2399 => conv_std_logic_vector(3, 8),
2400 => conv_std_logic_vector(3, 8),
2401 => conv_std_logic_vector(3, 8),
2402 => conv_std_logic_vector(3, 8),
2403 => conv_std_logic_vector(3, 8),
2404 => conv_std_logic_vector(3, 8),
2405 => conv_std_logic_vector(3, 8),
2406 => conv_std_logic_vector(3, 8),
2407 => conv_std_logic_vector(3, 8),
2408 => conv_std_logic_vector(3, 8),
2409 => conv_std_logic_vector(3, 8),
2410 => conv_std_logic_vector(3, 8),
2411 => conv_std_logic_vector(3, 8),
2412 => conv_std_logic_vector(3, 8),
2413 => conv_std_logic_vector(3, 8),
2414 => conv_std_logic_vector(3, 8),
2415 => conv_std_logic_vector(3, 8),
2416 => conv_std_logic_vector(3, 8),
2417 => conv_std_logic_vector(3, 8),
2418 => conv_std_logic_vector(4, 8),
2419 => conv_std_logic_vector(4, 8),
2420 => conv_std_logic_vector(4, 8),
2421 => conv_std_logic_vector(4, 8),
2422 => conv_std_logic_vector(4, 8),
2423 => conv_std_logic_vector(4, 8),
2424 => conv_std_logic_vector(4, 8),
2425 => conv_std_logic_vector(4, 8),
2426 => conv_std_logic_vector(4, 8),
2427 => conv_std_logic_vector(4, 8),
2428 => conv_std_logic_vector(4, 8),
2429 => conv_std_logic_vector(4, 8),
2430 => conv_std_logic_vector(4, 8),
2431 => conv_std_logic_vector(4, 8),
2432 => conv_std_logic_vector(4, 8),
2433 => conv_std_logic_vector(4, 8),
2434 => conv_std_logic_vector(4, 8),
2435 => conv_std_logic_vector(4, 8),
2436 => conv_std_logic_vector(4, 8),
2437 => conv_std_logic_vector(4, 8),
2438 => conv_std_logic_vector(4, 8),
2439 => conv_std_logic_vector(4, 8),
2440 => conv_std_logic_vector(4, 8),
2441 => conv_std_logic_vector(4, 8),
2442 => conv_std_logic_vector(4, 8),
2443 => conv_std_logic_vector(4, 8),
2444 => conv_std_logic_vector(4, 8),
2445 => conv_std_logic_vector(4, 8),
2446 => conv_std_logic_vector(4, 8),
2447 => conv_std_logic_vector(5, 8),
2448 => conv_std_logic_vector(5, 8),
2449 => conv_std_logic_vector(5, 8),
2450 => conv_std_logic_vector(5, 8),
2451 => conv_std_logic_vector(5, 8),
2452 => conv_std_logic_vector(5, 8),
2453 => conv_std_logic_vector(5, 8),
2454 => conv_std_logic_vector(5, 8),
2455 => conv_std_logic_vector(5, 8),
2456 => conv_std_logic_vector(5, 8),
2457 => conv_std_logic_vector(5, 8),
2458 => conv_std_logic_vector(5, 8),
2459 => conv_std_logic_vector(5, 8),
2460 => conv_std_logic_vector(5, 8),
2461 => conv_std_logic_vector(5, 8),
2462 => conv_std_logic_vector(5, 8),
2463 => conv_std_logic_vector(5, 8),
2464 => conv_std_logic_vector(5, 8),
2465 => conv_std_logic_vector(5, 8),
2466 => conv_std_logic_vector(5, 8),
2467 => conv_std_logic_vector(5, 8),
2468 => conv_std_logic_vector(5, 8),
2469 => conv_std_logic_vector(5, 8),
2470 => conv_std_logic_vector(5, 8),
2471 => conv_std_logic_vector(5, 8),
2472 => conv_std_logic_vector(5, 8),
2473 => conv_std_logic_vector(5, 8),
2474 => conv_std_logic_vector(5, 8),
2475 => conv_std_logic_vector(6, 8),
2476 => conv_std_logic_vector(6, 8),
2477 => conv_std_logic_vector(6, 8),
2478 => conv_std_logic_vector(6, 8),
2479 => conv_std_logic_vector(6, 8),
2480 => conv_std_logic_vector(6, 8),
2481 => conv_std_logic_vector(6, 8),
2482 => conv_std_logic_vector(6, 8),
2483 => conv_std_logic_vector(6, 8),
2484 => conv_std_logic_vector(6, 8),
2485 => conv_std_logic_vector(6, 8),
2486 => conv_std_logic_vector(6, 8),
2487 => conv_std_logic_vector(6, 8),
2488 => conv_std_logic_vector(6, 8),
2489 => conv_std_logic_vector(6, 8),
2490 => conv_std_logic_vector(6, 8),
2491 => conv_std_logic_vector(6, 8),
2492 => conv_std_logic_vector(6, 8),
2493 => conv_std_logic_vector(6, 8),
2494 => conv_std_logic_vector(6, 8),
2495 => conv_std_logic_vector(6, 8),
2496 => conv_std_logic_vector(6, 8),
2497 => conv_std_logic_vector(6, 8),
2498 => conv_std_logic_vector(6, 8),
2499 => conv_std_logic_vector(6, 8),
2500 => conv_std_logic_vector(6, 8),
2501 => conv_std_logic_vector(6, 8),
2502 => conv_std_logic_vector(6, 8),
2503 => conv_std_logic_vector(6, 8),
2504 => conv_std_logic_vector(7, 8),
2505 => conv_std_logic_vector(7, 8),
2506 => conv_std_logic_vector(7, 8),
2507 => conv_std_logic_vector(7, 8),
2508 => conv_std_logic_vector(7, 8),
2509 => conv_std_logic_vector(7, 8),
2510 => conv_std_logic_vector(7, 8),
2511 => conv_std_logic_vector(7, 8),
2512 => conv_std_logic_vector(7, 8),
2513 => conv_std_logic_vector(7, 8),
2514 => conv_std_logic_vector(7, 8),
2515 => conv_std_logic_vector(7, 8),
2516 => conv_std_logic_vector(7, 8),
2517 => conv_std_logic_vector(7, 8),
2518 => conv_std_logic_vector(7, 8),
2519 => conv_std_logic_vector(7, 8),
2520 => conv_std_logic_vector(7, 8),
2521 => conv_std_logic_vector(7, 8),
2522 => conv_std_logic_vector(7, 8),
2523 => conv_std_logic_vector(7, 8),
2524 => conv_std_logic_vector(7, 8),
2525 => conv_std_logic_vector(7, 8),
2526 => conv_std_logic_vector(7, 8),
2527 => conv_std_logic_vector(7, 8),
2528 => conv_std_logic_vector(7, 8),
2529 => conv_std_logic_vector(7, 8),
2530 => conv_std_logic_vector(7, 8),
2531 => conv_std_logic_vector(7, 8),
2532 => conv_std_logic_vector(8, 8),
2533 => conv_std_logic_vector(8, 8),
2534 => conv_std_logic_vector(8, 8),
2535 => conv_std_logic_vector(8, 8),
2536 => conv_std_logic_vector(8, 8),
2537 => conv_std_logic_vector(8, 8),
2538 => conv_std_logic_vector(8, 8),
2539 => conv_std_logic_vector(8, 8),
2540 => conv_std_logic_vector(8, 8),
2541 => conv_std_logic_vector(8, 8),
2542 => conv_std_logic_vector(8, 8),
2543 => conv_std_logic_vector(8, 8),
2544 => conv_std_logic_vector(8, 8),
2545 => conv_std_logic_vector(8, 8),
2546 => conv_std_logic_vector(8, 8),
2547 => conv_std_logic_vector(8, 8),
2548 => conv_std_logic_vector(8, 8),
2549 => conv_std_logic_vector(8, 8),
2550 => conv_std_logic_vector(8, 8),
2551 => conv_std_logic_vector(8, 8),
2552 => conv_std_logic_vector(8, 8),
2553 => conv_std_logic_vector(8, 8),
2554 => conv_std_logic_vector(8, 8),
2555 => conv_std_logic_vector(8, 8),
2556 => conv_std_logic_vector(8, 8),
2557 => conv_std_logic_vector(8, 8),
2558 => conv_std_logic_vector(8, 8),
2559 => conv_std_logic_vector(8, 8),
2560 => conv_std_logic_vector(0, 8),
2561 => conv_std_logic_vector(0, 8),
2562 => conv_std_logic_vector(0, 8),
2563 => conv_std_logic_vector(0, 8),
2564 => conv_std_logic_vector(0, 8),
2565 => conv_std_logic_vector(0, 8),
2566 => conv_std_logic_vector(0, 8),
2567 => conv_std_logic_vector(0, 8),
2568 => conv_std_logic_vector(0, 8),
2569 => conv_std_logic_vector(0, 8),
2570 => conv_std_logic_vector(0, 8),
2571 => conv_std_logic_vector(0, 8),
2572 => conv_std_logic_vector(0, 8),
2573 => conv_std_logic_vector(0, 8),
2574 => conv_std_logic_vector(0, 8),
2575 => conv_std_logic_vector(0, 8),
2576 => conv_std_logic_vector(0, 8),
2577 => conv_std_logic_vector(0, 8),
2578 => conv_std_logic_vector(0, 8),
2579 => conv_std_logic_vector(0, 8),
2580 => conv_std_logic_vector(0, 8),
2581 => conv_std_logic_vector(0, 8),
2582 => conv_std_logic_vector(0, 8),
2583 => conv_std_logic_vector(0, 8),
2584 => conv_std_logic_vector(0, 8),
2585 => conv_std_logic_vector(0, 8),
2586 => conv_std_logic_vector(1, 8),
2587 => conv_std_logic_vector(1, 8),
2588 => conv_std_logic_vector(1, 8),
2589 => conv_std_logic_vector(1, 8),
2590 => conv_std_logic_vector(1, 8),
2591 => conv_std_logic_vector(1, 8),
2592 => conv_std_logic_vector(1, 8),
2593 => conv_std_logic_vector(1, 8),
2594 => conv_std_logic_vector(1, 8),
2595 => conv_std_logic_vector(1, 8),
2596 => conv_std_logic_vector(1, 8),
2597 => conv_std_logic_vector(1, 8),
2598 => conv_std_logic_vector(1, 8),
2599 => conv_std_logic_vector(1, 8),
2600 => conv_std_logic_vector(1, 8),
2601 => conv_std_logic_vector(1, 8),
2602 => conv_std_logic_vector(1, 8),
2603 => conv_std_logic_vector(1, 8),
2604 => conv_std_logic_vector(1, 8),
2605 => conv_std_logic_vector(1, 8),
2606 => conv_std_logic_vector(1, 8),
2607 => conv_std_logic_vector(1, 8),
2608 => conv_std_logic_vector(1, 8),
2609 => conv_std_logic_vector(1, 8),
2610 => conv_std_logic_vector(1, 8),
2611 => conv_std_logic_vector(1, 8),
2612 => conv_std_logic_vector(2, 8),
2613 => conv_std_logic_vector(2, 8),
2614 => conv_std_logic_vector(2, 8),
2615 => conv_std_logic_vector(2, 8),
2616 => conv_std_logic_vector(2, 8),
2617 => conv_std_logic_vector(2, 8),
2618 => conv_std_logic_vector(2, 8),
2619 => conv_std_logic_vector(2, 8),
2620 => conv_std_logic_vector(2, 8),
2621 => conv_std_logic_vector(2, 8),
2622 => conv_std_logic_vector(2, 8),
2623 => conv_std_logic_vector(2, 8),
2624 => conv_std_logic_vector(2, 8),
2625 => conv_std_logic_vector(2, 8),
2626 => conv_std_logic_vector(2, 8),
2627 => conv_std_logic_vector(2, 8),
2628 => conv_std_logic_vector(2, 8),
2629 => conv_std_logic_vector(2, 8),
2630 => conv_std_logic_vector(2, 8),
2631 => conv_std_logic_vector(2, 8),
2632 => conv_std_logic_vector(2, 8),
2633 => conv_std_logic_vector(2, 8),
2634 => conv_std_logic_vector(2, 8),
2635 => conv_std_logic_vector(2, 8),
2636 => conv_std_logic_vector(2, 8),
2637 => conv_std_logic_vector(3, 8),
2638 => conv_std_logic_vector(3, 8),
2639 => conv_std_logic_vector(3, 8),
2640 => conv_std_logic_vector(3, 8),
2641 => conv_std_logic_vector(3, 8),
2642 => conv_std_logic_vector(3, 8),
2643 => conv_std_logic_vector(3, 8),
2644 => conv_std_logic_vector(3, 8),
2645 => conv_std_logic_vector(3, 8),
2646 => conv_std_logic_vector(3, 8),
2647 => conv_std_logic_vector(3, 8),
2648 => conv_std_logic_vector(3, 8),
2649 => conv_std_logic_vector(3, 8),
2650 => conv_std_logic_vector(3, 8),
2651 => conv_std_logic_vector(3, 8),
2652 => conv_std_logic_vector(3, 8),
2653 => conv_std_logic_vector(3, 8),
2654 => conv_std_logic_vector(3, 8),
2655 => conv_std_logic_vector(3, 8),
2656 => conv_std_logic_vector(3, 8),
2657 => conv_std_logic_vector(3, 8),
2658 => conv_std_logic_vector(3, 8),
2659 => conv_std_logic_vector(3, 8),
2660 => conv_std_logic_vector(3, 8),
2661 => conv_std_logic_vector(3, 8),
2662 => conv_std_logic_vector(3, 8),
2663 => conv_std_logic_vector(4, 8),
2664 => conv_std_logic_vector(4, 8),
2665 => conv_std_logic_vector(4, 8),
2666 => conv_std_logic_vector(4, 8),
2667 => conv_std_logic_vector(4, 8),
2668 => conv_std_logic_vector(4, 8),
2669 => conv_std_logic_vector(4, 8),
2670 => conv_std_logic_vector(4, 8),
2671 => conv_std_logic_vector(4, 8),
2672 => conv_std_logic_vector(4, 8),
2673 => conv_std_logic_vector(4, 8),
2674 => conv_std_logic_vector(4, 8),
2675 => conv_std_logic_vector(4, 8),
2676 => conv_std_logic_vector(4, 8),
2677 => conv_std_logic_vector(4, 8),
2678 => conv_std_logic_vector(4, 8),
2679 => conv_std_logic_vector(4, 8),
2680 => conv_std_logic_vector(4, 8),
2681 => conv_std_logic_vector(4, 8),
2682 => conv_std_logic_vector(4, 8),
2683 => conv_std_logic_vector(4, 8),
2684 => conv_std_logic_vector(4, 8),
2685 => conv_std_logic_vector(4, 8),
2686 => conv_std_logic_vector(4, 8),
2687 => conv_std_logic_vector(4, 8),
2688 => conv_std_logic_vector(5, 8),
2689 => conv_std_logic_vector(5, 8),
2690 => conv_std_logic_vector(5, 8),
2691 => conv_std_logic_vector(5, 8),
2692 => conv_std_logic_vector(5, 8),
2693 => conv_std_logic_vector(5, 8),
2694 => conv_std_logic_vector(5, 8),
2695 => conv_std_logic_vector(5, 8),
2696 => conv_std_logic_vector(5, 8),
2697 => conv_std_logic_vector(5, 8),
2698 => conv_std_logic_vector(5, 8),
2699 => conv_std_logic_vector(5, 8),
2700 => conv_std_logic_vector(5, 8),
2701 => conv_std_logic_vector(5, 8),
2702 => conv_std_logic_vector(5, 8),
2703 => conv_std_logic_vector(5, 8),
2704 => conv_std_logic_vector(5, 8),
2705 => conv_std_logic_vector(5, 8),
2706 => conv_std_logic_vector(5, 8),
2707 => conv_std_logic_vector(5, 8),
2708 => conv_std_logic_vector(5, 8),
2709 => conv_std_logic_vector(5, 8),
2710 => conv_std_logic_vector(5, 8),
2711 => conv_std_logic_vector(5, 8),
2712 => conv_std_logic_vector(5, 8),
2713 => conv_std_logic_vector(5, 8),
2714 => conv_std_logic_vector(6, 8),
2715 => conv_std_logic_vector(6, 8),
2716 => conv_std_logic_vector(6, 8),
2717 => conv_std_logic_vector(6, 8),
2718 => conv_std_logic_vector(6, 8),
2719 => conv_std_logic_vector(6, 8),
2720 => conv_std_logic_vector(6, 8),
2721 => conv_std_logic_vector(6, 8),
2722 => conv_std_logic_vector(6, 8),
2723 => conv_std_logic_vector(6, 8),
2724 => conv_std_logic_vector(6, 8),
2725 => conv_std_logic_vector(6, 8),
2726 => conv_std_logic_vector(6, 8),
2727 => conv_std_logic_vector(6, 8),
2728 => conv_std_logic_vector(6, 8),
2729 => conv_std_logic_vector(6, 8),
2730 => conv_std_logic_vector(6, 8),
2731 => conv_std_logic_vector(6, 8),
2732 => conv_std_logic_vector(6, 8),
2733 => conv_std_logic_vector(6, 8),
2734 => conv_std_logic_vector(6, 8),
2735 => conv_std_logic_vector(6, 8),
2736 => conv_std_logic_vector(6, 8),
2737 => conv_std_logic_vector(6, 8),
2738 => conv_std_logic_vector(6, 8),
2739 => conv_std_logic_vector(6, 8),
2740 => conv_std_logic_vector(7, 8),
2741 => conv_std_logic_vector(7, 8),
2742 => conv_std_logic_vector(7, 8),
2743 => conv_std_logic_vector(7, 8),
2744 => conv_std_logic_vector(7, 8),
2745 => conv_std_logic_vector(7, 8),
2746 => conv_std_logic_vector(7, 8),
2747 => conv_std_logic_vector(7, 8),
2748 => conv_std_logic_vector(7, 8),
2749 => conv_std_logic_vector(7, 8),
2750 => conv_std_logic_vector(7, 8),
2751 => conv_std_logic_vector(7, 8),
2752 => conv_std_logic_vector(7, 8),
2753 => conv_std_logic_vector(7, 8),
2754 => conv_std_logic_vector(7, 8),
2755 => conv_std_logic_vector(7, 8),
2756 => conv_std_logic_vector(7, 8),
2757 => conv_std_logic_vector(7, 8),
2758 => conv_std_logic_vector(7, 8),
2759 => conv_std_logic_vector(7, 8),
2760 => conv_std_logic_vector(7, 8),
2761 => conv_std_logic_vector(7, 8),
2762 => conv_std_logic_vector(7, 8),
2763 => conv_std_logic_vector(7, 8),
2764 => conv_std_logic_vector(7, 8),
2765 => conv_std_logic_vector(8, 8),
2766 => conv_std_logic_vector(8, 8),
2767 => conv_std_logic_vector(8, 8),
2768 => conv_std_logic_vector(8, 8),
2769 => conv_std_logic_vector(8, 8),
2770 => conv_std_logic_vector(8, 8),
2771 => conv_std_logic_vector(8, 8),
2772 => conv_std_logic_vector(8, 8),
2773 => conv_std_logic_vector(8, 8),
2774 => conv_std_logic_vector(8, 8),
2775 => conv_std_logic_vector(8, 8),
2776 => conv_std_logic_vector(8, 8),
2777 => conv_std_logic_vector(8, 8),
2778 => conv_std_logic_vector(8, 8),
2779 => conv_std_logic_vector(8, 8),
2780 => conv_std_logic_vector(8, 8),
2781 => conv_std_logic_vector(8, 8),
2782 => conv_std_logic_vector(8, 8),
2783 => conv_std_logic_vector(8, 8),
2784 => conv_std_logic_vector(8, 8),
2785 => conv_std_logic_vector(8, 8),
2786 => conv_std_logic_vector(8, 8),
2787 => conv_std_logic_vector(8, 8),
2788 => conv_std_logic_vector(8, 8),
2789 => conv_std_logic_vector(8, 8),
2790 => conv_std_logic_vector(8, 8),
2791 => conv_std_logic_vector(9, 8),
2792 => conv_std_logic_vector(9, 8),
2793 => conv_std_logic_vector(9, 8),
2794 => conv_std_logic_vector(9, 8),
2795 => conv_std_logic_vector(9, 8),
2796 => conv_std_logic_vector(9, 8),
2797 => conv_std_logic_vector(9, 8),
2798 => conv_std_logic_vector(9, 8),
2799 => conv_std_logic_vector(9, 8),
2800 => conv_std_logic_vector(9, 8),
2801 => conv_std_logic_vector(9, 8),
2802 => conv_std_logic_vector(9, 8),
2803 => conv_std_logic_vector(9, 8),
2804 => conv_std_logic_vector(9, 8),
2805 => conv_std_logic_vector(9, 8),
2806 => conv_std_logic_vector(9, 8),
2807 => conv_std_logic_vector(9, 8),
2808 => conv_std_logic_vector(9, 8),
2809 => conv_std_logic_vector(9, 8),
2810 => conv_std_logic_vector(9, 8),
2811 => conv_std_logic_vector(9, 8),
2812 => conv_std_logic_vector(9, 8),
2813 => conv_std_logic_vector(9, 8),
2814 => conv_std_logic_vector(9, 8),
2815 => conv_std_logic_vector(9, 8),
2816 => conv_std_logic_vector(0, 8),
2817 => conv_std_logic_vector(0, 8),
2818 => conv_std_logic_vector(0, 8),
2819 => conv_std_logic_vector(0, 8),
2820 => conv_std_logic_vector(0, 8),
2821 => conv_std_logic_vector(0, 8),
2822 => conv_std_logic_vector(0, 8),
2823 => conv_std_logic_vector(0, 8),
2824 => conv_std_logic_vector(0, 8),
2825 => conv_std_logic_vector(0, 8),
2826 => conv_std_logic_vector(0, 8),
2827 => conv_std_logic_vector(0, 8),
2828 => conv_std_logic_vector(0, 8),
2829 => conv_std_logic_vector(0, 8),
2830 => conv_std_logic_vector(0, 8),
2831 => conv_std_logic_vector(0, 8),
2832 => conv_std_logic_vector(0, 8),
2833 => conv_std_logic_vector(0, 8),
2834 => conv_std_logic_vector(0, 8),
2835 => conv_std_logic_vector(0, 8),
2836 => conv_std_logic_vector(0, 8),
2837 => conv_std_logic_vector(0, 8),
2838 => conv_std_logic_vector(0, 8),
2839 => conv_std_logic_vector(0, 8),
2840 => conv_std_logic_vector(1, 8),
2841 => conv_std_logic_vector(1, 8),
2842 => conv_std_logic_vector(1, 8),
2843 => conv_std_logic_vector(1, 8),
2844 => conv_std_logic_vector(1, 8),
2845 => conv_std_logic_vector(1, 8),
2846 => conv_std_logic_vector(1, 8),
2847 => conv_std_logic_vector(1, 8),
2848 => conv_std_logic_vector(1, 8),
2849 => conv_std_logic_vector(1, 8),
2850 => conv_std_logic_vector(1, 8),
2851 => conv_std_logic_vector(1, 8),
2852 => conv_std_logic_vector(1, 8),
2853 => conv_std_logic_vector(1, 8),
2854 => conv_std_logic_vector(1, 8),
2855 => conv_std_logic_vector(1, 8),
2856 => conv_std_logic_vector(1, 8),
2857 => conv_std_logic_vector(1, 8),
2858 => conv_std_logic_vector(1, 8),
2859 => conv_std_logic_vector(1, 8),
2860 => conv_std_logic_vector(1, 8),
2861 => conv_std_logic_vector(1, 8),
2862 => conv_std_logic_vector(1, 8),
2863 => conv_std_logic_vector(2, 8),
2864 => conv_std_logic_vector(2, 8),
2865 => conv_std_logic_vector(2, 8),
2866 => conv_std_logic_vector(2, 8),
2867 => conv_std_logic_vector(2, 8),
2868 => conv_std_logic_vector(2, 8),
2869 => conv_std_logic_vector(2, 8),
2870 => conv_std_logic_vector(2, 8),
2871 => conv_std_logic_vector(2, 8),
2872 => conv_std_logic_vector(2, 8),
2873 => conv_std_logic_vector(2, 8),
2874 => conv_std_logic_vector(2, 8),
2875 => conv_std_logic_vector(2, 8),
2876 => conv_std_logic_vector(2, 8),
2877 => conv_std_logic_vector(2, 8),
2878 => conv_std_logic_vector(2, 8),
2879 => conv_std_logic_vector(2, 8),
2880 => conv_std_logic_vector(2, 8),
2881 => conv_std_logic_vector(2, 8),
2882 => conv_std_logic_vector(2, 8),
2883 => conv_std_logic_vector(2, 8),
2884 => conv_std_logic_vector(2, 8),
2885 => conv_std_logic_vector(2, 8),
2886 => conv_std_logic_vector(3, 8),
2887 => conv_std_logic_vector(3, 8),
2888 => conv_std_logic_vector(3, 8),
2889 => conv_std_logic_vector(3, 8),
2890 => conv_std_logic_vector(3, 8),
2891 => conv_std_logic_vector(3, 8),
2892 => conv_std_logic_vector(3, 8),
2893 => conv_std_logic_vector(3, 8),
2894 => conv_std_logic_vector(3, 8),
2895 => conv_std_logic_vector(3, 8),
2896 => conv_std_logic_vector(3, 8),
2897 => conv_std_logic_vector(3, 8),
2898 => conv_std_logic_vector(3, 8),
2899 => conv_std_logic_vector(3, 8),
2900 => conv_std_logic_vector(3, 8),
2901 => conv_std_logic_vector(3, 8),
2902 => conv_std_logic_vector(3, 8),
2903 => conv_std_logic_vector(3, 8),
2904 => conv_std_logic_vector(3, 8),
2905 => conv_std_logic_vector(3, 8),
2906 => conv_std_logic_vector(3, 8),
2907 => conv_std_logic_vector(3, 8),
2908 => conv_std_logic_vector(3, 8),
2909 => conv_std_logic_vector(3, 8),
2910 => conv_std_logic_vector(4, 8),
2911 => conv_std_logic_vector(4, 8),
2912 => conv_std_logic_vector(4, 8),
2913 => conv_std_logic_vector(4, 8),
2914 => conv_std_logic_vector(4, 8),
2915 => conv_std_logic_vector(4, 8),
2916 => conv_std_logic_vector(4, 8),
2917 => conv_std_logic_vector(4, 8),
2918 => conv_std_logic_vector(4, 8),
2919 => conv_std_logic_vector(4, 8),
2920 => conv_std_logic_vector(4, 8),
2921 => conv_std_logic_vector(4, 8),
2922 => conv_std_logic_vector(4, 8),
2923 => conv_std_logic_vector(4, 8),
2924 => conv_std_logic_vector(4, 8),
2925 => conv_std_logic_vector(4, 8),
2926 => conv_std_logic_vector(4, 8),
2927 => conv_std_logic_vector(4, 8),
2928 => conv_std_logic_vector(4, 8),
2929 => conv_std_logic_vector(4, 8),
2930 => conv_std_logic_vector(4, 8),
2931 => conv_std_logic_vector(4, 8),
2932 => conv_std_logic_vector(4, 8),
2933 => conv_std_logic_vector(5, 8),
2934 => conv_std_logic_vector(5, 8),
2935 => conv_std_logic_vector(5, 8),
2936 => conv_std_logic_vector(5, 8),
2937 => conv_std_logic_vector(5, 8),
2938 => conv_std_logic_vector(5, 8),
2939 => conv_std_logic_vector(5, 8),
2940 => conv_std_logic_vector(5, 8),
2941 => conv_std_logic_vector(5, 8),
2942 => conv_std_logic_vector(5, 8),
2943 => conv_std_logic_vector(5, 8),
2944 => conv_std_logic_vector(5, 8),
2945 => conv_std_logic_vector(5, 8),
2946 => conv_std_logic_vector(5, 8),
2947 => conv_std_logic_vector(5, 8),
2948 => conv_std_logic_vector(5, 8),
2949 => conv_std_logic_vector(5, 8),
2950 => conv_std_logic_vector(5, 8),
2951 => conv_std_logic_vector(5, 8),
2952 => conv_std_logic_vector(5, 8),
2953 => conv_std_logic_vector(5, 8),
2954 => conv_std_logic_vector(5, 8),
2955 => conv_std_logic_vector(5, 8),
2956 => conv_std_logic_vector(6, 8),
2957 => conv_std_logic_vector(6, 8),
2958 => conv_std_logic_vector(6, 8),
2959 => conv_std_logic_vector(6, 8),
2960 => conv_std_logic_vector(6, 8),
2961 => conv_std_logic_vector(6, 8),
2962 => conv_std_logic_vector(6, 8),
2963 => conv_std_logic_vector(6, 8),
2964 => conv_std_logic_vector(6, 8),
2965 => conv_std_logic_vector(6, 8),
2966 => conv_std_logic_vector(6, 8),
2967 => conv_std_logic_vector(6, 8),
2968 => conv_std_logic_vector(6, 8),
2969 => conv_std_logic_vector(6, 8),
2970 => conv_std_logic_vector(6, 8),
2971 => conv_std_logic_vector(6, 8),
2972 => conv_std_logic_vector(6, 8),
2973 => conv_std_logic_vector(6, 8),
2974 => conv_std_logic_vector(6, 8),
2975 => conv_std_logic_vector(6, 8),
2976 => conv_std_logic_vector(6, 8),
2977 => conv_std_logic_vector(6, 8),
2978 => conv_std_logic_vector(6, 8),
2979 => conv_std_logic_vector(7, 8),
2980 => conv_std_logic_vector(7, 8),
2981 => conv_std_logic_vector(7, 8),
2982 => conv_std_logic_vector(7, 8),
2983 => conv_std_logic_vector(7, 8),
2984 => conv_std_logic_vector(7, 8),
2985 => conv_std_logic_vector(7, 8),
2986 => conv_std_logic_vector(7, 8),
2987 => conv_std_logic_vector(7, 8),
2988 => conv_std_logic_vector(7, 8),
2989 => conv_std_logic_vector(7, 8),
2990 => conv_std_logic_vector(7, 8),
2991 => conv_std_logic_vector(7, 8),
2992 => conv_std_logic_vector(7, 8),
2993 => conv_std_logic_vector(7, 8),
2994 => conv_std_logic_vector(7, 8),
2995 => conv_std_logic_vector(7, 8),
2996 => conv_std_logic_vector(7, 8),
2997 => conv_std_logic_vector(7, 8),
2998 => conv_std_logic_vector(7, 8),
2999 => conv_std_logic_vector(7, 8),
3000 => conv_std_logic_vector(7, 8),
3001 => conv_std_logic_vector(7, 8),
3002 => conv_std_logic_vector(7, 8),
3003 => conv_std_logic_vector(8, 8),
3004 => conv_std_logic_vector(8, 8),
3005 => conv_std_logic_vector(8, 8),
3006 => conv_std_logic_vector(8, 8),
3007 => conv_std_logic_vector(8, 8),
3008 => conv_std_logic_vector(8, 8),
3009 => conv_std_logic_vector(8, 8),
3010 => conv_std_logic_vector(8, 8),
3011 => conv_std_logic_vector(8, 8),
3012 => conv_std_logic_vector(8, 8),
3013 => conv_std_logic_vector(8, 8),
3014 => conv_std_logic_vector(8, 8),
3015 => conv_std_logic_vector(8, 8),
3016 => conv_std_logic_vector(8, 8),
3017 => conv_std_logic_vector(8, 8),
3018 => conv_std_logic_vector(8, 8),
3019 => conv_std_logic_vector(8, 8),
3020 => conv_std_logic_vector(8, 8),
3021 => conv_std_logic_vector(8, 8),
3022 => conv_std_logic_vector(8, 8),
3023 => conv_std_logic_vector(8, 8),
3024 => conv_std_logic_vector(8, 8),
3025 => conv_std_logic_vector(8, 8),
3026 => conv_std_logic_vector(9, 8),
3027 => conv_std_logic_vector(9, 8),
3028 => conv_std_logic_vector(9, 8),
3029 => conv_std_logic_vector(9, 8),
3030 => conv_std_logic_vector(9, 8),
3031 => conv_std_logic_vector(9, 8),
3032 => conv_std_logic_vector(9, 8),
3033 => conv_std_logic_vector(9, 8),
3034 => conv_std_logic_vector(9, 8),
3035 => conv_std_logic_vector(9, 8),
3036 => conv_std_logic_vector(9, 8),
3037 => conv_std_logic_vector(9, 8),
3038 => conv_std_logic_vector(9, 8),
3039 => conv_std_logic_vector(9, 8),
3040 => conv_std_logic_vector(9, 8),
3041 => conv_std_logic_vector(9, 8),
3042 => conv_std_logic_vector(9, 8),
3043 => conv_std_logic_vector(9, 8),
3044 => conv_std_logic_vector(9, 8),
3045 => conv_std_logic_vector(9, 8),
3046 => conv_std_logic_vector(9, 8),
3047 => conv_std_logic_vector(9, 8),
3048 => conv_std_logic_vector(9, 8),
3049 => conv_std_logic_vector(10, 8),
3050 => conv_std_logic_vector(10, 8),
3051 => conv_std_logic_vector(10, 8),
3052 => conv_std_logic_vector(10, 8),
3053 => conv_std_logic_vector(10, 8),
3054 => conv_std_logic_vector(10, 8),
3055 => conv_std_logic_vector(10, 8),
3056 => conv_std_logic_vector(10, 8),
3057 => conv_std_logic_vector(10, 8),
3058 => conv_std_logic_vector(10, 8),
3059 => conv_std_logic_vector(10, 8),
3060 => conv_std_logic_vector(10, 8),
3061 => conv_std_logic_vector(10, 8),
3062 => conv_std_logic_vector(10, 8),
3063 => conv_std_logic_vector(10, 8),
3064 => conv_std_logic_vector(10, 8),
3065 => conv_std_logic_vector(10, 8),
3066 => conv_std_logic_vector(10, 8),
3067 => conv_std_logic_vector(10, 8),
3068 => conv_std_logic_vector(10, 8),
3069 => conv_std_logic_vector(10, 8),
3070 => conv_std_logic_vector(10, 8),
3071 => conv_std_logic_vector(10, 8),
3072 => conv_std_logic_vector(0, 8),
3073 => conv_std_logic_vector(0, 8),
3074 => conv_std_logic_vector(0, 8),
3075 => conv_std_logic_vector(0, 8),
3076 => conv_std_logic_vector(0, 8),
3077 => conv_std_logic_vector(0, 8),
3078 => conv_std_logic_vector(0, 8),
3079 => conv_std_logic_vector(0, 8),
3080 => conv_std_logic_vector(0, 8),
3081 => conv_std_logic_vector(0, 8),
3082 => conv_std_logic_vector(0, 8),
3083 => conv_std_logic_vector(0, 8),
3084 => conv_std_logic_vector(0, 8),
3085 => conv_std_logic_vector(0, 8),
3086 => conv_std_logic_vector(0, 8),
3087 => conv_std_logic_vector(0, 8),
3088 => conv_std_logic_vector(0, 8),
3089 => conv_std_logic_vector(0, 8),
3090 => conv_std_logic_vector(0, 8),
3091 => conv_std_logic_vector(0, 8),
3092 => conv_std_logic_vector(0, 8),
3093 => conv_std_logic_vector(0, 8),
3094 => conv_std_logic_vector(1, 8),
3095 => conv_std_logic_vector(1, 8),
3096 => conv_std_logic_vector(1, 8),
3097 => conv_std_logic_vector(1, 8),
3098 => conv_std_logic_vector(1, 8),
3099 => conv_std_logic_vector(1, 8),
3100 => conv_std_logic_vector(1, 8),
3101 => conv_std_logic_vector(1, 8),
3102 => conv_std_logic_vector(1, 8),
3103 => conv_std_logic_vector(1, 8),
3104 => conv_std_logic_vector(1, 8),
3105 => conv_std_logic_vector(1, 8),
3106 => conv_std_logic_vector(1, 8),
3107 => conv_std_logic_vector(1, 8),
3108 => conv_std_logic_vector(1, 8),
3109 => conv_std_logic_vector(1, 8),
3110 => conv_std_logic_vector(1, 8),
3111 => conv_std_logic_vector(1, 8),
3112 => conv_std_logic_vector(1, 8),
3113 => conv_std_logic_vector(1, 8),
3114 => conv_std_logic_vector(1, 8),
3115 => conv_std_logic_vector(2, 8),
3116 => conv_std_logic_vector(2, 8),
3117 => conv_std_logic_vector(2, 8),
3118 => conv_std_logic_vector(2, 8),
3119 => conv_std_logic_vector(2, 8),
3120 => conv_std_logic_vector(2, 8),
3121 => conv_std_logic_vector(2, 8),
3122 => conv_std_logic_vector(2, 8),
3123 => conv_std_logic_vector(2, 8),
3124 => conv_std_logic_vector(2, 8),
3125 => conv_std_logic_vector(2, 8),
3126 => conv_std_logic_vector(2, 8),
3127 => conv_std_logic_vector(2, 8),
3128 => conv_std_logic_vector(2, 8),
3129 => conv_std_logic_vector(2, 8),
3130 => conv_std_logic_vector(2, 8),
3131 => conv_std_logic_vector(2, 8),
3132 => conv_std_logic_vector(2, 8),
3133 => conv_std_logic_vector(2, 8),
3134 => conv_std_logic_vector(2, 8),
3135 => conv_std_logic_vector(2, 8),
3136 => conv_std_logic_vector(3, 8),
3137 => conv_std_logic_vector(3, 8),
3138 => conv_std_logic_vector(3, 8),
3139 => conv_std_logic_vector(3, 8),
3140 => conv_std_logic_vector(3, 8),
3141 => conv_std_logic_vector(3, 8),
3142 => conv_std_logic_vector(3, 8),
3143 => conv_std_logic_vector(3, 8),
3144 => conv_std_logic_vector(3, 8),
3145 => conv_std_logic_vector(3, 8),
3146 => conv_std_logic_vector(3, 8),
3147 => conv_std_logic_vector(3, 8),
3148 => conv_std_logic_vector(3, 8),
3149 => conv_std_logic_vector(3, 8),
3150 => conv_std_logic_vector(3, 8),
3151 => conv_std_logic_vector(3, 8),
3152 => conv_std_logic_vector(3, 8),
3153 => conv_std_logic_vector(3, 8),
3154 => conv_std_logic_vector(3, 8),
3155 => conv_std_logic_vector(3, 8),
3156 => conv_std_logic_vector(3, 8),
3157 => conv_std_logic_vector(3, 8),
3158 => conv_std_logic_vector(4, 8),
3159 => conv_std_logic_vector(4, 8),
3160 => conv_std_logic_vector(4, 8),
3161 => conv_std_logic_vector(4, 8),
3162 => conv_std_logic_vector(4, 8),
3163 => conv_std_logic_vector(4, 8),
3164 => conv_std_logic_vector(4, 8),
3165 => conv_std_logic_vector(4, 8),
3166 => conv_std_logic_vector(4, 8),
3167 => conv_std_logic_vector(4, 8),
3168 => conv_std_logic_vector(4, 8),
3169 => conv_std_logic_vector(4, 8),
3170 => conv_std_logic_vector(4, 8),
3171 => conv_std_logic_vector(4, 8),
3172 => conv_std_logic_vector(4, 8),
3173 => conv_std_logic_vector(4, 8),
3174 => conv_std_logic_vector(4, 8),
3175 => conv_std_logic_vector(4, 8),
3176 => conv_std_logic_vector(4, 8),
3177 => conv_std_logic_vector(4, 8),
3178 => conv_std_logic_vector(4, 8),
3179 => conv_std_logic_vector(5, 8),
3180 => conv_std_logic_vector(5, 8),
3181 => conv_std_logic_vector(5, 8),
3182 => conv_std_logic_vector(5, 8),
3183 => conv_std_logic_vector(5, 8),
3184 => conv_std_logic_vector(5, 8),
3185 => conv_std_logic_vector(5, 8),
3186 => conv_std_logic_vector(5, 8),
3187 => conv_std_logic_vector(5, 8),
3188 => conv_std_logic_vector(5, 8),
3189 => conv_std_logic_vector(5, 8),
3190 => conv_std_logic_vector(5, 8),
3191 => conv_std_logic_vector(5, 8),
3192 => conv_std_logic_vector(5, 8),
3193 => conv_std_logic_vector(5, 8),
3194 => conv_std_logic_vector(5, 8),
3195 => conv_std_logic_vector(5, 8),
3196 => conv_std_logic_vector(5, 8),
3197 => conv_std_logic_vector(5, 8),
3198 => conv_std_logic_vector(5, 8),
3199 => conv_std_logic_vector(5, 8),
3200 => conv_std_logic_vector(6, 8),
3201 => conv_std_logic_vector(6, 8),
3202 => conv_std_logic_vector(6, 8),
3203 => conv_std_logic_vector(6, 8),
3204 => conv_std_logic_vector(6, 8),
3205 => conv_std_logic_vector(6, 8),
3206 => conv_std_logic_vector(6, 8),
3207 => conv_std_logic_vector(6, 8),
3208 => conv_std_logic_vector(6, 8),
3209 => conv_std_logic_vector(6, 8),
3210 => conv_std_logic_vector(6, 8),
3211 => conv_std_logic_vector(6, 8),
3212 => conv_std_logic_vector(6, 8),
3213 => conv_std_logic_vector(6, 8),
3214 => conv_std_logic_vector(6, 8),
3215 => conv_std_logic_vector(6, 8),
3216 => conv_std_logic_vector(6, 8),
3217 => conv_std_logic_vector(6, 8),
3218 => conv_std_logic_vector(6, 8),
3219 => conv_std_logic_vector(6, 8),
3220 => conv_std_logic_vector(6, 8),
3221 => conv_std_logic_vector(6, 8),
3222 => conv_std_logic_vector(7, 8),
3223 => conv_std_logic_vector(7, 8),
3224 => conv_std_logic_vector(7, 8),
3225 => conv_std_logic_vector(7, 8),
3226 => conv_std_logic_vector(7, 8),
3227 => conv_std_logic_vector(7, 8),
3228 => conv_std_logic_vector(7, 8),
3229 => conv_std_logic_vector(7, 8),
3230 => conv_std_logic_vector(7, 8),
3231 => conv_std_logic_vector(7, 8),
3232 => conv_std_logic_vector(7, 8),
3233 => conv_std_logic_vector(7, 8),
3234 => conv_std_logic_vector(7, 8),
3235 => conv_std_logic_vector(7, 8),
3236 => conv_std_logic_vector(7, 8),
3237 => conv_std_logic_vector(7, 8),
3238 => conv_std_logic_vector(7, 8),
3239 => conv_std_logic_vector(7, 8),
3240 => conv_std_logic_vector(7, 8),
3241 => conv_std_logic_vector(7, 8),
3242 => conv_std_logic_vector(7, 8),
3243 => conv_std_logic_vector(8, 8),
3244 => conv_std_logic_vector(8, 8),
3245 => conv_std_logic_vector(8, 8),
3246 => conv_std_logic_vector(8, 8),
3247 => conv_std_logic_vector(8, 8),
3248 => conv_std_logic_vector(8, 8),
3249 => conv_std_logic_vector(8, 8),
3250 => conv_std_logic_vector(8, 8),
3251 => conv_std_logic_vector(8, 8),
3252 => conv_std_logic_vector(8, 8),
3253 => conv_std_logic_vector(8, 8),
3254 => conv_std_logic_vector(8, 8),
3255 => conv_std_logic_vector(8, 8),
3256 => conv_std_logic_vector(8, 8),
3257 => conv_std_logic_vector(8, 8),
3258 => conv_std_logic_vector(8, 8),
3259 => conv_std_logic_vector(8, 8),
3260 => conv_std_logic_vector(8, 8),
3261 => conv_std_logic_vector(8, 8),
3262 => conv_std_logic_vector(8, 8),
3263 => conv_std_logic_vector(8, 8),
3264 => conv_std_logic_vector(9, 8),
3265 => conv_std_logic_vector(9, 8),
3266 => conv_std_logic_vector(9, 8),
3267 => conv_std_logic_vector(9, 8),
3268 => conv_std_logic_vector(9, 8),
3269 => conv_std_logic_vector(9, 8),
3270 => conv_std_logic_vector(9, 8),
3271 => conv_std_logic_vector(9, 8),
3272 => conv_std_logic_vector(9, 8),
3273 => conv_std_logic_vector(9, 8),
3274 => conv_std_logic_vector(9, 8),
3275 => conv_std_logic_vector(9, 8),
3276 => conv_std_logic_vector(9, 8),
3277 => conv_std_logic_vector(9, 8),
3278 => conv_std_logic_vector(9, 8),
3279 => conv_std_logic_vector(9, 8),
3280 => conv_std_logic_vector(9, 8),
3281 => conv_std_logic_vector(9, 8),
3282 => conv_std_logic_vector(9, 8),
3283 => conv_std_logic_vector(9, 8),
3284 => conv_std_logic_vector(9, 8),
3285 => conv_std_logic_vector(9, 8),
3286 => conv_std_logic_vector(10, 8),
3287 => conv_std_logic_vector(10, 8),
3288 => conv_std_logic_vector(10, 8),
3289 => conv_std_logic_vector(10, 8),
3290 => conv_std_logic_vector(10, 8),
3291 => conv_std_logic_vector(10, 8),
3292 => conv_std_logic_vector(10, 8),
3293 => conv_std_logic_vector(10, 8),
3294 => conv_std_logic_vector(10, 8),
3295 => conv_std_logic_vector(10, 8),
3296 => conv_std_logic_vector(10, 8),
3297 => conv_std_logic_vector(10, 8),
3298 => conv_std_logic_vector(10, 8),
3299 => conv_std_logic_vector(10, 8),
3300 => conv_std_logic_vector(10, 8),
3301 => conv_std_logic_vector(10, 8),
3302 => conv_std_logic_vector(10, 8),
3303 => conv_std_logic_vector(10, 8),
3304 => conv_std_logic_vector(10, 8),
3305 => conv_std_logic_vector(10, 8),
3306 => conv_std_logic_vector(10, 8),
3307 => conv_std_logic_vector(11, 8),
3308 => conv_std_logic_vector(11, 8),
3309 => conv_std_logic_vector(11, 8),
3310 => conv_std_logic_vector(11, 8),
3311 => conv_std_logic_vector(11, 8),
3312 => conv_std_logic_vector(11, 8),
3313 => conv_std_logic_vector(11, 8),
3314 => conv_std_logic_vector(11, 8),
3315 => conv_std_logic_vector(11, 8),
3316 => conv_std_logic_vector(11, 8),
3317 => conv_std_logic_vector(11, 8),
3318 => conv_std_logic_vector(11, 8),
3319 => conv_std_logic_vector(11, 8),
3320 => conv_std_logic_vector(11, 8),
3321 => conv_std_logic_vector(11, 8),
3322 => conv_std_logic_vector(11, 8),
3323 => conv_std_logic_vector(11, 8),
3324 => conv_std_logic_vector(11, 8),
3325 => conv_std_logic_vector(11, 8),
3326 => conv_std_logic_vector(11, 8),
3327 => conv_std_logic_vector(11, 8),
3328 => conv_std_logic_vector(0, 8),
3329 => conv_std_logic_vector(0, 8),
3330 => conv_std_logic_vector(0, 8),
3331 => conv_std_logic_vector(0, 8),
3332 => conv_std_logic_vector(0, 8),
3333 => conv_std_logic_vector(0, 8),
3334 => conv_std_logic_vector(0, 8),
3335 => conv_std_logic_vector(0, 8),
3336 => conv_std_logic_vector(0, 8),
3337 => conv_std_logic_vector(0, 8),
3338 => conv_std_logic_vector(0, 8),
3339 => conv_std_logic_vector(0, 8),
3340 => conv_std_logic_vector(0, 8),
3341 => conv_std_logic_vector(0, 8),
3342 => conv_std_logic_vector(0, 8),
3343 => conv_std_logic_vector(0, 8),
3344 => conv_std_logic_vector(0, 8),
3345 => conv_std_logic_vector(0, 8),
3346 => conv_std_logic_vector(0, 8),
3347 => conv_std_logic_vector(0, 8),
3348 => conv_std_logic_vector(1, 8),
3349 => conv_std_logic_vector(1, 8),
3350 => conv_std_logic_vector(1, 8),
3351 => conv_std_logic_vector(1, 8),
3352 => conv_std_logic_vector(1, 8),
3353 => conv_std_logic_vector(1, 8),
3354 => conv_std_logic_vector(1, 8),
3355 => conv_std_logic_vector(1, 8),
3356 => conv_std_logic_vector(1, 8),
3357 => conv_std_logic_vector(1, 8),
3358 => conv_std_logic_vector(1, 8),
3359 => conv_std_logic_vector(1, 8),
3360 => conv_std_logic_vector(1, 8),
3361 => conv_std_logic_vector(1, 8),
3362 => conv_std_logic_vector(1, 8),
3363 => conv_std_logic_vector(1, 8),
3364 => conv_std_logic_vector(1, 8),
3365 => conv_std_logic_vector(1, 8),
3366 => conv_std_logic_vector(1, 8),
3367 => conv_std_logic_vector(1, 8),
3368 => conv_std_logic_vector(2, 8),
3369 => conv_std_logic_vector(2, 8),
3370 => conv_std_logic_vector(2, 8),
3371 => conv_std_logic_vector(2, 8),
3372 => conv_std_logic_vector(2, 8),
3373 => conv_std_logic_vector(2, 8),
3374 => conv_std_logic_vector(2, 8),
3375 => conv_std_logic_vector(2, 8),
3376 => conv_std_logic_vector(2, 8),
3377 => conv_std_logic_vector(2, 8),
3378 => conv_std_logic_vector(2, 8),
3379 => conv_std_logic_vector(2, 8),
3380 => conv_std_logic_vector(2, 8),
3381 => conv_std_logic_vector(2, 8),
3382 => conv_std_logic_vector(2, 8),
3383 => conv_std_logic_vector(2, 8),
3384 => conv_std_logic_vector(2, 8),
3385 => conv_std_logic_vector(2, 8),
3386 => conv_std_logic_vector(2, 8),
3387 => conv_std_logic_vector(2, 8),
3388 => conv_std_logic_vector(3, 8),
3389 => conv_std_logic_vector(3, 8),
3390 => conv_std_logic_vector(3, 8),
3391 => conv_std_logic_vector(3, 8),
3392 => conv_std_logic_vector(3, 8),
3393 => conv_std_logic_vector(3, 8),
3394 => conv_std_logic_vector(3, 8),
3395 => conv_std_logic_vector(3, 8),
3396 => conv_std_logic_vector(3, 8),
3397 => conv_std_logic_vector(3, 8),
3398 => conv_std_logic_vector(3, 8),
3399 => conv_std_logic_vector(3, 8),
3400 => conv_std_logic_vector(3, 8),
3401 => conv_std_logic_vector(3, 8),
3402 => conv_std_logic_vector(3, 8),
3403 => conv_std_logic_vector(3, 8),
3404 => conv_std_logic_vector(3, 8),
3405 => conv_std_logic_vector(3, 8),
3406 => conv_std_logic_vector(3, 8),
3407 => conv_std_logic_vector(4, 8),
3408 => conv_std_logic_vector(4, 8),
3409 => conv_std_logic_vector(4, 8),
3410 => conv_std_logic_vector(4, 8),
3411 => conv_std_logic_vector(4, 8),
3412 => conv_std_logic_vector(4, 8),
3413 => conv_std_logic_vector(4, 8),
3414 => conv_std_logic_vector(4, 8),
3415 => conv_std_logic_vector(4, 8),
3416 => conv_std_logic_vector(4, 8),
3417 => conv_std_logic_vector(4, 8),
3418 => conv_std_logic_vector(4, 8),
3419 => conv_std_logic_vector(4, 8),
3420 => conv_std_logic_vector(4, 8),
3421 => conv_std_logic_vector(4, 8),
3422 => conv_std_logic_vector(4, 8),
3423 => conv_std_logic_vector(4, 8),
3424 => conv_std_logic_vector(4, 8),
3425 => conv_std_logic_vector(4, 8),
3426 => conv_std_logic_vector(4, 8),
3427 => conv_std_logic_vector(5, 8),
3428 => conv_std_logic_vector(5, 8),
3429 => conv_std_logic_vector(5, 8),
3430 => conv_std_logic_vector(5, 8),
3431 => conv_std_logic_vector(5, 8),
3432 => conv_std_logic_vector(5, 8),
3433 => conv_std_logic_vector(5, 8),
3434 => conv_std_logic_vector(5, 8),
3435 => conv_std_logic_vector(5, 8),
3436 => conv_std_logic_vector(5, 8),
3437 => conv_std_logic_vector(5, 8),
3438 => conv_std_logic_vector(5, 8),
3439 => conv_std_logic_vector(5, 8),
3440 => conv_std_logic_vector(5, 8),
3441 => conv_std_logic_vector(5, 8),
3442 => conv_std_logic_vector(5, 8),
3443 => conv_std_logic_vector(5, 8),
3444 => conv_std_logic_vector(5, 8),
3445 => conv_std_logic_vector(5, 8),
3446 => conv_std_logic_vector(5, 8),
3447 => conv_std_logic_vector(6, 8),
3448 => conv_std_logic_vector(6, 8),
3449 => conv_std_logic_vector(6, 8),
3450 => conv_std_logic_vector(6, 8),
3451 => conv_std_logic_vector(6, 8),
3452 => conv_std_logic_vector(6, 8),
3453 => conv_std_logic_vector(6, 8),
3454 => conv_std_logic_vector(6, 8),
3455 => conv_std_logic_vector(6, 8),
3456 => conv_std_logic_vector(6, 8),
3457 => conv_std_logic_vector(6, 8),
3458 => conv_std_logic_vector(6, 8),
3459 => conv_std_logic_vector(6, 8),
3460 => conv_std_logic_vector(6, 8),
3461 => conv_std_logic_vector(6, 8),
3462 => conv_std_logic_vector(6, 8),
3463 => conv_std_logic_vector(6, 8),
3464 => conv_std_logic_vector(6, 8),
3465 => conv_std_logic_vector(6, 8),
3466 => conv_std_logic_vector(7, 8),
3467 => conv_std_logic_vector(7, 8),
3468 => conv_std_logic_vector(7, 8),
3469 => conv_std_logic_vector(7, 8),
3470 => conv_std_logic_vector(7, 8),
3471 => conv_std_logic_vector(7, 8),
3472 => conv_std_logic_vector(7, 8),
3473 => conv_std_logic_vector(7, 8),
3474 => conv_std_logic_vector(7, 8),
3475 => conv_std_logic_vector(7, 8),
3476 => conv_std_logic_vector(7, 8),
3477 => conv_std_logic_vector(7, 8),
3478 => conv_std_logic_vector(7, 8),
3479 => conv_std_logic_vector(7, 8),
3480 => conv_std_logic_vector(7, 8),
3481 => conv_std_logic_vector(7, 8),
3482 => conv_std_logic_vector(7, 8),
3483 => conv_std_logic_vector(7, 8),
3484 => conv_std_logic_vector(7, 8),
3485 => conv_std_logic_vector(7, 8),
3486 => conv_std_logic_vector(8, 8),
3487 => conv_std_logic_vector(8, 8),
3488 => conv_std_logic_vector(8, 8),
3489 => conv_std_logic_vector(8, 8),
3490 => conv_std_logic_vector(8, 8),
3491 => conv_std_logic_vector(8, 8),
3492 => conv_std_logic_vector(8, 8),
3493 => conv_std_logic_vector(8, 8),
3494 => conv_std_logic_vector(8, 8),
3495 => conv_std_logic_vector(8, 8),
3496 => conv_std_logic_vector(8, 8),
3497 => conv_std_logic_vector(8, 8),
3498 => conv_std_logic_vector(8, 8),
3499 => conv_std_logic_vector(8, 8),
3500 => conv_std_logic_vector(8, 8),
3501 => conv_std_logic_vector(8, 8),
3502 => conv_std_logic_vector(8, 8),
3503 => conv_std_logic_vector(8, 8),
3504 => conv_std_logic_vector(8, 8),
3505 => conv_std_logic_vector(8, 8),
3506 => conv_std_logic_vector(9, 8),
3507 => conv_std_logic_vector(9, 8),
3508 => conv_std_logic_vector(9, 8),
3509 => conv_std_logic_vector(9, 8),
3510 => conv_std_logic_vector(9, 8),
3511 => conv_std_logic_vector(9, 8),
3512 => conv_std_logic_vector(9, 8),
3513 => conv_std_logic_vector(9, 8),
3514 => conv_std_logic_vector(9, 8),
3515 => conv_std_logic_vector(9, 8),
3516 => conv_std_logic_vector(9, 8),
3517 => conv_std_logic_vector(9, 8),
3518 => conv_std_logic_vector(9, 8),
3519 => conv_std_logic_vector(9, 8),
3520 => conv_std_logic_vector(9, 8),
3521 => conv_std_logic_vector(9, 8),
3522 => conv_std_logic_vector(9, 8),
3523 => conv_std_logic_vector(9, 8),
3524 => conv_std_logic_vector(9, 8),
3525 => conv_std_logic_vector(10, 8),
3526 => conv_std_logic_vector(10, 8),
3527 => conv_std_logic_vector(10, 8),
3528 => conv_std_logic_vector(10, 8),
3529 => conv_std_logic_vector(10, 8),
3530 => conv_std_logic_vector(10, 8),
3531 => conv_std_logic_vector(10, 8),
3532 => conv_std_logic_vector(10, 8),
3533 => conv_std_logic_vector(10, 8),
3534 => conv_std_logic_vector(10, 8),
3535 => conv_std_logic_vector(10, 8),
3536 => conv_std_logic_vector(10, 8),
3537 => conv_std_logic_vector(10, 8),
3538 => conv_std_logic_vector(10, 8),
3539 => conv_std_logic_vector(10, 8),
3540 => conv_std_logic_vector(10, 8),
3541 => conv_std_logic_vector(10, 8),
3542 => conv_std_logic_vector(10, 8),
3543 => conv_std_logic_vector(10, 8),
3544 => conv_std_logic_vector(10, 8),
3545 => conv_std_logic_vector(11, 8),
3546 => conv_std_logic_vector(11, 8),
3547 => conv_std_logic_vector(11, 8),
3548 => conv_std_logic_vector(11, 8),
3549 => conv_std_logic_vector(11, 8),
3550 => conv_std_logic_vector(11, 8),
3551 => conv_std_logic_vector(11, 8),
3552 => conv_std_logic_vector(11, 8),
3553 => conv_std_logic_vector(11, 8),
3554 => conv_std_logic_vector(11, 8),
3555 => conv_std_logic_vector(11, 8),
3556 => conv_std_logic_vector(11, 8),
3557 => conv_std_logic_vector(11, 8),
3558 => conv_std_logic_vector(11, 8),
3559 => conv_std_logic_vector(11, 8),
3560 => conv_std_logic_vector(11, 8),
3561 => conv_std_logic_vector(11, 8),
3562 => conv_std_logic_vector(11, 8),
3563 => conv_std_logic_vector(11, 8),
3564 => conv_std_logic_vector(11, 8),
3565 => conv_std_logic_vector(12, 8),
3566 => conv_std_logic_vector(12, 8),
3567 => conv_std_logic_vector(12, 8),
3568 => conv_std_logic_vector(12, 8),
3569 => conv_std_logic_vector(12, 8),
3570 => conv_std_logic_vector(12, 8),
3571 => conv_std_logic_vector(12, 8),
3572 => conv_std_logic_vector(12, 8),
3573 => conv_std_logic_vector(12, 8),
3574 => conv_std_logic_vector(12, 8),
3575 => conv_std_logic_vector(12, 8),
3576 => conv_std_logic_vector(12, 8),
3577 => conv_std_logic_vector(12, 8),
3578 => conv_std_logic_vector(12, 8),
3579 => conv_std_logic_vector(12, 8),
3580 => conv_std_logic_vector(12, 8),
3581 => conv_std_logic_vector(12, 8),
3582 => conv_std_logic_vector(12, 8),
3583 => conv_std_logic_vector(12, 8),
3584 => conv_std_logic_vector(0, 8),
3585 => conv_std_logic_vector(0, 8),
3586 => conv_std_logic_vector(0, 8),
3587 => conv_std_logic_vector(0, 8),
3588 => conv_std_logic_vector(0, 8),
3589 => conv_std_logic_vector(0, 8),
3590 => conv_std_logic_vector(0, 8),
3591 => conv_std_logic_vector(0, 8),
3592 => conv_std_logic_vector(0, 8),
3593 => conv_std_logic_vector(0, 8),
3594 => conv_std_logic_vector(0, 8),
3595 => conv_std_logic_vector(0, 8),
3596 => conv_std_logic_vector(0, 8),
3597 => conv_std_logic_vector(0, 8),
3598 => conv_std_logic_vector(0, 8),
3599 => conv_std_logic_vector(0, 8),
3600 => conv_std_logic_vector(0, 8),
3601 => conv_std_logic_vector(0, 8),
3602 => conv_std_logic_vector(0, 8),
3603 => conv_std_logic_vector(1, 8),
3604 => conv_std_logic_vector(1, 8),
3605 => conv_std_logic_vector(1, 8),
3606 => conv_std_logic_vector(1, 8),
3607 => conv_std_logic_vector(1, 8),
3608 => conv_std_logic_vector(1, 8),
3609 => conv_std_logic_vector(1, 8),
3610 => conv_std_logic_vector(1, 8),
3611 => conv_std_logic_vector(1, 8),
3612 => conv_std_logic_vector(1, 8),
3613 => conv_std_logic_vector(1, 8),
3614 => conv_std_logic_vector(1, 8),
3615 => conv_std_logic_vector(1, 8),
3616 => conv_std_logic_vector(1, 8),
3617 => conv_std_logic_vector(1, 8),
3618 => conv_std_logic_vector(1, 8),
3619 => conv_std_logic_vector(1, 8),
3620 => conv_std_logic_vector(1, 8),
3621 => conv_std_logic_vector(2, 8),
3622 => conv_std_logic_vector(2, 8),
3623 => conv_std_logic_vector(2, 8),
3624 => conv_std_logic_vector(2, 8),
3625 => conv_std_logic_vector(2, 8),
3626 => conv_std_logic_vector(2, 8),
3627 => conv_std_logic_vector(2, 8),
3628 => conv_std_logic_vector(2, 8),
3629 => conv_std_logic_vector(2, 8),
3630 => conv_std_logic_vector(2, 8),
3631 => conv_std_logic_vector(2, 8),
3632 => conv_std_logic_vector(2, 8),
3633 => conv_std_logic_vector(2, 8),
3634 => conv_std_logic_vector(2, 8),
3635 => conv_std_logic_vector(2, 8),
3636 => conv_std_logic_vector(2, 8),
3637 => conv_std_logic_vector(2, 8),
3638 => conv_std_logic_vector(2, 8),
3639 => conv_std_logic_vector(3, 8),
3640 => conv_std_logic_vector(3, 8),
3641 => conv_std_logic_vector(3, 8),
3642 => conv_std_logic_vector(3, 8),
3643 => conv_std_logic_vector(3, 8),
3644 => conv_std_logic_vector(3, 8),
3645 => conv_std_logic_vector(3, 8),
3646 => conv_std_logic_vector(3, 8),
3647 => conv_std_logic_vector(3, 8),
3648 => conv_std_logic_vector(3, 8),
3649 => conv_std_logic_vector(3, 8),
3650 => conv_std_logic_vector(3, 8),
3651 => conv_std_logic_vector(3, 8),
3652 => conv_std_logic_vector(3, 8),
3653 => conv_std_logic_vector(3, 8),
3654 => conv_std_logic_vector(3, 8),
3655 => conv_std_logic_vector(3, 8),
3656 => conv_std_logic_vector(3, 8),
3657 => conv_std_logic_vector(3, 8),
3658 => conv_std_logic_vector(4, 8),
3659 => conv_std_logic_vector(4, 8),
3660 => conv_std_logic_vector(4, 8),
3661 => conv_std_logic_vector(4, 8),
3662 => conv_std_logic_vector(4, 8),
3663 => conv_std_logic_vector(4, 8),
3664 => conv_std_logic_vector(4, 8),
3665 => conv_std_logic_vector(4, 8),
3666 => conv_std_logic_vector(4, 8),
3667 => conv_std_logic_vector(4, 8),
3668 => conv_std_logic_vector(4, 8),
3669 => conv_std_logic_vector(4, 8),
3670 => conv_std_logic_vector(4, 8),
3671 => conv_std_logic_vector(4, 8),
3672 => conv_std_logic_vector(4, 8),
3673 => conv_std_logic_vector(4, 8),
3674 => conv_std_logic_vector(4, 8),
3675 => conv_std_logic_vector(4, 8),
3676 => conv_std_logic_vector(5, 8),
3677 => conv_std_logic_vector(5, 8),
3678 => conv_std_logic_vector(5, 8),
3679 => conv_std_logic_vector(5, 8),
3680 => conv_std_logic_vector(5, 8),
3681 => conv_std_logic_vector(5, 8),
3682 => conv_std_logic_vector(5, 8),
3683 => conv_std_logic_vector(5, 8),
3684 => conv_std_logic_vector(5, 8),
3685 => conv_std_logic_vector(5, 8),
3686 => conv_std_logic_vector(5, 8),
3687 => conv_std_logic_vector(5, 8),
3688 => conv_std_logic_vector(5, 8),
3689 => conv_std_logic_vector(5, 8),
3690 => conv_std_logic_vector(5, 8),
3691 => conv_std_logic_vector(5, 8),
3692 => conv_std_logic_vector(5, 8),
3693 => conv_std_logic_vector(5, 8),
3694 => conv_std_logic_vector(6, 8),
3695 => conv_std_logic_vector(6, 8),
3696 => conv_std_logic_vector(6, 8),
3697 => conv_std_logic_vector(6, 8),
3698 => conv_std_logic_vector(6, 8),
3699 => conv_std_logic_vector(6, 8),
3700 => conv_std_logic_vector(6, 8),
3701 => conv_std_logic_vector(6, 8),
3702 => conv_std_logic_vector(6, 8),
3703 => conv_std_logic_vector(6, 8),
3704 => conv_std_logic_vector(6, 8),
3705 => conv_std_logic_vector(6, 8),
3706 => conv_std_logic_vector(6, 8),
3707 => conv_std_logic_vector(6, 8),
3708 => conv_std_logic_vector(6, 8),
3709 => conv_std_logic_vector(6, 8),
3710 => conv_std_logic_vector(6, 8),
3711 => conv_std_logic_vector(6, 8),
3712 => conv_std_logic_vector(7, 8),
3713 => conv_std_logic_vector(7, 8),
3714 => conv_std_logic_vector(7, 8),
3715 => conv_std_logic_vector(7, 8),
3716 => conv_std_logic_vector(7, 8),
3717 => conv_std_logic_vector(7, 8),
3718 => conv_std_logic_vector(7, 8),
3719 => conv_std_logic_vector(7, 8),
3720 => conv_std_logic_vector(7, 8),
3721 => conv_std_logic_vector(7, 8),
3722 => conv_std_logic_vector(7, 8),
3723 => conv_std_logic_vector(7, 8),
3724 => conv_std_logic_vector(7, 8),
3725 => conv_std_logic_vector(7, 8),
3726 => conv_std_logic_vector(7, 8),
3727 => conv_std_logic_vector(7, 8),
3728 => conv_std_logic_vector(7, 8),
3729 => conv_std_logic_vector(7, 8),
3730 => conv_std_logic_vector(7, 8),
3731 => conv_std_logic_vector(8, 8),
3732 => conv_std_logic_vector(8, 8),
3733 => conv_std_logic_vector(8, 8),
3734 => conv_std_logic_vector(8, 8),
3735 => conv_std_logic_vector(8, 8),
3736 => conv_std_logic_vector(8, 8),
3737 => conv_std_logic_vector(8, 8),
3738 => conv_std_logic_vector(8, 8),
3739 => conv_std_logic_vector(8, 8),
3740 => conv_std_logic_vector(8, 8),
3741 => conv_std_logic_vector(8, 8),
3742 => conv_std_logic_vector(8, 8),
3743 => conv_std_logic_vector(8, 8),
3744 => conv_std_logic_vector(8, 8),
3745 => conv_std_logic_vector(8, 8),
3746 => conv_std_logic_vector(8, 8),
3747 => conv_std_logic_vector(8, 8),
3748 => conv_std_logic_vector(8, 8),
3749 => conv_std_logic_vector(9, 8),
3750 => conv_std_logic_vector(9, 8),
3751 => conv_std_logic_vector(9, 8),
3752 => conv_std_logic_vector(9, 8),
3753 => conv_std_logic_vector(9, 8),
3754 => conv_std_logic_vector(9, 8),
3755 => conv_std_logic_vector(9, 8),
3756 => conv_std_logic_vector(9, 8),
3757 => conv_std_logic_vector(9, 8),
3758 => conv_std_logic_vector(9, 8),
3759 => conv_std_logic_vector(9, 8),
3760 => conv_std_logic_vector(9, 8),
3761 => conv_std_logic_vector(9, 8),
3762 => conv_std_logic_vector(9, 8),
3763 => conv_std_logic_vector(9, 8),
3764 => conv_std_logic_vector(9, 8),
3765 => conv_std_logic_vector(9, 8),
3766 => conv_std_logic_vector(9, 8),
3767 => conv_std_logic_vector(10, 8),
3768 => conv_std_logic_vector(10, 8),
3769 => conv_std_logic_vector(10, 8),
3770 => conv_std_logic_vector(10, 8),
3771 => conv_std_logic_vector(10, 8),
3772 => conv_std_logic_vector(10, 8),
3773 => conv_std_logic_vector(10, 8),
3774 => conv_std_logic_vector(10, 8),
3775 => conv_std_logic_vector(10, 8),
3776 => conv_std_logic_vector(10, 8),
3777 => conv_std_logic_vector(10, 8),
3778 => conv_std_logic_vector(10, 8),
3779 => conv_std_logic_vector(10, 8),
3780 => conv_std_logic_vector(10, 8),
3781 => conv_std_logic_vector(10, 8),
3782 => conv_std_logic_vector(10, 8),
3783 => conv_std_logic_vector(10, 8),
3784 => conv_std_logic_vector(10, 8),
3785 => conv_std_logic_vector(10, 8),
3786 => conv_std_logic_vector(11, 8),
3787 => conv_std_logic_vector(11, 8),
3788 => conv_std_logic_vector(11, 8),
3789 => conv_std_logic_vector(11, 8),
3790 => conv_std_logic_vector(11, 8),
3791 => conv_std_logic_vector(11, 8),
3792 => conv_std_logic_vector(11, 8),
3793 => conv_std_logic_vector(11, 8),
3794 => conv_std_logic_vector(11, 8),
3795 => conv_std_logic_vector(11, 8),
3796 => conv_std_logic_vector(11, 8),
3797 => conv_std_logic_vector(11, 8),
3798 => conv_std_logic_vector(11, 8),
3799 => conv_std_logic_vector(11, 8),
3800 => conv_std_logic_vector(11, 8),
3801 => conv_std_logic_vector(11, 8),
3802 => conv_std_logic_vector(11, 8),
3803 => conv_std_logic_vector(11, 8),
3804 => conv_std_logic_vector(12, 8),
3805 => conv_std_logic_vector(12, 8),
3806 => conv_std_logic_vector(12, 8),
3807 => conv_std_logic_vector(12, 8),
3808 => conv_std_logic_vector(12, 8),
3809 => conv_std_logic_vector(12, 8),
3810 => conv_std_logic_vector(12, 8),
3811 => conv_std_logic_vector(12, 8),
3812 => conv_std_logic_vector(12, 8),
3813 => conv_std_logic_vector(12, 8),
3814 => conv_std_logic_vector(12, 8),
3815 => conv_std_logic_vector(12, 8),
3816 => conv_std_logic_vector(12, 8),
3817 => conv_std_logic_vector(12, 8),
3818 => conv_std_logic_vector(12, 8),
3819 => conv_std_logic_vector(12, 8),
3820 => conv_std_logic_vector(12, 8),
3821 => conv_std_logic_vector(12, 8),
3822 => conv_std_logic_vector(13, 8),
3823 => conv_std_logic_vector(13, 8),
3824 => conv_std_logic_vector(13, 8),
3825 => conv_std_logic_vector(13, 8),
3826 => conv_std_logic_vector(13, 8),
3827 => conv_std_logic_vector(13, 8),
3828 => conv_std_logic_vector(13, 8),
3829 => conv_std_logic_vector(13, 8),
3830 => conv_std_logic_vector(13, 8),
3831 => conv_std_logic_vector(13, 8),
3832 => conv_std_logic_vector(13, 8),
3833 => conv_std_logic_vector(13, 8),
3834 => conv_std_logic_vector(13, 8),
3835 => conv_std_logic_vector(13, 8),
3836 => conv_std_logic_vector(13, 8),
3837 => conv_std_logic_vector(13, 8),
3838 => conv_std_logic_vector(13, 8),
3839 => conv_std_logic_vector(13, 8),
3840 => conv_std_logic_vector(0, 8),
3841 => conv_std_logic_vector(0, 8),
3842 => conv_std_logic_vector(0, 8),
3843 => conv_std_logic_vector(0, 8),
3844 => conv_std_logic_vector(0, 8),
3845 => conv_std_logic_vector(0, 8),
3846 => conv_std_logic_vector(0, 8),
3847 => conv_std_logic_vector(0, 8),
3848 => conv_std_logic_vector(0, 8),
3849 => conv_std_logic_vector(0, 8),
3850 => conv_std_logic_vector(0, 8),
3851 => conv_std_logic_vector(0, 8),
3852 => conv_std_logic_vector(0, 8),
3853 => conv_std_logic_vector(0, 8),
3854 => conv_std_logic_vector(0, 8),
3855 => conv_std_logic_vector(0, 8),
3856 => conv_std_logic_vector(0, 8),
3857 => conv_std_logic_vector(0, 8),
3858 => conv_std_logic_vector(1, 8),
3859 => conv_std_logic_vector(1, 8),
3860 => conv_std_logic_vector(1, 8),
3861 => conv_std_logic_vector(1, 8),
3862 => conv_std_logic_vector(1, 8),
3863 => conv_std_logic_vector(1, 8),
3864 => conv_std_logic_vector(1, 8),
3865 => conv_std_logic_vector(1, 8),
3866 => conv_std_logic_vector(1, 8),
3867 => conv_std_logic_vector(1, 8),
3868 => conv_std_logic_vector(1, 8),
3869 => conv_std_logic_vector(1, 8),
3870 => conv_std_logic_vector(1, 8),
3871 => conv_std_logic_vector(1, 8),
3872 => conv_std_logic_vector(1, 8),
3873 => conv_std_logic_vector(1, 8),
3874 => conv_std_logic_vector(1, 8),
3875 => conv_std_logic_vector(2, 8),
3876 => conv_std_logic_vector(2, 8),
3877 => conv_std_logic_vector(2, 8),
3878 => conv_std_logic_vector(2, 8),
3879 => conv_std_logic_vector(2, 8),
3880 => conv_std_logic_vector(2, 8),
3881 => conv_std_logic_vector(2, 8),
3882 => conv_std_logic_vector(2, 8),
3883 => conv_std_logic_vector(2, 8),
3884 => conv_std_logic_vector(2, 8),
3885 => conv_std_logic_vector(2, 8),
3886 => conv_std_logic_vector(2, 8),
3887 => conv_std_logic_vector(2, 8),
3888 => conv_std_logic_vector(2, 8),
3889 => conv_std_logic_vector(2, 8),
3890 => conv_std_logic_vector(2, 8),
3891 => conv_std_logic_vector(2, 8),
3892 => conv_std_logic_vector(3, 8),
3893 => conv_std_logic_vector(3, 8),
3894 => conv_std_logic_vector(3, 8),
3895 => conv_std_logic_vector(3, 8),
3896 => conv_std_logic_vector(3, 8),
3897 => conv_std_logic_vector(3, 8),
3898 => conv_std_logic_vector(3, 8),
3899 => conv_std_logic_vector(3, 8),
3900 => conv_std_logic_vector(3, 8),
3901 => conv_std_logic_vector(3, 8),
3902 => conv_std_logic_vector(3, 8),
3903 => conv_std_logic_vector(3, 8),
3904 => conv_std_logic_vector(3, 8),
3905 => conv_std_logic_vector(3, 8),
3906 => conv_std_logic_vector(3, 8),
3907 => conv_std_logic_vector(3, 8),
3908 => conv_std_logic_vector(3, 8),
3909 => conv_std_logic_vector(4, 8),
3910 => conv_std_logic_vector(4, 8),
3911 => conv_std_logic_vector(4, 8),
3912 => conv_std_logic_vector(4, 8),
3913 => conv_std_logic_vector(4, 8),
3914 => conv_std_logic_vector(4, 8),
3915 => conv_std_logic_vector(4, 8),
3916 => conv_std_logic_vector(4, 8),
3917 => conv_std_logic_vector(4, 8),
3918 => conv_std_logic_vector(4, 8),
3919 => conv_std_logic_vector(4, 8),
3920 => conv_std_logic_vector(4, 8),
3921 => conv_std_logic_vector(4, 8),
3922 => conv_std_logic_vector(4, 8),
3923 => conv_std_logic_vector(4, 8),
3924 => conv_std_logic_vector(4, 8),
3925 => conv_std_logic_vector(4, 8),
3926 => conv_std_logic_vector(5, 8),
3927 => conv_std_logic_vector(5, 8),
3928 => conv_std_logic_vector(5, 8),
3929 => conv_std_logic_vector(5, 8),
3930 => conv_std_logic_vector(5, 8),
3931 => conv_std_logic_vector(5, 8),
3932 => conv_std_logic_vector(5, 8),
3933 => conv_std_logic_vector(5, 8),
3934 => conv_std_logic_vector(5, 8),
3935 => conv_std_logic_vector(5, 8),
3936 => conv_std_logic_vector(5, 8),
3937 => conv_std_logic_vector(5, 8),
3938 => conv_std_logic_vector(5, 8),
3939 => conv_std_logic_vector(5, 8),
3940 => conv_std_logic_vector(5, 8),
3941 => conv_std_logic_vector(5, 8),
3942 => conv_std_logic_vector(5, 8),
3943 => conv_std_logic_vector(6, 8),
3944 => conv_std_logic_vector(6, 8),
3945 => conv_std_logic_vector(6, 8),
3946 => conv_std_logic_vector(6, 8),
3947 => conv_std_logic_vector(6, 8),
3948 => conv_std_logic_vector(6, 8),
3949 => conv_std_logic_vector(6, 8),
3950 => conv_std_logic_vector(6, 8),
3951 => conv_std_logic_vector(6, 8),
3952 => conv_std_logic_vector(6, 8),
3953 => conv_std_logic_vector(6, 8),
3954 => conv_std_logic_vector(6, 8),
3955 => conv_std_logic_vector(6, 8),
3956 => conv_std_logic_vector(6, 8),
3957 => conv_std_logic_vector(6, 8),
3958 => conv_std_logic_vector(6, 8),
3959 => conv_std_logic_vector(6, 8),
3960 => conv_std_logic_vector(7, 8),
3961 => conv_std_logic_vector(7, 8),
3962 => conv_std_logic_vector(7, 8),
3963 => conv_std_logic_vector(7, 8),
3964 => conv_std_logic_vector(7, 8),
3965 => conv_std_logic_vector(7, 8),
3966 => conv_std_logic_vector(7, 8),
3967 => conv_std_logic_vector(7, 8),
3968 => conv_std_logic_vector(7, 8),
3969 => conv_std_logic_vector(7, 8),
3970 => conv_std_logic_vector(7, 8),
3971 => conv_std_logic_vector(7, 8),
3972 => conv_std_logic_vector(7, 8),
3973 => conv_std_logic_vector(7, 8),
3974 => conv_std_logic_vector(7, 8),
3975 => conv_std_logic_vector(7, 8),
3976 => conv_std_logic_vector(7, 8),
3977 => conv_std_logic_vector(8, 8),
3978 => conv_std_logic_vector(8, 8),
3979 => conv_std_logic_vector(8, 8),
3980 => conv_std_logic_vector(8, 8),
3981 => conv_std_logic_vector(8, 8),
3982 => conv_std_logic_vector(8, 8),
3983 => conv_std_logic_vector(8, 8),
3984 => conv_std_logic_vector(8, 8),
3985 => conv_std_logic_vector(8, 8),
3986 => conv_std_logic_vector(8, 8),
3987 => conv_std_logic_vector(8, 8),
3988 => conv_std_logic_vector(8, 8),
3989 => conv_std_logic_vector(8, 8),
3990 => conv_std_logic_vector(8, 8),
3991 => conv_std_logic_vector(8, 8),
3992 => conv_std_logic_vector(8, 8),
3993 => conv_std_logic_vector(8, 8),
3994 => conv_std_logic_vector(9, 8),
3995 => conv_std_logic_vector(9, 8),
3996 => conv_std_logic_vector(9, 8),
3997 => conv_std_logic_vector(9, 8),
3998 => conv_std_logic_vector(9, 8),
3999 => conv_std_logic_vector(9, 8),
4000 => conv_std_logic_vector(9, 8),
4001 => conv_std_logic_vector(9, 8),
4002 => conv_std_logic_vector(9, 8),
4003 => conv_std_logic_vector(9, 8),
4004 => conv_std_logic_vector(9, 8),
4005 => conv_std_logic_vector(9, 8),
4006 => conv_std_logic_vector(9, 8),
4007 => conv_std_logic_vector(9, 8),
4008 => conv_std_logic_vector(9, 8),
4009 => conv_std_logic_vector(9, 8),
4010 => conv_std_logic_vector(9, 8),
4011 => conv_std_logic_vector(10, 8),
4012 => conv_std_logic_vector(10, 8),
4013 => conv_std_logic_vector(10, 8),
4014 => conv_std_logic_vector(10, 8),
4015 => conv_std_logic_vector(10, 8),
4016 => conv_std_logic_vector(10, 8),
4017 => conv_std_logic_vector(10, 8),
4018 => conv_std_logic_vector(10, 8),
4019 => conv_std_logic_vector(10, 8),
4020 => conv_std_logic_vector(10, 8),
4021 => conv_std_logic_vector(10, 8),
4022 => conv_std_logic_vector(10, 8),
4023 => conv_std_logic_vector(10, 8),
4024 => conv_std_logic_vector(10, 8),
4025 => conv_std_logic_vector(10, 8),
4026 => conv_std_logic_vector(10, 8),
4027 => conv_std_logic_vector(10, 8),
4028 => conv_std_logic_vector(11, 8),
4029 => conv_std_logic_vector(11, 8),
4030 => conv_std_logic_vector(11, 8),
4031 => conv_std_logic_vector(11, 8),
4032 => conv_std_logic_vector(11, 8),
4033 => conv_std_logic_vector(11, 8),
4034 => conv_std_logic_vector(11, 8),
4035 => conv_std_logic_vector(11, 8),
4036 => conv_std_logic_vector(11, 8),
4037 => conv_std_logic_vector(11, 8),
4038 => conv_std_logic_vector(11, 8),
4039 => conv_std_logic_vector(11, 8),
4040 => conv_std_logic_vector(11, 8),
4041 => conv_std_logic_vector(11, 8),
4042 => conv_std_logic_vector(11, 8),
4043 => conv_std_logic_vector(11, 8),
4044 => conv_std_logic_vector(11, 8),
4045 => conv_std_logic_vector(12, 8),
4046 => conv_std_logic_vector(12, 8),
4047 => conv_std_logic_vector(12, 8),
4048 => conv_std_logic_vector(12, 8),
4049 => conv_std_logic_vector(12, 8),
4050 => conv_std_logic_vector(12, 8),
4051 => conv_std_logic_vector(12, 8),
4052 => conv_std_logic_vector(12, 8),
4053 => conv_std_logic_vector(12, 8),
4054 => conv_std_logic_vector(12, 8),
4055 => conv_std_logic_vector(12, 8),
4056 => conv_std_logic_vector(12, 8),
4057 => conv_std_logic_vector(12, 8),
4058 => conv_std_logic_vector(12, 8),
4059 => conv_std_logic_vector(12, 8),
4060 => conv_std_logic_vector(12, 8),
4061 => conv_std_logic_vector(12, 8),
4062 => conv_std_logic_vector(13, 8),
4063 => conv_std_logic_vector(13, 8),
4064 => conv_std_logic_vector(13, 8),
4065 => conv_std_logic_vector(13, 8),
4066 => conv_std_logic_vector(13, 8),
4067 => conv_std_logic_vector(13, 8),
4068 => conv_std_logic_vector(13, 8),
4069 => conv_std_logic_vector(13, 8),
4070 => conv_std_logic_vector(13, 8),
4071 => conv_std_logic_vector(13, 8),
4072 => conv_std_logic_vector(13, 8),
4073 => conv_std_logic_vector(13, 8),
4074 => conv_std_logic_vector(13, 8),
4075 => conv_std_logic_vector(13, 8),
4076 => conv_std_logic_vector(13, 8),
4077 => conv_std_logic_vector(13, 8),
4078 => conv_std_logic_vector(13, 8),
4079 => conv_std_logic_vector(14, 8),
4080 => conv_std_logic_vector(14, 8),
4081 => conv_std_logic_vector(14, 8),
4082 => conv_std_logic_vector(14, 8),
4083 => conv_std_logic_vector(14, 8),
4084 => conv_std_logic_vector(14, 8),
4085 => conv_std_logic_vector(14, 8),
4086 => conv_std_logic_vector(14, 8),
4087 => conv_std_logic_vector(14, 8),
4088 => conv_std_logic_vector(14, 8),
4089 => conv_std_logic_vector(14, 8),
4090 => conv_std_logic_vector(14, 8),
4091 => conv_std_logic_vector(14, 8),
4092 => conv_std_logic_vector(14, 8),
4093 => conv_std_logic_vector(14, 8),
4094 => conv_std_logic_vector(14, 8),
4095 => conv_std_logic_vector(14, 8),
4096 => conv_std_logic_vector(0, 8),
4097 => conv_std_logic_vector(0, 8),
4098 => conv_std_logic_vector(0, 8),
4099 => conv_std_logic_vector(0, 8),
4100 => conv_std_logic_vector(0, 8),
4101 => conv_std_logic_vector(0, 8),
4102 => conv_std_logic_vector(0, 8),
4103 => conv_std_logic_vector(0, 8),
4104 => conv_std_logic_vector(0, 8),
4105 => conv_std_logic_vector(0, 8),
4106 => conv_std_logic_vector(0, 8),
4107 => conv_std_logic_vector(0, 8),
4108 => conv_std_logic_vector(0, 8),
4109 => conv_std_logic_vector(0, 8),
4110 => conv_std_logic_vector(0, 8),
4111 => conv_std_logic_vector(0, 8),
4112 => conv_std_logic_vector(1, 8),
4113 => conv_std_logic_vector(1, 8),
4114 => conv_std_logic_vector(1, 8),
4115 => conv_std_logic_vector(1, 8),
4116 => conv_std_logic_vector(1, 8),
4117 => conv_std_logic_vector(1, 8),
4118 => conv_std_logic_vector(1, 8),
4119 => conv_std_logic_vector(1, 8),
4120 => conv_std_logic_vector(1, 8),
4121 => conv_std_logic_vector(1, 8),
4122 => conv_std_logic_vector(1, 8),
4123 => conv_std_logic_vector(1, 8),
4124 => conv_std_logic_vector(1, 8),
4125 => conv_std_logic_vector(1, 8),
4126 => conv_std_logic_vector(1, 8),
4127 => conv_std_logic_vector(1, 8),
4128 => conv_std_logic_vector(2, 8),
4129 => conv_std_logic_vector(2, 8),
4130 => conv_std_logic_vector(2, 8),
4131 => conv_std_logic_vector(2, 8),
4132 => conv_std_logic_vector(2, 8),
4133 => conv_std_logic_vector(2, 8),
4134 => conv_std_logic_vector(2, 8),
4135 => conv_std_logic_vector(2, 8),
4136 => conv_std_logic_vector(2, 8),
4137 => conv_std_logic_vector(2, 8),
4138 => conv_std_logic_vector(2, 8),
4139 => conv_std_logic_vector(2, 8),
4140 => conv_std_logic_vector(2, 8),
4141 => conv_std_logic_vector(2, 8),
4142 => conv_std_logic_vector(2, 8),
4143 => conv_std_logic_vector(2, 8),
4144 => conv_std_logic_vector(3, 8),
4145 => conv_std_logic_vector(3, 8),
4146 => conv_std_logic_vector(3, 8),
4147 => conv_std_logic_vector(3, 8),
4148 => conv_std_logic_vector(3, 8),
4149 => conv_std_logic_vector(3, 8),
4150 => conv_std_logic_vector(3, 8),
4151 => conv_std_logic_vector(3, 8),
4152 => conv_std_logic_vector(3, 8),
4153 => conv_std_logic_vector(3, 8),
4154 => conv_std_logic_vector(3, 8),
4155 => conv_std_logic_vector(3, 8),
4156 => conv_std_logic_vector(3, 8),
4157 => conv_std_logic_vector(3, 8),
4158 => conv_std_logic_vector(3, 8),
4159 => conv_std_logic_vector(3, 8),
4160 => conv_std_logic_vector(4, 8),
4161 => conv_std_logic_vector(4, 8),
4162 => conv_std_logic_vector(4, 8),
4163 => conv_std_logic_vector(4, 8),
4164 => conv_std_logic_vector(4, 8),
4165 => conv_std_logic_vector(4, 8),
4166 => conv_std_logic_vector(4, 8),
4167 => conv_std_logic_vector(4, 8),
4168 => conv_std_logic_vector(4, 8),
4169 => conv_std_logic_vector(4, 8),
4170 => conv_std_logic_vector(4, 8),
4171 => conv_std_logic_vector(4, 8),
4172 => conv_std_logic_vector(4, 8),
4173 => conv_std_logic_vector(4, 8),
4174 => conv_std_logic_vector(4, 8),
4175 => conv_std_logic_vector(4, 8),
4176 => conv_std_logic_vector(5, 8),
4177 => conv_std_logic_vector(5, 8),
4178 => conv_std_logic_vector(5, 8),
4179 => conv_std_logic_vector(5, 8),
4180 => conv_std_logic_vector(5, 8),
4181 => conv_std_logic_vector(5, 8),
4182 => conv_std_logic_vector(5, 8),
4183 => conv_std_logic_vector(5, 8),
4184 => conv_std_logic_vector(5, 8),
4185 => conv_std_logic_vector(5, 8),
4186 => conv_std_logic_vector(5, 8),
4187 => conv_std_logic_vector(5, 8),
4188 => conv_std_logic_vector(5, 8),
4189 => conv_std_logic_vector(5, 8),
4190 => conv_std_logic_vector(5, 8),
4191 => conv_std_logic_vector(5, 8),
4192 => conv_std_logic_vector(6, 8),
4193 => conv_std_logic_vector(6, 8),
4194 => conv_std_logic_vector(6, 8),
4195 => conv_std_logic_vector(6, 8),
4196 => conv_std_logic_vector(6, 8),
4197 => conv_std_logic_vector(6, 8),
4198 => conv_std_logic_vector(6, 8),
4199 => conv_std_logic_vector(6, 8),
4200 => conv_std_logic_vector(6, 8),
4201 => conv_std_logic_vector(6, 8),
4202 => conv_std_logic_vector(6, 8),
4203 => conv_std_logic_vector(6, 8),
4204 => conv_std_logic_vector(6, 8),
4205 => conv_std_logic_vector(6, 8),
4206 => conv_std_logic_vector(6, 8),
4207 => conv_std_logic_vector(6, 8),
4208 => conv_std_logic_vector(7, 8),
4209 => conv_std_logic_vector(7, 8),
4210 => conv_std_logic_vector(7, 8),
4211 => conv_std_logic_vector(7, 8),
4212 => conv_std_logic_vector(7, 8),
4213 => conv_std_logic_vector(7, 8),
4214 => conv_std_logic_vector(7, 8),
4215 => conv_std_logic_vector(7, 8),
4216 => conv_std_logic_vector(7, 8),
4217 => conv_std_logic_vector(7, 8),
4218 => conv_std_logic_vector(7, 8),
4219 => conv_std_logic_vector(7, 8),
4220 => conv_std_logic_vector(7, 8),
4221 => conv_std_logic_vector(7, 8),
4222 => conv_std_logic_vector(7, 8),
4223 => conv_std_logic_vector(7, 8),
4224 => conv_std_logic_vector(8, 8),
4225 => conv_std_logic_vector(8, 8),
4226 => conv_std_logic_vector(8, 8),
4227 => conv_std_logic_vector(8, 8),
4228 => conv_std_logic_vector(8, 8),
4229 => conv_std_logic_vector(8, 8),
4230 => conv_std_logic_vector(8, 8),
4231 => conv_std_logic_vector(8, 8),
4232 => conv_std_logic_vector(8, 8),
4233 => conv_std_logic_vector(8, 8),
4234 => conv_std_logic_vector(8, 8),
4235 => conv_std_logic_vector(8, 8),
4236 => conv_std_logic_vector(8, 8),
4237 => conv_std_logic_vector(8, 8),
4238 => conv_std_logic_vector(8, 8),
4239 => conv_std_logic_vector(8, 8),
4240 => conv_std_logic_vector(9, 8),
4241 => conv_std_logic_vector(9, 8),
4242 => conv_std_logic_vector(9, 8),
4243 => conv_std_logic_vector(9, 8),
4244 => conv_std_logic_vector(9, 8),
4245 => conv_std_logic_vector(9, 8),
4246 => conv_std_logic_vector(9, 8),
4247 => conv_std_logic_vector(9, 8),
4248 => conv_std_logic_vector(9, 8),
4249 => conv_std_logic_vector(9, 8),
4250 => conv_std_logic_vector(9, 8),
4251 => conv_std_logic_vector(9, 8),
4252 => conv_std_logic_vector(9, 8),
4253 => conv_std_logic_vector(9, 8),
4254 => conv_std_logic_vector(9, 8),
4255 => conv_std_logic_vector(9, 8),
4256 => conv_std_logic_vector(10, 8),
4257 => conv_std_logic_vector(10, 8),
4258 => conv_std_logic_vector(10, 8),
4259 => conv_std_logic_vector(10, 8),
4260 => conv_std_logic_vector(10, 8),
4261 => conv_std_logic_vector(10, 8),
4262 => conv_std_logic_vector(10, 8),
4263 => conv_std_logic_vector(10, 8),
4264 => conv_std_logic_vector(10, 8),
4265 => conv_std_logic_vector(10, 8),
4266 => conv_std_logic_vector(10, 8),
4267 => conv_std_logic_vector(10, 8),
4268 => conv_std_logic_vector(10, 8),
4269 => conv_std_logic_vector(10, 8),
4270 => conv_std_logic_vector(10, 8),
4271 => conv_std_logic_vector(10, 8),
4272 => conv_std_logic_vector(11, 8),
4273 => conv_std_logic_vector(11, 8),
4274 => conv_std_logic_vector(11, 8),
4275 => conv_std_logic_vector(11, 8),
4276 => conv_std_logic_vector(11, 8),
4277 => conv_std_logic_vector(11, 8),
4278 => conv_std_logic_vector(11, 8),
4279 => conv_std_logic_vector(11, 8),
4280 => conv_std_logic_vector(11, 8),
4281 => conv_std_logic_vector(11, 8),
4282 => conv_std_logic_vector(11, 8),
4283 => conv_std_logic_vector(11, 8),
4284 => conv_std_logic_vector(11, 8),
4285 => conv_std_logic_vector(11, 8),
4286 => conv_std_logic_vector(11, 8),
4287 => conv_std_logic_vector(11, 8),
4288 => conv_std_logic_vector(12, 8),
4289 => conv_std_logic_vector(12, 8),
4290 => conv_std_logic_vector(12, 8),
4291 => conv_std_logic_vector(12, 8),
4292 => conv_std_logic_vector(12, 8),
4293 => conv_std_logic_vector(12, 8),
4294 => conv_std_logic_vector(12, 8),
4295 => conv_std_logic_vector(12, 8),
4296 => conv_std_logic_vector(12, 8),
4297 => conv_std_logic_vector(12, 8),
4298 => conv_std_logic_vector(12, 8),
4299 => conv_std_logic_vector(12, 8),
4300 => conv_std_logic_vector(12, 8),
4301 => conv_std_logic_vector(12, 8),
4302 => conv_std_logic_vector(12, 8),
4303 => conv_std_logic_vector(12, 8),
4304 => conv_std_logic_vector(13, 8),
4305 => conv_std_logic_vector(13, 8),
4306 => conv_std_logic_vector(13, 8),
4307 => conv_std_logic_vector(13, 8),
4308 => conv_std_logic_vector(13, 8),
4309 => conv_std_logic_vector(13, 8),
4310 => conv_std_logic_vector(13, 8),
4311 => conv_std_logic_vector(13, 8),
4312 => conv_std_logic_vector(13, 8),
4313 => conv_std_logic_vector(13, 8),
4314 => conv_std_logic_vector(13, 8),
4315 => conv_std_logic_vector(13, 8),
4316 => conv_std_logic_vector(13, 8),
4317 => conv_std_logic_vector(13, 8),
4318 => conv_std_logic_vector(13, 8),
4319 => conv_std_logic_vector(13, 8),
4320 => conv_std_logic_vector(14, 8),
4321 => conv_std_logic_vector(14, 8),
4322 => conv_std_logic_vector(14, 8),
4323 => conv_std_logic_vector(14, 8),
4324 => conv_std_logic_vector(14, 8),
4325 => conv_std_logic_vector(14, 8),
4326 => conv_std_logic_vector(14, 8),
4327 => conv_std_logic_vector(14, 8),
4328 => conv_std_logic_vector(14, 8),
4329 => conv_std_logic_vector(14, 8),
4330 => conv_std_logic_vector(14, 8),
4331 => conv_std_logic_vector(14, 8),
4332 => conv_std_logic_vector(14, 8),
4333 => conv_std_logic_vector(14, 8),
4334 => conv_std_logic_vector(14, 8),
4335 => conv_std_logic_vector(14, 8),
4336 => conv_std_logic_vector(15, 8),
4337 => conv_std_logic_vector(15, 8),
4338 => conv_std_logic_vector(15, 8),
4339 => conv_std_logic_vector(15, 8),
4340 => conv_std_logic_vector(15, 8),
4341 => conv_std_logic_vector(15, 8),
4342 => conv_std_logic_vector(15, 8),
4343 => conv_std_logic_vector(15, 8),
4344 => conv_std_logic_vector(15, 8),
4345 => conv_std_logic_vector(15, 8),
4346 => conv_std_logic_vector(15, 8),
4347 => conv_std_logic_vector(15, 8),
4348 => conv_std_logic_vector(15, 8),
4349 => conv_std_logic_vector(15, 8),
4350 => conv_std_logic_vector(15, 8),
4351 => conv_std_logic_vector(15, 8),
4352 => conv_std_logic_vector(0, 8),
4353 => conv_std_logic_vector(0, 8),
4354 => conv_std_logic_vector(0, 8),
4355 => conv_std_logic_vector(0, 8),
4356 => conv_std_logic_vector(0, 8),
4357 => conv_std_logic_vector(0, 8),
4358 => conv_std_logic_vector(0, 8),
4359 => conv_std_logic_vector(0, 8),
4360 => conv_std_logic_vector(0, 8),
4361 => conv_std_logic_vector(0, 8),
4362 => conv_std_logic_vector(0, 8),
4363 => conv_std_logic_vector(0, 8),
4364 => conv_std_logic_vector(0, 8),
4365 => conv_std_logic_vector(0, 8),
4366 => conv_std_logic_vector(0, 8),
4367 => conv_std_logic_vector(0, 8),
4368 => conv_std_logic_vector(1, 8),
4369 => conv_std_logic_vector(1, 8),
4370 => conv_std_logic_vector(1, 8),
4371 => conv_std_logic_vector(1, 8),
4372 => conv_std_logic_vector(1, 8),
4373 => conv_std_logic_vector(1, 8),
4374 => conv_std_logic_vector(1, 8),
4375 => conv_std_logic_vector(1, 8),
4376 => conv_std_logic_vector(1, 8),
4377 => conv_std_logic_vector(1, 8),
4378 => conv_std_logic_vector(1, 8),
4379 => conv_std_logic_vector(1, 8),
4380 => conv_std_logic_vector(1, 8),
4381 => conv_std_logic_vector(1, 8),
4382 => conv_std_logic_vector(1, 8),
4383 => conv_std_logic_vector(2, 8),
4384 => conv_std_logic_vector(2, 8),
4385 => conv_std_logic_vector(2, 8),
4386 => conv_std_logic_vector(2, 8),
4387 => conv_std_logic_vector(2, 8),
4388 => conv_std_logic_vector(2, 8),
4389 => conv_std_logic_vector(2, 8),
4390 => conv_std_logic_vector(2, 8),
4391 => conv_std_logic_vector(2, 8),
4392 => conv_std_logic_vector(2, 8),
4393 => conv_std_logic_vector(2, 8),
4394 => conv_std_logic_vector(2, 8),
4395 => conv_std_logic_vector(2, 8),
4396 => conv_std_logic_vector(2, 8),
4397 => conv_std_logic_vector(2, 8),
4398 => conv_std_logic_vector(3, 8),
4399 => conv_std_logic_vector(3, 8),
4400 => conv_std_logic_vector(3, 8),
4401 => conv_std_logic_vector(3, 8),
4402 => conv_std_logic_vector(3, 8),
4403 => conv_std_logic_vector(3, 8),
4404 => conv_std_logic_vector(3, 8),
4405 => conv_std_logic_vector(3, 8),
4406 => conv_std_logic_vector(3, 8),
4407 => conv_std_logic_vector(3, 8),
4408 => conv_std_logic_vector(3, 8),
4409 => conv_std_logic_vector(3, 8),
4410 => conv_std_logic_vector(3, 8),
4411 => conv_std_logic_vector(3, 8),
4412 => conv_std_logic_vector(3, 8),
4413 => conv_std_logic_vector(4, 8),
4414 => conv_std_logic_vector(4, 8),
4415 => conv_std_logic_vector(4, 8),
4416 => conv_std_logic_vector(4, 8),
4417 => conv_std_logic_vector(4, 8),
4418 => conv_std_logic_vector(4, 8),
4419 => conv_std_logic_vector(4, 8),
4420 => conv_std_logic_vector(4, 8),
4421 => conv_std_logic_vector(4, 8),
4422 => conv_std_logic_vector(4, 8),
4423 => conv_std_logic_vector(4, 8),
4424 => conv_std_logic_vector(4, 8),
4425 => conv_std_logic_vector(4, 8),
4426 => conv_std_logic_vector(4, 8),
4427 => conv_std_logic_vector(4, 8),
4428 => conv_std_logic_vector(5, 8),
4429 => conv_std_logic_vector(5, 8),
4430 => conv_std_logic_vector(5, 8),
4431 => conv_std_logic_vector(5, 8),
4432 => conv_std_logic_vector(5, 8),
4433 => conv_std_logic_vector(5, 8),
4434 => conv_std_logic_vector(5, 8),
4435 => conv_std_logic_vector(5, 8),
4436 => conv_std_logic_vector(5, 8),
4437 => conv_std_logic_vector(5, 8),
4438 => conv_std_logic_vector(5, 8),
4439 => conv_std_logic_vector(5, 8),
4440 => conv_std_logic_vector(5, 8),
4441 => conv_std_logic_vector(5, 8),
4442 => conv_std_logic_vector(5, 8),
4443 => conv_std_logic_vector(6, 8),
4444 => conv_std_logic_vector(6, 8),
4445 => conv_std_logic_vector(6, 8),
4446 => conv_std_logic_vector(6, 8),
4447 => conv_std_logic_vector(6, 8),
4448 => conv_std_logic_vector(6, 8),
4449 => conv_std_logic_vector(6, 8),
4450 => conv_std_logic_vector(6, 8),
4451 => conv_std_logic_vector(6, 8),
4452 => conv_std_logic_vector(6, 8),
4453 => conv_std_logic_vector(6, 8),
4454 => conv_std_logic_vector(6, 8),
4455 => conv_std_logic_vector(6, 8),
4456 => conv_std_logic_vector(6, 8),
4457 => conv_std_logic_vector(6, 8),
4458 => conv_std_logic_vector(7, 8),
4459 => conv_std_logic_vector(7, 8),
4460 => conv_std_logic_vector(7, 8),
4461 => conv_std_logic_vector(7, 8),
4462 => conv_std_logic_vector(7, 8),
4463 => conv_std_logic_vector(7, 8),
4464 => conv_std_logic_vector(7, 8),
4465 => conv_std_logic_vector(7, 8),
4466 => conv_std_logic_vector(7, 8),
4467 => conv_std_logic_vector(7, 8),
4468 => conv_std_logic_vector(7, 8),
4469 => conv_std_logic_vector(7, 8),
4470 => conv_std_logic_vector(7, 8),
4471 => conv_std_logic_vector(7, 8),
4472 => conv_std_logic_vector(7, 8),
4473 => conv_std_logic_vector(8, 8),
4474 => conv_std_logic_vector(8, 8),
4475 => conv_std_logic_vector(8, 8),
4476 => conv_std_logic_vector(8, 8),
4477 => conv_std_logic_vector(8, 8),
4478 => conv_std_logic_vector(8, 8),
4479 => conv_std_logic_vector(8, 8),
4480 => conv_std_logic_vector(8, 8),
4481 => conv_std_logic_vector(8, 8),
4482 => conv_std_logic_vector(8, 8),
4483 => conv_std_logic_vector(8, 8),
4484 => conv_std_logic_vector(8, 8),
4485 => conv_std_logic_vector(8, 8),
4486 => conv_std_logic_vector(8, 8),
4487 => conv_std_logic_vector(8, 8),
4488 => conv_std_logic_vector(9, 8),
4489 => conv_std_logic_vector(9, 8),
4490 => conv_std_logic_vector(9, 8),
4491 => conv_std_logic_vector(9, 8),
4492 => conv_std_logic_vector(9, 8),
4493 => conv_std_logic_vector(9, 8),
4494 => conv_std_logic_vector(9, 8),
4495 => conv_std_logic_vector(9, 8),
4496 => conv_std_logic_vector(9, 8),
4497 => conv_std_logic_vector(9, 8),
4498 => conv_std_logic_vector(9, 8),
4499 => conv_std_logic_vector(9, 8),
4500 => conv_std_logic_vector(9, 8),
4501 => conv_std_logic_vector(9, 8),
4502 => conv_std_logic_vector(9, 8),
4503 => conv_std_logic_vector(10, 8),
4504 => conv_std_logic_vector(10, 8),
4505 => conv_std_logic_vector(10, 8),
4506 => conv_std_logic_vector(10, 8),
4507 => conv_std_logic_vector(10, 8),
4508 => conv_std_logic_vector(10, 8),
4509 => conv_std_logic_vector(10, 8),
4510 => conv_std_logic_vector(10, 8),
4511 => conv_std_logic_vector(10, 8),
4512 => conv_std_logic_vector(10, 8),
4513 => conv_std_logic_vector(10, 8),
4514 => conv_std_logic_vector(10, 8),
4515 => conv_std_logic_vector(10, 8),
4516 => conv_std_logic_vector(10, 8),
4517 => conv_std_logic_vector(10, 8),
4518 => conv_std_logic_vector(11, 8),
4519 => conv_std_logic_vector(11, 8),
4520 => conv_std_logic_vector(11, 8),
4521 => conv_std_logic_vector(11, 8),
4522 => conv_std_logic_vector(11, 8),
4523 => conv_std_logic_vector(11, 8),
4524 => conv_std_logic_vector(11, 8),
4525 => conv_std_logic_vector(11, 8),
4526 => conv_std_logic_vector(11, 8),
4527 => conv_std_logic_vector(11, 8),
4528 => conv_std_logic_vector(11, 8),
4529 => conv_std_logic_vector(11, 8),
4530 => conv_std_logic_vector(11, 8),
4531 => conv_std_logic_vector(11, 8),
4532 => conv_std_logic_vector(11, 8),
4533 => conv_std_logic_vector(12, 8),
4534 => conv_std_logic_vector(12, 8),
4535 => conv_std_logic_vector(12, 8),
4536 => conv_std_logic_vector(12, 8),
4537 => conv_std_logic_vector(12, 8),
4538 => conv_std_logic_vector(12, 8),
4539 => conv_std_logic_vector(12, 8),
4540 => conv_std_logic_vector(12, 8),
4541 => conv_std_logic_vector(12, 8),
4542 => conv_std_logic_vector(12, 8),
4543 => conv_std_logic_vector(12, 8),
4544 => conv_std_logic_vector(12, 8),
4545 => conv_std_logic_vector(12, 8),
4546 => conv_std_logic_vector(12, 8),
4547 => conv_std_logic_vector(12, 8),
4548 => conv_std_logic_vector(13, 8),
4549 => conv_std_logic_vector(13, 8),
4550 => conv_std_logic_vector(13, 8),
4551 => conv_std_logic_vector(13, 8),
4552 => conv_std_logic_vector(13, 8),
4553 => conv_std_logic_vector(13, 8),
4554 => conv_std_logic_vector(13, 8),
4555 => conv_std_logic_vector(13, 8),
4556 => conv_std_logic_vector(13, 8),
4557 => conv_std_logic_vector(13, 8),
4558 => conv_std_logic_vector(13, 8),
4559 => conv_std_logic_vector(13, 8),
4560 => conv_std_logic_vector(13, 8),
4561 => conv_std_logic_vector(13, 8),
4562 => conv_std_logic_vector(13, 8),
4563 => conv_std_logic_vector(14, 8),
4564 => conv_std_logic_vector(14, 8),
4565 => conv_std_logic_vector(14, 8),
4566 => conv_std_logic_vector(14, 8),
4567 => conv_std_logic_vector(14, 8),
4568 => conv_std_logic_vector(14, 8),
4569 => conv_std_logic_vector(14, 8),
4570 => conv_std_logic_vector(14, 8),
4571 => conv_std_logic_vector(14, 8),
4572 => conv_std_logic_vector(14, 8),
4573 => conv_std_logic_vector(14, 8),
4574 => conv_std_logic_vector(14, 8),
4575 => conv_std_logic_vector(14, 8),
4576 => conv_std_logic_vector(14, 8),
4577 => conv_std_logic_vector(14, 8),
4578 => conv_std_logic_vector(15, 8),
4579 => conv_std_logic_vector(15, 8),
4580 => conv_std_logic_vector(15, 8),
4581 => conv_std_logic_vector(15, 8),
4582 => conv_std_logic_vector(15, 8),
4583 => conv_std_logic_vector(15, 8),
4584 => conv_std_logic_vector(15, 8),
4585 => conv_std_logic_vector(15, 8),
4586 => conv_std_logic_vector(15, 8),
4587 => conv_std_logic_vector(15, 8),
4588 => conv_std_logic_vector(15, 8),
4589 => conv_std_logic_vector(15, 8),
4590 => conv_std_logic_vector(15, 8),
4591 => conv_std_logic_vector(15, 8),
4592 => conv_std_logic_vector(15, 8),
4593 => conv_std_logic_vector(16, 8),
4594 => conv_std_logic_vector(16, 8),
4595 => conv_std_logic_vector(16, 8),
4596 => conv_std_logic_vector(16, 8),
4597 => conv_std_logic_vector(16, 8),
4598 => conv_std_logic_vector(16, 8),
4599 => conv_std_logic_vector(16, 8),
4600 => conv_std_logic_vector(16, 8),
4601 => conv_std_logic_vector(16, 8),
4602 => conv_std_logic_vector(16, 8),
4603 => conv_std_logic_vector(16, 8),
4604 => conv_std_logic_vector(16, 8),
4605 => conv_std_logic_vector(16, 8),
4606 => conv_std_logic_vector(16, 8),
4607 => conv_std_logic_vector(16, 8),
4608 => conv_std_logic_vector(0, 8),
4609 => conv_std_logic_vector(0, 8),
4610 => conv_std_logic_vector(0, 8),
4611 => conv_std_logic_vector(0, 8),
4612 => conv_std_logic_vector(0, 8),
4613 => conv_std_logic_vector(0, 8),
4614 => conv_std_logic_vector(0, 8),
4615 => conv_std_logic_vector(0, 8),
4616 => conv_std_logic_vector(0, 8),
4617 => conv_std_logic_vector(0, 8),
4618 => conv_std_logic_vector(0, 8),
4619 => conv_std_logic_vector(0, 8),
4620 => conv_std_logic_vector(0, 8),
4621 => conv_std_logic_vector(0, 8),
4622 => conv_std_logic_vector(0, 8),
4623 => conv_std_logic_vector(1, 8),
4624 => conv_std_logic_vector(1, 8),
4625 => conv_std_logic_vector(1, 8),
4626 => conv_std_logic_vector(1, 8),
4627 => conv_std_logic_vector(1, 8),
4628 => conv_std_logic_vector(1, 8),
4629 => conv_std_logic_vector(1, 8),
4630 => conv_std_logic_vector(1, 8),
4631 => conv_std_logic_vector(1, 8),
4632 => conv_std_logic_vector(1, 8),
4633 => conv_std_logic_vector(1, 8),
4634 => conv_std_logic_vector(1, 8),
4635 => conv_std_logic_vector(1, 8),
4636 => conv_std_logic_vector(1, 8),
4637 => conv_std_logic_vector(2, 8),
4638 => conv_std_logic_vector(2, 8),
4639 => conv_std_logic_vector(2, 8),
4640 => conv_std_logic_vector(2, 8),
4641 => conv_std_logic_vector(2, 8),
4642 => conv_std_logic_vector(2, 8),
4643 => conv_std_logic_vector(2, 8),
4644 => conv_std_logic_vector(2, 8),
4645 => conv_std_logic_vector(2, 8),
4646 => conv_std_logic_vector(2, 8),
4647 => conv_std_logic_vector(2, 8),
4648 => conv_std_logic_vector(2, 8),
4649 => conv_std_logic_vector(2, 8),
4650 => conv_std_logic_vector(2, 8),
4651 => conv_std_logic_vector(3, 8),
4652 => conv_std_logic_vector(3, 8),
4653 => conv_std_logic_vector(3, 8),
4654 => conv_std_logic_vector(3, 8),
4655 => conv_std_logic_vector(3, 8),
4656 => conv_std_logic_vector(3, 8),
4657 => conv_std_logic_vector(3, 8),
4658 => conv_std_logic_vector(3, 8),
4659 => conv_std_logic_vector(3, 8),
4660 => conv_std_logic_vector(3, 8),
4661 => conv_std_logic_vector(3, 8),
4662 => conv_std_logic_vector(3, 8),
4663 => conv_std_logic_vector(3, 8),
4664 => conv_std_logic_vector(3, 8),
4665 => conv_std_logic_vector(4, 8),
4666 => conv_std_logic_vector(4, 8),
4667 => conv_std_logic_vector(4, 8),
4668 => conv_std_logic_vector(4, 8),
4669 => conv_std_logic_vector(4, 8),
4670 => conv_std_logic_vector(4, 8),
4671 => conv_std_logic_vector(4, 8),
4672 => conv_std_logic_vector(4, 8),
4673 => conv_std_logic_vector(4, 8),
4674 => conv_std_logic_vector(4, 8),
4675 => conv_std_logic_vector(4, 8),
4676 => conv_std_logic_vector(4, 8),
4677 => conv_std_logic_vector(4, 8),
4678 => conv_std_logic_vector(4, 8),
4679 => conv_std_logic_vector(4, 8),
4680 => conv_std_logic_vector(5, 8),
4681 => conv_std_logic_vector(5, 8),
4682 => conv_std_logic_vector(5, 8),
4683 => conv_std_logic_vector(5, 8),
4684 => conv_std_logic_vector(5, 8),
4685 => conv_std_logic_vector(5, 8),
4686 => conv_std_logic_vector(5, 8),
4687 => conv_std_logic_vector(5, 8),
4688 => conv_std_logic_vector(5, 8),
4689 => conv_std_logic_vector(5, 8),
4690 => conv_std_logic_vector(5, 8),
4691 => conv_std_logic_vector(5, 8),
4692 => conv_std_logic_vector(5, 8),
4693 => conv_std_logic_vector(5, 8),
4694 => conv_std_logic_vector(6, 8),
4695 => conv_std_logic_vector(6, 8),
4696 => conv_std_logic_vector(6, 8),
4697 => conv_std_logic_vector(6, 8),
4698 => conv_std_logic_vector(6, 8),
4699 => conv_std_logic_vector(6, 8),
4700 => conv_std_logic_vector(6, 8),
4701 => conv_std_logic_vector(6, 8),
4702 => conv_std_logic_vector(6, 8),
4703 => conv_std_logic_vector(6, 8),
4704 => conv_std_logic_vector(6, 8),
4705 => conv_std_logic_vector(6, 8),
4706 => conv_std_logic_vector(6, 8),
4707 => conv_std_logic_vector(6, 8),
4708 => conv_std_logic_vector(7, 8),
4709 => conv_std_logic_vector(7, 8),
4710 => conv_std_logic_vector(7, 8),
4711 => conv_std_logic_vector(7, 8),
4712 => conv_std_logic_vector(7, 8),
4713 => conv_std_logic_vector(7, 8),
4714 => conv_std_logic_vector(7, 8),
4715 => conv_std_logic_vector(7, 8),
4716 => conv_std_logic_vector(7, 8),
4717 => conv_std_logic_vector(7, 8),
4718 => conv_std_logic_vector(7, 8),
4719 => conv_std_logic_vector(7, 8),
4720 => conv_std_logic_vector(7, 8),
4721 => conv_std_logic_vector(7, 8),
4722 => conv_std_logic_vector(8, 8),
4723 => conv_std_logic_vector(8, 8),
4724 => conv_std_logic_vector(8, 8),
4725 => conv_std_logic_vector(8, 8),
4726 => conv_std_logic_vector(8, 8),
4727 => conv_std_logic_vector(8, 8),
4728 => conv_std_logic_vector(8, 8),
4729 => conv_std_logic_vector(8, 8),
4730 => conv_std_logic_vector(8, 8),
4731 => conv_std_logic_vector(8, 8),
4732 => conv_std_logic_vector(8, 8),
4733 => conv_std_logic_vector(8, 8),
4734 => conv_std_logic_vector(8, 8),
4735 => conv_std_logic_vector(8, 8),
4736 => conv_std_logic_vector(9, 8),
4737 => conv_std_logic_vector(9, 8),
4738 => conv_std_logic_vector(9, 8),
4739 => conv_std_logic_vector(9, 8),
4740 => conv_std_logic_vector(9, 8),
4741 => conv_std_logic_vector(9, 8),
4742 => conv_std_logic_vector(9, 8),
4743 => conv_std_logic_vector(9, 8),
4744 => conv_std_logic_vector(9, 8),
4745 => conv_std_logic_vector(9, 8),
4746 => conv_std_logic_vector(9, 8),
4747 => conv_std_logic_vector(9, 8),
4748 => conv_std_logic_vector(9, 8),
4749 => conv_std_logic_vector(9, 8),
4750 => conv_std_logic_vector(9, 8),
4751 => conv_std_logic_vector(10, 8),
4752 => conv_std_logic_vector(10, 8),
4753 => conv_std_logic_vector(10, 8),
4754 => conv_std_logic_vector(10, 8),
4755 => conv_std_logic_vector(10, 8),
4756 => conv_std_logic_vector(10, 8),
4757 => conv_std_logic_vector(10, 8),
4758 => conv_std_logic_vector(10, 8),
4759 => conv_std_logic_vector(10, 8),
4760 => conv_std_logic_vector(10, 8),
4761 => conv_std_logic_vector(10, 8),
4762 => conv_std_logic_vector(10, 8),
4763 => conv_std_logic_vector(10, 8),
4764 => conv_std_logic_vector(10, 8),
4765 => conv_std_logic_vector(11, 8),
4766 => conv_std_logic_vector(11, 8),
4767 => conv_std_logic_vector(11, 8),
4768 => conv_std_logic_vector(11, 8),
4769 => conv_std_logic_vector(11, 8),
4770 => conv_std_logic_vector(11, 8),
4771 => conv_std_logic_vector(11, 8),
4772 => conv_std_logic_vector(11, 8),
4773 => conv_std_logic_vector(11, 8),
4774 => conv_std_logic_vector(11, 8),
4775 => conv_std_logic_vector(11, 8),
4776 => conv_std_logic_vector(11, 8),
4777 => conv_std_logic_vector(11, 8),
4778 => conv_std_logic_vector(11, 8),
4779 => conv_std_logic_vector(12, 8),
4780 => conv_std_logic_vector(12, 8),
4781 => conv_std_logic_vector(12, 8),
4782 => conv_std_logic_vector(12, 8),
4783 => conv_std_logic_vector(12, 8),
4784 => conv_std_logic_vector(12, 8),
4785 => conv_std_logic_vector(12, 8),
4786 => conv_std_logic_vector(12, 8),
4787 => conv_std_logic_vector(12, 8),
4788 => conv_std_logic_vector(12, 8),
4789 => conv_std_logic_vector(12, 8),
4790 => conv_std_logic_vector(12, 8),
4791 => conv_std_logic_vector(12, 8),
4792 => conv_std_logic_vector(12, 8),
4793 => conv_std_logic_vector(13, 8),
4794 => conv_std_logic_vector(13, 8),
4795 => conv_std_logic_vector(13, 8),
4796 => conv_std_logic_vector(13, 8),
4797 => conv_std_logic_vector(13, 8),
4798 => conv_std_logic_vector(13, 8),
4799 => conv_std_logic_vector(13, 8),
4800 => conv_std_logic_vector(13, 8),
4801 => conv_std_logic_vector(13, 8),
4802 => conv_std_logic_vector(13, 8),
4803 => conv_std_logic_vector(13, 8),
4804 => conv_std_logic_vector(13, 8),
4805 => conv_std_logic_vector(13, 8),
4806 => conv_std_logic_vector(13, 8),
4807 => conv_std_logic_vector(13, 8),
4808 => conv_std_logic_vector(14, 8),
4809 => conv_std_logic_vector(14, 8),
4810 => conv_std_logic_vector(14, 8),
4811 => conv_std_logic_vector(14, 8),
4812 => conv_std_logic_vector(14, 8),
4813 => conv_std_logic_vector(14, 8),
4814 => conv_std_logic_vector(14, 8),
4815 => conv_std_logic_vector(14, 8),
4816 => conv_std_logic_vector(14, 8),
4817 => conv_std_logic_vector(14, 8),
4818 => conv_std_logic_vector(14, 8),
4819 => conv_std_logic_vector(14, 8),
4820 => conv_std_logic_vector(14, 8),
4821 => conv_std_logic_vector(14, 8),
4822 => conv_std_logic_vector(15, 8),
4823 => conv_std_logic_vector(15, 8),
4824 => conv_std_logic_vector(15, 8),
4825 => conv_std_logic_vector(15, 8),
4826 => conv_std_logic_vector(15, 8),
4827 => conv_std_logic_vector(15, 8),
4828 => conv_std_logic_vector(15, 8),
4829 => conv_std_logic_vector(15, 8),
4830 => conv_std_logic_vector(15, 8),
4831 => conv_std_logic_vector(15, 8),
4832 => conv_std_logic_vector(15, 8),
4833 => conv_std_logic_vector(15, 8),
4834 => conv_std_logic_vector(15, 8),
4835 => conv_std_logic_vector(15, 8),
4836 => conv_std_logic_vector(16, 8),
4837 => conv_std_logic_vector(16, 8),
4838 => conv_std_logic_vector(16, 8),
4839 => conv_std_logic_vector(16, 8),
4840 => conv_std_logic_vector(16, 8),
4841 => conv_std_logic_vector(16, 8),
4842 => conv_std_logic_vector(16, 8),
4843 => conv_std_logic_vector(16, 8),
4844 => conv_std_logic_vector(16, 8),
4845 => conv_std_logic_vector(16, 8),
4846 => conv_std_logic_vector(16, 8),
4847 => conv_std_logic_vector(16, 8),
4848 => conv_std_logic_vector(16, 8),
4849 => conv_std_logic_vector(16, 8),
4850 => conv_std_logic_vector(17, 8),
4851 => conv_std_logic_vector(17, 8),
4852 => conv_std_logic_vector(17, 8),
4853 => conv_std_logic_vector(17, 8),
4854 => conv_std_logic_vector(17, 8),
4855 => conv_std_logic_vector(17, 8),
4856 => conv_std_logic_vector(17, 8),
4857 => conv_std_logic_vector(17, 8),
4858 => conv_std_logic_vector(17, 8),
4859 => conv_std_logic_vector(17, 8),
4860 => conv_std_logic_vector(17, 8),
4861 => conv_std_logic_vector(17, 8),
4862 => conv_std_logic_vector(17, 8),
4863 => conv_std_logic_vector(17, 8),
4864 => conv_std_logic_vector(0, 8),
4865 => conv_std_logic_vector(0, 8),
4866 => conv_std_logic_vector(0, 8),
4867 => conv_std_logic_vector(0, 8),
4868 => conv_std_logic_vector(0, 8),
4869 => conv_std_logic_vector(0, 8),
4870 => conv_std_logic_vector(0, 8),
4871 => conv_std_logic_vector(0, 8),
4872 => conv_std_logic_vector(0, 8),
4873 => conv_std_logic_vector(0, 8),
4874 => conv_std_logic_vector(0, 8),
4875 => conv_std_logic_vector(0, 8),
4876 => conv_std_logic_vector(0, 8),
4877 => conv_std_logic_vector(0, 8),
4878 => conv_std_logic_vector(1, 8),
4879 => conv_std_logic_vector(1, 8),
4880 => conv_std_logic_vector(1, 8),
4881 => conv_std_logic_vector(1, 8),
4882 => conv_std_logic_vector(1, 8),
4883 => conv_std_logic_vector(1, 8),
4884 => conv_std_logic_vector(1, 8),
4885 => conv_std_logic_vector(1, 8),
4886 => conv_std_logic_vector(1, 8),
4887 => conv_std_logic_vector(1, 8),
4888 => conv_std_logic_vector(1, 8),
4889 => conv_std_logic_vector(1, 8),
4890 => conv_std_logic_vector(1, 8),
4891 => conv_std_logic_vector(2, 8),
4892 => conv_std_logic_vector(2, 8),
4893 => conv_std_logic_vector(2, 8),
4894 => conv_std_logic_vector(2, 8),
4895 => conv_std_logic_vector(2, 8),
4896 => conv_std_logic_vector(2, 8),
4897 => conv_std_logic_vector(2, 8),
4898 => conv_std_logic_vector(2, 8),
4899 => conv_std_logic_vector(2, 8),
4900 => conv_std_logic_vector(2, 8),
4901 => conv_std_logic_vector(2, 8),
4902 => conv_std_logic_vector(2, 8),
4903 => conv_std_logic_vector(2, 8),
4904 => conv_std_logic_vector(2, 8),
4905 => conv_std_logic_vector(3, 8),
4906 => conv_std_logic_vector(3, 8),
4907 => conv_std_logic_vector(3, 8),
4908 => conv_std_logic_vector(3, 8),
4909 => conv_std_logic_vector(3, 8),
4910 => conv_std_logic_vector(3, 8),
4911 => conv_std_logic_vector(3, 8),
4912 => conv_std_logic_vector(3, 8),
4913 => conv_std_logic_vector(3, 8),
4914 => conv_std_logic_vector(3, 8),
4915 => conv_std_logic_vector(3, 8),
4916 => conv_std_logic_vector(3, 8),
4917 => conv_std_logic_vector(3, 8),
4918 => conv_std_logic_vector(4, 8),
4919 => conv_std_logic_vector(4, 8),
4920 => conv_std_logic_vector(4, 8),
4921 => conv_std_logic_vector(4, 8),
4922 => conv_std_logic_vector(4, 8),
4923 => conv_std_logic_vector(4, 8),
4924 => conv_std_logic_vector(4, 8),
4925 => conv_std_logic_vector(4, 8),
4926 => conv_std_logic_vector(4, 8),
4927 => conv_std_logic_vector(4, 8),
4928 => conv_std_logic_vector(4, 8),
4929 => conv_std_logic_vector(4, 8),
4930 => conv_std_logic_vector(4, 8),
4931 => conv_std_logic_vector(4, 8),
4932 => conv_std_logic_vector(5, 8),
4933 => conv_std_logic_vector(5, 8),
4934 => conv_std_logic_vector(5, 8),
4935 => conv_std_logic_vector(5, 8),
4936 => conv_std_logic_vector(5, 8),
4937 => conv_std_logic_vector(5, 8),
4938 => conv_std_logic_vector(5, 8),
4939 => conv_std_logic_vector(5, 8),
4940 => conv_std_logic_vector(5, 8),
4941 => conv_std_logic_vector(5, 8),
4942 => conv_std_logic_vector(5, 8),
4943 => conv_std_logic_vector(5, 8),
4944 => conv_std_logic_vector(5, 8),
4945 => conv_std_logic_vector(6, 8),
4946 => conv_std_logic_vector(6, 8),
4947 => conv_std_logic_vector(6, 8),
4948 => conv_std_logic_vector(6, 8),
4949 => conv_std_logic_vector(6, 8),
4950 => conv_std_logic_vector(6, 8),
4951 => conv_std_logic_vector(6, 8),
4952 => conv_std_logic_vector(6, 8),
4953 => conv_std_logic_vector(6, 8),
4954 => conv_std_logic_vector(6, 8),
4955 => conv_std_logic_vector(6, 8),
4956 => conv_std_logic_vector(6, 8),
4957 => conv_std_logic_vector(6, 8),
4958 => conv_std_logic_vector(6, 8),
4959 => conv_std_logic_vector(7, 8),
4960 => conv_std_logic_vector(7, 8),
4961 => conv_std_logic_vector(7, 8),
4962 => conv_std_logic_vector(7, 8),
4963 => conv_std_logic_vector(7, 8),
4964 => conv_std_logic_vector(7, 8),
4965 => conv_std_logic_vector(7, 8),
4966 => conv_std_logic_vector(7, 8),
4967 => conv_std_logic_vector(7, 8),
4968 => conv_std_logic_vector(7, 8),
4969 => conv_std_logic_vector(7, 8),
4970 => conv_std_logic_vector(7, 8),
4971 => conv_std_logic_vector(7, 8),
4972 => conv_std_logic_vector(8, 8),
4973 => conv_std_logic_vector(8, 8),
4974 => conv_std_logic_vector(8, 8),
4975 => conv_std_logic_vector(8, 8),
4976 => conv_std_logic_vector(8, 8),
4977 => conv_std_logic_vector(8, 8),
4978 => conv_std_logic_vector(8, 8),
4979 => conv_std_logic_vector(8, 8),
4980 => conv_std_logic_vector(8, 8),
4981 => conv_std_logic_vector(8, 8),
4982 => conv_std_logic_vector(8, 8),
4983 => conv_std_logic_vector(8, 8),
4984 => conv_std_logic_vector(8, 8),
4985 => conv_std_logic_vector(8, 8),
4986 => conv_std_logic_vector(9, 8),
4987 => conv_std_logic_vector(9, 8),
4988 => conv_std_logic_vector(9, 8),
4989 => conv_std_logic_vector(9, 8),
4990 => conv_std_logic_vector(9, 8),
4991 => conv_std_logic_vector(9, 8),
4992 => conv_std_logic_vector(9, 8),
4993 => conv_std_logic_vector(9, 8),
4994 => conv_std_logic_vector(9, 8),
4995 => conv_std_logic_vector(9, 8),
4996 => conv_std_logic_vector(9, 8),
4997 => conv_std_logic_vector(9, 8),
4998 => conv_std_logic_vector(9, 8),
4999 => conv_std_logic_vector(10, 8),
5000 => conv_std_logic_vector(10, 8),
5001 => conv_std_logic_vector(10, 8),
5002 => conv_std_logic_vector(10, 8),
5003 => conv_std_logic_vector(10, 8),
5004 => conv_std_logic_vector(10, 8),
5005 => conv_std_logic_vector(10, 8),
5006 => conv_std_logic_vector(10, 8),
5007 => conv_std_logic_vector(10, 8),
5008 => conv_std_logic_vector(10, 8),
5009 => conv_std_logic_vector(10, 8),
5010 => conv_std_logic_vector(10, 8),
5011 => conv_std_logic_vector(10, 8),
5012 => conv_std_logic_vector(10, 8),
5013 => conv_std_logic_vector(11, 8),
5014 => conv_std_logic_vector(11, 8),
5015 => conv_std_logic_vector(11, 8),
5016 => conv_std_logic_vector(11, 8),
5017 => conv_std_logic_vector(11, 8),
5018 => conv_std_logic_vector(11, 8),
5019 => conv_std_logic_vector(11, 8),
5020 => conv_std_logic_vector(11, 8),
5021 => conv_std_logic_vector(11, 8),
5022 => conv_std_logic_vector(11, 8),
5023 => conv_std_logic_vector(11, 8),
5024 => conv_std_logic_vector(11, 8),
5025 => conv_std_logic_vector(11, 8),
5026 => conv_std_logic_vector(12, 8),
5027 => conv_std_logic_vector(12, 8),
5028 => conv_std_logic_vector(12, 8),
5029 => conv_std_logic_vector(12, 8),
5030 => conv_std_logic_vector(12, 8),
5031 => conv_std_logic_vector(12, 8),
5032 => conv_std_logic_vector(12, 8),
5033 => conv_std_logic_vector(12, 8),
5034 => conv_std_logic_vector(12, 8),
5035 => conv_std_logic_vector(12, 8),
5036 => conv_std_logic_vector(12, 8),
5037 => conv_std_logic_vector(12, 8),
5038 => conv_std_logic_vector(12, 8),
5039 => conv_std_logic_vector(12, 8),
5040 => conv_std_logic_vector(13, 8),
5041 => conv_std_logic_vector(13, 8),
5042 => conv_std_logic_vector(13, 8),
5043 => conv_std_logic_vector(13, 8),
5044 => conv_std_logic_vector(13, 8),
5045 => conv_std_logic_vector(13, 8),
5046 => conv_std_logic_vector(13, 8),
5047 => conv_std_logic_vector(13, 8),
5048 => conv_std_logic_vector(13, 8),
5049 => conv_std_logic_vector(13, 8),
5050 => conv_std_logic_vector(13, 8),
5051 => conv_std_logic_vector(13, 8),
5052 => conv_std_logic_vector(13, 8),
5053 => conv_std_logic_vector(14, 8),
5054 => conv_std_logic_vector(14, 8),
5055 => conv_std_logic_vector(14, 8),
5056 => conv_std_logic_vector(14, 8),
5057 => conv_std_logic_vector(14, 8),
5058 => conv_std_logic_vector(14, 8),
5059 => conv_std_logic_vector(14, 8),
5060 => conv_std_logic_vector(14, 8),
5061 => conv_std_logic_vector(14, 8),
5062 => conv_std_logic_vector(14, 8),
5063 => conv_std_logic_vector(14, 8),
5064 => conv_std_logic_vector(14, 8),
5065 => conv_std_logic_vector(14, 8),
5066 => conv_std_logic_vector(14, 8),
5067 => conv_std_logic_vector(15, 8),
5068 => conv_std_logic_vector(15, 8),
5069 => conv_std_logic_vector(15, 8),
5070 => conv_std_logic_vector(15, 8),
5071 => conv_std_logic_vector(15, 8),
5072 => conv_std_logic_vector(15, 8),
5073 => conv_std_logic_vector(15, 8),
5074 => conv_std_logic_vector(15, 8),
5075 => conv_std_logic_vector(15, 8),
5076 => conv_std_logic_vector(15, 8),
5077 => conv_std_logic_vector(15, 8),
5078 => conv_std_logic_vector(15, 8),
5079 => conv_std_logic_vector(15, 8),
5080 => conv_std_logic_vector(16, 8),
5081 => conv_std_logic_vector(16, 8),
5082 => conv_std_logic_vector(16, 8),
5083 => conv_std_logic_vector(16, 8),
5084 => conv_std_logic_vector(16, 8),
5085 => conv_std_logic_vector(16, 8),
5086 => conv_std_logic_vector(16, 8),
5087 => conv_std_logic_vector(16, 8),
5088 => conv_std_logic_vector(16, 8),
5089 => conv_std_logic_vector(16, 8),
5090 => conv_std_logic_vector(16, 8),
5091 => conv_std_logic_vector(16, 8),
5092 => conv_std_logic_vector(16, 8),
5093 => conv_std_logic_vector(16, 8),
5094 => conv_std_logic_vector(17, 8),
5095 => conv_std_logic_vector(17, 8),
5096 => conv_std_logic_vector(17, 8),
5097 => conv_std_logic_vector(17, 8),
5098 => conv_std_logic_vector(17, 8),
5099 => conv_std_logic_vector(17, 8),
5100 => conv_std_logic_vector(17, 8),
5101 => conv_std_logic_vector(17, 8),
5102 => conv_std_logic_vector(17, 8),
5103 => conv_std_logic_vector(17, 8),
5104 => conv_std_logic_vector(17, 8),
5105 => conv_std_logic_vector(17, 8),
5106 => conv_std_logic_vector(17, 8),
5107 => conv_std_logic_vector(18, 8),
5108 => conv_std_logic_vector(18, 8),
5109 => conv_std_logic_vector(18, 8),
5110 => conv_std_logic_vector(18, 8),
5111 => conv_std_logic_vector(18, 8),
5112 => conv_std_logic_vector(18, 8),
5113 => conv_std_logic_vector(18, 8),
5114 => conv_std_logic_vector(18, 8),
5115 => conv_std_logic_vector(18, 8),
5116 => conv_std_logic_vector(18, 8),
5117 => conv_std_logic_vector(18, 8),
5118 => conv_std_logic_vector(18, 8),
5119 => conv_std_logic_vector(18, 8),
5120 => conv_std_logic_vector(0, 8),
5121 => conv_std_logic_vector(0, 8),
5122 => conv_std_logic_vector(0, 8),
5123 => conv_std_logic_vector(0, 8),
5124 => conv_std_logic_vector(0, 8),
5125 => conv_std_logic_vector(0, 8),
5126 => conv_std_logic_vector(0, 8),
5127 => conv_std_logic_vector(0, 8),
5128 => conv_std_logic_vector(0, 8),
5129 => conv_std_logic_vector(0, 8),
5130 => conv_std_logic_vector(0, 8),
5131 => conv_std_logic_vector(0, 8),
5132 => conv_std_logic_vector(0, 8),
5133 => conv_std_logic_vector(1, 8),
5134 => conv_std_logic_vector(1, 8),
5135 => conv_std_logic_vector(1, 8),
5136 => conv_std_logic_vector(1, 8),
5137 => conv_std_logic_vector(1, 8),
5138 => conv_std_logic_vector(1, 8),
5139 => conv_std_logic_vector(1, 8),
5140 => conv_std_logic_vector(1, 8),
5141 => conv_std_logic_vector(1, 8),
5142 => conv_std_logic_vector(1, 8),
5143 => conv_std_logic_vector(1, 8),
5144 => conv_std_logic_vector(1, 8),
5145 => conv_std_logic_vector(1, 8),
5146 => conv_std_logic_vector(2, 8),
5147 => conv_std_logic_vector(2, 8),
5148 => conv_std_logic_vector(2, 8),
5149 => conv_std_logic_vector(2, 8),
5150 => conv_std_logic_vector(2, 8),
5151 => conv_std_logic_vector(2, 8),
5152 => conv_std_logic_vector(2, 8),
5153 => conv_std_logic_vector(2, 8),
5154 => conv_std_logic_vector(2, 8),
5155 => conv_std_logic_vector(2, 8),
5156 => conv_std_logic_vector(2, 8),
5157 => conv_std_logic_vector(2, 8),
5158 => conv_std_logic_vector(2, 8),
5159 => conv_std_logic_vector(3, 8),
5160 => conv_std_logic_vector(3, 8),
5161 => conv_std_logic_vector(3, 8),
5162 => conv_std_logic_vector(3, 8),
5163 => conv_std_logic_vector(3, 8),
5164 => conv_std_logic_vector(3, 8),
5165 => conv_std_logic_vector(3, 8),
5166 => conv_std_logic_vector(3, 8),
5167 => conv_std_logic_vector(3, 8),
5168 => conv_std_logic_vector(3, 8),
5169 => conv_std_logic_vector(3, 8),
5170 => conv_std_logic_vector(3, 8),
5171 => conv_std_logic_vector(3, 8),
5172 => conv_std_logic_vector(4, 8),
5173 => conv_std_logic_vector(4, 8),
5174 => conv_std_logic_vector(4, 8),
5175 => conv_std_logic_vector(4, 8),
5176 => conv_std_logic_vector(4, 8),
5177 => conv_std_logic_vector(4, 8),
5178 => conv_std_logic_vector(4, 8),
5179 => conv_std_logic_vector(4, 8),
5180 => conv_std_logic_vector(4, 8),
5181 => conv_std_logic_vector(4, 8),
5182 => conv_std_logic_vector(4, 8),
5183 => conv_std_logic_vector(4, 8),
5184 => conv_std_logic_vector(5, 8),
5185 => conv_std_logic_vector(5, 8),
5186 => conv_std_logic_vector(5, 8),
5187 => conv_std_logic_vector(5, 8),
5188 => conv_std_logic_vector(5, 8),
5189 => conv_std_logic_vector(5, 8),
5190 => conv_std_logic_vector(5, 8),
5191 => conv_std_logic_vector(5, 8),
5192 => conv_std_logic_vector(5, 8),
5193 => conv_std_logic_vector(5, 8),
5194 => conv_std_logic_vector(5, 8),
5195 => conv_std_logic_vector(5, 8),
5196 => conv_std_logic_vector(5, 8),
5197 => conv_std_logic_vector(6, 8),
5198 => conv_std_logic_vector(6, 8),
5199 => conv_std_logic_vector(6, 8),
5200 => conv_std_logic_vector(6, 8),
5201 => conv_std_logic_vector(6, 8),
5202 => conv_std_logic_vector(6, 8),
5203 => conv_std_logic_vector(6, 8),
5204 => conv_std_logic_vector(6, 8),
5205 => conv_std_logic_vector(6, 8),
5206 => conv_std_logic_vector(6, 8),
5207 => conv_std_logic_vector(6, 8),
5208 => conv_std_logic_vector(6, 8),
5209 => conv_std_logic_vector(6, 8),
5210 => conv_std_logic_vector(7, 8),
5211 => conv_std_logic_vector(7, 8),
5212 => conv_std_logic_vector(7, 8),
5213 => conv_std_logic_vector(7, 8),
5214 => conv_std_logic_vector(7, 8),
5215 => conv_std_logic_vector(7, 8),
5216 => conv_std_logic_vector(7, 8),
5217 => conv_std_logic_vector(7, 8),
5218 => conv_std_logic_vector(7, 8),
5219 => conv_std_logic_vector(7, 8),
5220 => conv_std_logic_vector(7, 8),
5221 => conv_std_logic_vector(7, 8),
5222 => conv_std_logic_vector(7, 8),
5223 => conv_std_logic_vector(8, 8),
5224 => conv_std_logic_vector(8, 8),
5225 => conv_std_logic_vector(8, 8),
5226 => conv_std_logic_vector(8, 8),
5227 => conv_std_logic_vector(8, 8),
5228 => conv_std_logic_vector(8, 8),
5229 => conv_std_logic_vector(8, 8),
5230 => conv_std_logic_vector(8, 8),
5231 => conv_std_logic_vector(8, 8),
5232 => conv_std_logic_vector(8, 8),
5233 => conv_std_logic_vector(8, 8),
5234 => conv_std_logic_vector(8, 8),
5235 => conv_std_logic_vector(8, 8),
5236 => conv_std_logic_vector(9, 8),
5237 => conv_std_logic_vector(9, 8),
5238 => conv_std_logic_vector(9, 8),
5239 => conv_std_logic_vector(9, 8),
5240 => conv_std_logic_vector(9, 8),
5241 => conv_std_logic_vector(9, 8),
5242 => conv_std_logic_vector(9, 8),
5243 => conv_std_logic_vector(9, 8),
5244 => conv_std_logic_vector(9, 8),
5245 => conv_std_logic_vector(9, 8),
5246 => conv_std_logic_vector(9, 8),
5247 => conv_std_logic_vector(9, 8),
5248 => conv_std_logic_vector(10, 8),
5249 => conv_std_logic_vector(10, 8),
5250 => conv_std_logic_vector(10, 8),
5251 => conv_std_logic_vector(10, 8),
5252 => conv_std_logic_vector(10, 8),
5253 => conv_std_logic_vector(10, 8),
5254 => conv_std_logic_vector(10, 8),
5255 => conv_std_logic_vector(10, 8),
5256 => conv_std_logic_vector(10, 8),
5257 => conv_std_logic_vector(10, 8),
5258 => conv_std_logic_vector(10, 8),
5259 => conv_std_logic_vector(10, 8),
5260 => conv_std_logic_vector(10, 8),
5261 => conv_std_logic_vector(11, 8),
5262 => conv_std_logic_vector(11, 8),
5263 => conv_std_logic_vector(11, 8),
5264 => conv_std_logic_vector(11, 8),
5265 => conv_std_logic_vector(11, 8),
5266 => conv_std_logic_vector(11, 8),
5267 => conv_std_logic_vector(11, 8),
5268 => conv_std_logic_vector(11, 8),
5269 => conv_std_logic_vector(11, 8),
5270 => conv_std_logic_vector(11, 8),
5271 => conv_std_logic_vector(11, 8),
5272 => conv_std_logic_vector(11, 8),
5273 => conv_std_logic_vector(11, 8),
5274 => conv_std_logic_vector(12, 8),
5275 => conv_std_logic_vector(12, 8),
5276 => conv_std_logic_vector(12, 8),
5277 => conv_std_logic_vector(12, 8),
5278 => conv_std_logic_vector(12, 8),
5279 => conv_std_logic_vector(12, 8),
5280 => conv_std_logic_vector(12, 8),
5281 => conv_std_logic_vector(12, 8),
5282 => conv_std_logic_vector(12, 8),
5283 => conv_std_logic_vector(12, 8),
5284 => conv_std_logic_vector(12, 8),
5285 => conv_std_logic_vector(12, 8),
5286 => conv_std_logic_vector(12, 8),
5287 => conv_std_logic_vector(13, 8),
5288 => conv_std_logic_vector(13, 8),
5289 => conv_std_logic_vector(13, 8),
5290 => conv_std_logic_vector(13, 8),
5291 => conv_std_logic_vector(13, 8),
5292 => conv_std_logic_vector(13, 8),
5293 => conv_std_logic_vector(13, 8),
5294 => conv_std_logic_vector(13, 8),
5295 => conv_std_logic_vector(13, 8),
5296 => conv_std_logic_vector(13, 8),
5297 => conv_std_logic_vector(13, 8),
5298 => conv_std_logic_vector(13, 8),
5299 => conv_std_logic_vector(13, 8),
5300 => conv_std_logic_vector(14, 8),
5301 => conv_std_logic_vector(14, 8),
5302 => conv_std_logic_vector(14, 8),
5303 => conv_std_logic_vector(14, 8),
5304 => conv_std_logic_vector(14, 8),
5305 => conv_std_logic_vector(14, 8),
5306 => conv_std_logic_vector(14, 8),
5307 => conv_std_logic_vector(14, 8),
5308 => conv_std_logic_vector(14, 8),
5309 => conv_std_logic_vector(14, 8),
5310 => conv_std_logic_vector(14, 8),
5311 => conv_std_logic_vector(14, 8),
5312 => conv_std_logic_vector(15, 8),
5313 => conv_std_logic_vector(15, 8),
5314 => conv_std_logic_vector(15, 8),
5315 => conv_std_logic_vector(15, 8),
5316 => conv_std_logic_vector(15, 8),
5317 => conv_std_logic_vector(15, 8),
5318 => conv_std_logic_vector(15, 8),
5319 => conv_std_logic_vector(15, 8),
5320 => conv_std_logic_vector(15, 8),
5321 => conv_std_logic_vector(15, 8),
5322 => conv_std_logic_vector(15, 8),
5323 => conv_std_logic_vector(15, 8),
5324 => conv_std_logic_vector(15, 8),
5325 => conv_std_logic_vector(16, 8),
5326 => conv_std_logic_vector(16, 8),
5327 => conv_std_logic_vector(16, 8),
5328 => conv_std_logic_vector(16, 8),
5329 => conv_std_logic_vector(16, 8),
5330 => conv_std_logic_vector(16, 8),
5331 => conv_std_logic_vector(16, 8),
5332 => conv_std_logic_vector(16, 8),
5333 => conv_std_logic_vector(16, 8),
5334 => conv_std_logic_vector(16, 8),
5335 => conv_std_logic_vector(16, 8),
5336 => conv_std_logic_vector(16, 8),
5337 => conv_std_logic_vector(16, 8),
5338 => conv_std_logic_vector(17, 8),
5339 => conv_std_logic_vector(17, 8),
5340 => conv_std_logic_vector(17, 8),
5341 => conv_std_logic_vector(17, 8),
5342 => conv_std_logic_vector(17, 8),
5343 => conv_std_logic_vector(17, 8),
5344 => conv_std_logic_vector(17, 8),
5345 => conv_std_logic_vector(17, 8),
5346 => conv_std_logic_vector(17, 8),
5347 => conv_std_logic_vector(17, 8),
5348 => conv_std_logic_vector(17, 8),
5349 => conv_std_logic_vector(17, 8),
5350 => conv_std_logic_vector(17, 8),
5351 => conv_std_logic_vector(18, 8),
5352 => conv_std_logic_vector(18, 8),
5353 => conv_std_logic_vector(18, 8),
5354 => conv_std_logic_vector(18, 8),
5355 => conv_std_logic_vector(18, 8),
5356 => conv_std_logic_vector(18, 8),
5357 => conv_std_logic_vector(18, 8),
5358 => conv_std_logic_vector(18, 8),
5359 => conv_std_logic_vector(18, 8),
5360 => conv_std_logic_vector(18, 8),
5361 => conv_std_logic_vector(18, 8),
5362 => conv_std_logic_vector(18, 8),
5363 => conv_std_logic_vector(18, 8),
5364 => conv_std_logic_vector(19, 8),
5365 => conv_std_logic_vector(19, 8),
5366 => conv_std_logic_vector(19, 8),
5367 => conv_std_logic_vector(19, 8),
5368 => conv_std_logic_vector(19, 8),
5369 => conv_std_logic_vector(19, 8),
5370 => conv_std_logic_vector(19, 8),
5371 => conv_std_logic_vector(19, 8),
5372 => conv_std_logic_vector(19, 8),
5373 => conv_std_logic_vector(19, 8),
5374 => conv_std_logic_vector(19, 8),
5375 => conv_std_logic_vector(19, 8),
5376 => conv_std_logic_vector(0, 8),
5377 => conv_std_logic_vector(0, 8),
5378 => conv_std_logic_vector(0, 8),
5379 => conv_std_logic_vector(0, 8),
5380 => conv_std_logic_vector(0, 8),
5381 => conv_std_logic_vector(0, 8),
5382 => conv_std_logic_vector(0, 8),
5383 => conv_std_logic_vector(0, 8),
5384 => conv_std_logic_vector(0, 8),
5385 => conv_std_logic_vector(0, 8),
5386 => conv_std_logic_vector(0, 8),
5387 => conv_std_logic_vector(0, 8),
5388 => conv_std_logic_vector(0, 8),
5389 => conv_std_logic_vector(1, 8),
5390 => conv_std_logic_vector(1, 8),
5391 => conv_std_logic_vector(1, 8),
5392 => conv_std_logic_vector(1, 8),
5393 => conv_std_logic_vector(1, 8),
5394 => conv_std_logic_vector(1, 8),
5395 => conv_std_logic_vector(1, 8),
5396 => conv_std_logic_vector(1, 8),
5397 => conv_std_logic_vector(1, 8),
5398 => conv_std_logic_vector(1, 8),
5399 => conv_std_logic_vector(1, 8),
5400 => conv_std_logic_vector(1, 8),
5401 => conv_std_logic_vector(2, 8),
5402 => conv_std_logic_vector(2, 8),
5403 => conv_std_logic_vector(2, 8),
5404 => conv_std_logic_vector(2, 8),
5405 => conv_std_logic_vector(2, 8),
5406 => conv_std_logic_vector(2, 8),
5407 => conv_std_logic_vector(2, 8),
5408 => conv_std_logic_vector(2, 8),
5409 => conv_std_logic_vector(2, 8),
5410 => conv_std_logic_vector(2, 8),
5411 => conv_std_logic_vector(2, 8),
5412 => conv_std_logic_vector(2, 8),
5413 => conv_std_logic_vector(3, 8),
5414 => conv_std_logic_vector(3, 8),
5415 => conv_std_logic_vector(3, 8),
5416 => conv_std_logic_vector(3, 8),
5417 => conv_std_logic_vector(3, 8),
5418 => conv_std_logic_vector(3, 8),
5419 => conv_std_logic_vector(3, 8),
5420 => conv_std_logic_vector(3, 8),
5421 => conv_std_logic_vector(3, 8),
5422 => conv_std_logic_vector(3, 8),
5423 => conv_std_logic_vector(3, 8),
5424 => conv_std_logic_vector(3, 8),
5425 => conv_std_logic_vector(4, 8),
5426 => conv_std_logic_vector(4, 8),
5427 => conv_std_logic_vector(4, 8),
5428 => conv_std_logic_vector(4, 8),
5429 => conv_std_logic_vector(4, 8),
5430 => conv_std_logic_vector(4, 8),
5431 => conv_std_logic_vector(4, 8),
5432 => conv_std_logic_vector(4, 8),
5433 => conv_std_logic_vector(4, 8),
5434 => conv_std_logic_vector(4, 8),
5435 => conv_std_logic_vector(4, 8),
5436 => conv_std_logic_vector(4, 8),
5437 => conv_std_logic_vector(5, 8),
5438 => conv_std_logic_vector(5, 8),
5439 => conv_std_logic_vector(5, 8),
5440 => conv_std_logic_vector(5, 8),
5441 => conv_std_logic_vector(5, 8),
5442 => conv_std_logic_vector(5, 8),
5443 => conv_std_logic_vector(5, 8),
5444 => conv_std_logic_vector(5, 8),
5445 => conv_std_logic_vector(5, 8),
5446 => conv_std_logic_vector(5, 8),
5447 => conv_std_logic_vector(5, 8),
5448 => conv_std_logic_vector(5, 8),
5449 => conv_std_logic_vector(5, 8),
5450 => conv_std_logic_vector(6, 8),
5451 => conv_std_logic_vector(6, 8),
5452 => conv_std_logic_vector(6, 8),
5453 => conv_std_logic_vector(6, 8),
5454 => conv_std_logic_vector(6, 8),
5455 => conv_std_logic_vector(6, 8),
5456 => conv_std_logic_vector(6, 8),
5457 => conv_std_logic_vector(6, 8),
5458 => conv_std_logic_vector(6, 8),
5459 => conv_std_logic_vector(6, 8),
5460 => conv_std_logic_vector(6, 8),
5461 => conv_std_logic_vector(6, 8),
5462 => conv_std_logic_vector(7, 8),
5463 => conv_std_logic_vector(7, 8),
5464 => conv_std_logic_vector(7, 8),
5465 => conv_std_logic_vector(7, 8),
5466 => conv_std_logic_vector(7, 8),
5467 => conv_std_logic_vector(7, 8),
5468 => conv_std_logic_vector(7, 8),
5469 => conv_std_logic_vector(7, 8),
5470 => conv_std_logic_vector(7, 8),
5471 => conv_std_logic_vector(7, 8),
5472 => conv_std_logic_vector(7, 8),
5473 => conv_std_logic_vector(7, 8),
5474 => conv_std_logic_vector(8, 8),
5475 => conv_std_logic_vector(8, 8),
5476 => conv_std_logic_vector(8, 8),
5477 => conv_std_logic_vector(8, 8),
5478 => conv_std_logic_vector(8, 8),
5479 => conv_std_logic_vector(8, 8),
5480 => conv_std_logic_vector(8, 8),
5481 => conv_std_logic_vector(8, 8),
5482 => conv_std_logic_vector(8, 8),
5483 => conv_std_logic_vector(8, 8),
5484 => conv_std_logic_vector(8, 8),
5485 => conv_std_logic_vector(8, 8),
5486 => conv_std_logic_vector(9, 8),
5487 => conv_std_logic_vector(9, 8),
5488 => conv_std_logic_vector(9, 8),
5489 => conv_std_logic_vector(9, 8),
5490 => conv_std_logic_vector(9, 8),
5491 => conv_std_logic_vector(9, 8),
5492 => conv_std_logic_vector(9, 8),
5493 => conv_std_logic_vector(9, 8),
5494 => conv_std_logic_vector(9, 8),
5495 => conv_std_logic_vector(9, 8),
5496 => conv_std_logic_vector(9, 8),
5497 => conv_std_logic_vector(9, 8),
5498 => conv_std_logic_vector(10, 8),
5499 => conv_std_logic_vector(10, 8),
5500 => conv_std_logic_vector(10, 8),
5501 => conv_std_logic_vector(10, 8),
5502 => conv_std_logic_vector(10, 8),
5503 => conv_std_logic_vector(10, 8),
5504 => conv_std_logic_vector(10, 8),
5505 => conv_std_logic_vector(10, 8),
5506 => conv_std_logic_vector(10, 8),
5507 => conv_std_logic_vector(10, 8),
5508 => conv_std_logic_vector(10, 8),
5509 => conv_std_logic_vector(10, 8),
5510 => conv_std_logic_vector(10, 8),
5511 => conv_std_logic_vector(11, 8),
5512 => conv_std_logic_vector(11, 8),
5513 => conv_std_logic_vector(11, 8),
5514 => conv_std_logic_vector(11, 8),
5515 => conv_std_logic_vector(11, 8),
5516 => conv_std_logic_vector(11, 8),
5517 => conv_std_logic_vector(11, 8),
5518 => conv_std_logic_vector(11, 8),
5519 => conv_std_logic_vector(11, 8),
5520 => conv_std_logic_vector(11, 8),
5521 => conv_std_logic_vector(11, 8),
5522 => conv_std_logic_vector(11, 8),
5523 => conv_std_logic_vector(12, 8),
5524 => conv_std_logic_vector(12, 8),
5525 => conv_std_logic_vector(12, 8),
5526 => conv_std_logic_vector(12, 8),
5527 => conv_std_logic_vector(12, 8),
5528 => conv_std_logic_vector(12, 8),
5529 => conv_std_logic_vector(12, 8),
5530 => conv_std_logic_vector(12, 8),
5531 => conv_std_logic_vector(12, 8),
5532 => conv_std_logic_vector(12, 8),
5533 => conv_std_logic_vector(12, 8),
5534 => conv_std_logic_vector(12, 8),
5535 => conv_std_logic_vector(13, 8),
5536 => conv_std_logic_vector(13, 8),
5537 => conv_std_logic_vector(13, 8),
5538 => conv_std_logic_vector(13, 8),
5539 => conv_std_logic_vector(13, 8),
5540 => conv_std_logic_vector(13, 8),
5541 => conv_std_logic_vector(13, 8),
5542 => conv_std_logic_vector(13, 8),
5543 => conv_std_logic_vector(13, 8),
5544 => conv_std_logic_vector(13, 8),
5545 => conv_std_logic_vector(13, 8),
5546 => conv_std_logic_vector(13, 8),
5547 => conv_std_logic_vector(14, 8),
5548 => conv_std_logic_vector(14, 8),
5549 => conv_std_logic_vector(14, 8),
5550 => conv_std_logic_vector(14, 8),
5551 => conv_std_logic_vector(14, 8),
5552 => conv_std_logic_vector(14, 8),
5553 => conv_std_logic_vector(14, 8),
5554 => conv_std_logic_vector(14, 8),
5555 => conv_std_logic_vector(14, 8),
5556 => conv_std_logic_vector(14, 8),
5557 => conv_std_logic_vector(14, 8),
5558 => conv_std_logic_vector(14, 8),
5559 => conv_std_logic_vector(15, 8),
5560 => conv_std_logic_vector(15, 8),
5561 => conv_std_logic_vector(15, 8),
5562 => conv_std_logic_vector(15, 8),
5563 => conv_std_logic_vector(15, 8),
5564 => conv_std_logic_vector(15, 8),
5565 => conv_std_logic_vector(15, 8),
5566 => conv_std_logic_vector(15, 8),
5567 => conv_std_logic_vector(15, 8),
5568 => conv_std_logic_vector(15, 8),
5569 => conv_std_logic_vector(15, 8),
5570 => conv_std_logic_vector(15, 8),
5571 => conv_std_logic_vector(15, 8),
5572 => conv_std_logic_vector(16, 8),
5573 => conv_std_logic_vector(16, 8),
5574 => conv_std_logic_vector(16, 8),
5575 => conv_std_logic_vector(16, 8),
5576 => conv_std_logic_vector(16, 8),
5577 => conv_std_logic_vector(16, 8),
5578 => conv_std_logic_vector(16, 8),
5579 => conv_std_logic_vector(16, 8),
5580 => conv_std_logic_vector(16, 8),
5581 => conv_std_logic_vector(16, 8),
5582 => conv_std_logic_vector(16, 8),
5583 => conv_std_logic_vector(16, 8),
5584 => conv_std_logic_vector(17, 8),
5585 => conv_std_logic_vector(17, 8),
5586 => conv_std_logic_vector(17, 8),
5587 => conv_std_logic_vector(17, 8),
5588 => conv_std_logic_vector(17, 8),
5589 => conv_std_logic_vector(17, 8),
5590 => conv_std_logic_vector(17, 8),
5591 => conv_std_logic_vector(17, 8),
5592 => conv_std_logic_vector(17, 8),
5593 => conv_std_logic_vector(17, 8),
5594 => conv_std_logic_vector(17, 8),
5595 => conv_std_logic_vector(17, 8),
5596 => conv_std_logic_vector(18, 8),
5597 => conv_std_logic_vector(18, 8),
5598 => conv_std_logic_vector(18, 8),
5599 => conv_std_logic_vector(18, 8),
5600 => conv_std_logic_vector(18, 8),
5601 => conv_std_logic_vector(18, 8),
5602 => conv_std_logic_vector(18, 8),
5603 => conv_std_logic_vector(18, 8),
5604 => conv_std_logic_vector(18, 8),
5605 => conv_std_logic_vector(18, 8),
5606 => conv_std_logic_vector(18, 8),
5607 => conv_std_logic_vector(18, 8),
5608 => conv_std_logic_vector(19, 8),
5609 => conv_std_logic_vector(19, 8),
5610 => conv_std_logic_vector(19, 8),
5611 => conv_std_logic_vector(19, 8),
5612 => conv_std_logic_vector(19, 8),
5613 => conv_std_logic_vector(19, 8),
5614 => conv_std_logic_vector(19, 8),
5615 => conv_std_logic_vector(19, 8),
5616 => conv_std_logic_vector(19, 8),
5617 => conv_std_logic_vector(19, 8),
5618 => conv_std_logic_vector(19, 8),
5619 => conv_std_logic_vector(19, 8),
5620 => conv_std_logic_vector(20, 8),
5621 => conv_std_logic_vector(20, 8),
5622 => conv_std_logic_vector(20, 8),
5623 => conv_std_logic_vector(20, 8),
5624 => conv_std_logic_vector(20, 8),
5625 => conv_std_logic_vector(20, 8),
5626 => conv_std_logic_vector(20, 8),
5627 => conv_std_logic_vector(20, 8),
5628 => conv_std_logic_vector(20, 8),
5629 => conv_std_logic_vector(20, 8),
5630 => conv_std_logic_vector(20, 8),
5631 => conv_std_logic_vector(20, 8),
5632 => conv_std_logic_vector(0, 8),
5633 => conv_std_logic_vector(0, 8),
5634 => conv_std_logic_vector(0, 8),
5635 => conv_std_logic_vector(0, 8),
5636 => conv_std_logic_vector(0, 8),
5637 => conv_std_logic_vector(0, 8),
5638 => conv_std_logic_vector(0, 8),
5639 => conv_std_logic_vector(0, 8),
5640 => conv_std_logic_vector(0, 8),
5641 => conv_std_logic_vector(0, 8),
5642 => conv_std_logic_vector(0, 8),
5643 => conv_std_logic_vector(0, 8),
5644 => conv_std_logic_vector(1, 8),
5645 => conv_std_logic_vector(1, 8),
5646 => conv_std_logic_vector(1, 8),
5647 => conv_std_logic_vector(1, 8),
5648 => conv_std_logic_vector(1, 8),
5649 => conv_std_logic_vector(1, 8),
5650 => conv_std_logic_vector(1, 8),
5651 => conv_std_logic_vector(1, 8),
5652 => conv_std_logic_vector(1, 8),
5653 => conv_std_logic_vector(1, 8),
5654 => conv_std_logic_vector(1, 8),
5655 => conv_std_logic_vector(1, 8),
5656 => conv_std_logic_vector(2, 8),
5657 => conv_std_logic_vector(2, 8),
5658 => conv_std_logic_vector(2, 8),
5659 => conv_std_logic_vector(2, 8),
5660 => conv_std_logic_vector(2, 8),
5661 => conv_std_logic_vector(2, 8),
5662 => conv_std_logic_vector(2, 8),
5663 => conv_std_logic_vector(2, 8),
5664 => conv_std_logic_vector(2, 8),
5665 => conv_std_logic_vector(2, 8),
5666 => conv_std_logic_vector(2, 8),
5667 => conv_std_logic_vector(3, 8),
5668 => conv_std_logic_vector(3, 8),
5669 => conv_std_logic_vector(3, 8),
5670 => conv_std_logic_vector(3, 8),
5671 => conv_std_logic_vector(3, 8),
5672 => conv_std_logic_vector(3, 8),
5673 => conv_std_logic_vector(3, 8),
5674 => conv_std_logic_vector(3, 8),
5675 => conv_std_logic_vector(3, 8),
5676 => conv_std_logic_vector(3, 8),
5677 => conv_std_logic_vector(3, 8),
5678 => conv_std_logic_vector(3, 8),
5679 => conv_std_logic_vector(4, 8),
5680 => conv_std_logic_vector(4, 8),
5681 => conv_std_logic_vector(4, 8),
5682 => conv_std_logic_vector(4, 8),
5683 => conv_std_logic_vector(4, 8),
5684 => conv_std_logic_vector(4, 8),
5685 => conv_std_logic_vector(4, 8),
5686 => conv_std_logic_vector(4, 8),
5687 => conv_std_logic_vector(4, 8),
5688 => conv_std_logic_vector(4, 8),
5689 => conv_std_logic_vector(4, 8),
5690 => conv_std_logic_vector(4, 8),
5691 => conv_std_logic_vector(5, 8),
5692 => conv_std_logic_vector(5, 8),
5693 => conv_std_logic_vector(5, 8),
5694 => conv_std_logic_vector(5, 8),
5695 => conv_std_logic_vector(5, 8),
5696 => conv_std_logic_vector(5, 8),
5697 => conv_std_logic_vector(5, 8),
5698 => conv_std_logic_vector(5, 8),
5699 => conv_std_logic_vector(5, 8),
5700 => conv_std_logic_vector(5, 8),
5701 => conv_std_logic_vector(5, 8),
5702 => conv_std_logic_vector(6, 8),
5703 => conv_std_logic_vector(6, 8),
5704 => conv_std_logic_vector(6, 8),
5705 => conv_std_logic_vector(6, 8),
5706 => conv_std_logic_vector(6, 8),
5707 => conv_std_logic_vector(6, 8),
5708 => conv_std_logic_vector(6, 8),
5709 => conv_std_logic_vector(6, 8),
5710 => conv_std_logic_vector(6, 8),
5711 => conv_std_logic_vector(6, 8),
5712 => conv_std_logic_vector(6, 8),
5713 => conv_std_logic_vector(6, 8),
5714 => conv_std_logic_vector(7, 8),
5715 => conv_std_logic_vector(7, 8),
5716 => conv_std_logic_vector(7, 8),
5717 => conv_std_logic_vector(7, 8),
5718 => conv_std_logic_vector(7, 8),
5719 => conv_std_logic_vector(7, 8),
5720 => conv_std_logic_vector(7, 8),
5721 => conv_std_logic_vector(7, 8),
5722 => conv_std_logic_vector(7, 8),
5723 => conv_std_logic_vector(7, 8),
5724 => conv_std_logic_vector(7, 8),
5725 => conv_std_logic_vector(7, 8),
5726 => conv_std_logic_vector(8, 8),
5727 => conv_std_logic_vector(8, 8),
5728 => conv_std_logic_vector(8, 8),
5729 => conv_std_logic_vector(8, 8),
5730 => conv_std_logic_vector(8, 8),
5731 => conv_std_logic_vector(8, 8),
5732 => conv_std_logic_vector(8, 8),
5733 => conv_std_logic_vector(8, 8),
5734 => conv_std_logic_vector(8, 8),
5735 => conv_std_logic_vector(8, 8),
5736 => conv_std_logic_vector(8, 8),
5737 => conv_std_logic_vector(9, 8),
5738 => conv_std_logic_vector(9, 8),
5739 => conv_std_logic_vector(9, 8),
5740 => conv_std_logic_vector(9, 8),
5741 => conv_std_logic_vector(9, 8),
5742 => conv_std_logic_vector(9, 8),
5743 => conv_std_logic_vector(9, 8),
5744 => conv_std_logic_vector(9, 8),
5745 => conv_std_logic_vector(9, 8),
5746 => conv_std_logic_vector(9, 8),
5747 => conv_std_logic_vector(9, 8),
5748 => conv_std_logic_vector(9, 8),
5749 => conv_std_logic_vector(10, 8),
5750 => conv_std_logic_vector(10, 8),
5751 => conv_std_logic_vector(10, 8),
5752 => conv_std_logic_vector(10, 8),
5753 => conv_std_logic_vector(10, 8),
5754 => conv_std_logic_vector(10, 8),
5755 => conv_std_logic_vector(10, 8),
5756 => conv_std_logic_vector(10, 8),
5757 => conv_std_logic_vector(10, 8),
5758 => conv_std_logic_vector(10, 8),
5759 => conv_std_logic_vector(10, 8),
5760 => conv_std_logic_vector(11, 8),
5761 => conv_std_logic_vector(11, 8),
5762 => conv_std_logic_vector(11, 8),
5763 => conv_std_logic_vector(11, 8),
5764 => conv_std_logic_vector(11, 8),
5765 => conv_std_logic_vector(11, 8),
5766 => conv_std_logic_vector(11, 8),
5767 => conv_std_logic_vector(11, 8),
5768 => conv_std_logic_vector(11, 8),
5769 => conv_std_logic_vector(11, 8),
5770 => conv_std_logic_vector(11, 8),
5771 => conv_std_logic_vector(11, 8),
5772 => conv_std_logic_vector(12, 8),
5773 => conv_std_logic_vector(12, 8),
5774 => conv_std_logic_vector(12, 8),
5775 => conv_std_logic_vector(12, 8),
5776 => conv_std_logic_vector(12, 8),
5777 => conv_std_logic_vector(12, 8),
5778 => conv_std_logic_vector(12, 8),
5779 => conv_std_logic_vector(12, 8),
5780 => conv_std_logic_vector(12, 8),
5781 => conv_std_logic_vector(12, 8),
5782 => conv_std_logic_vector(12, 8),
5783 => conv_std_logic_vector(12, 8),
5784 => conv_std_logic_vector(13, 8),
5785 => conv_std_logic_vector(13, 8),
5786 => conv_std_logic_vector(13, 8),
5787 => conv_std_logic_vector(13, 8),
5788 => conv_std_logic_vector(13, 8),
5789 => conv_std_logic_vector(13, 8),
5790 => conv_std_logic_vector(13, 8),
5791 => conv_std_logic_vector(13, 8),
5792 => conv_std_logic_vector(13, 8),
5793 => conv_std_logic_vector(13, 8),
5794 => conv_std_logic_vector(13, 8),
5795 => conv_std_logic_vector(14, 8),
5796 => conv_std_logic_vector(14, 8),
5797 => conv_std_logic_vector(14, 8),
5798 => conv_std_logic_vector(14, 8),
5799 => conv_std_logic_vector(14, 8),
5800 => conv_std_logic_vector(14, 8),
5801 => conv_std_logic_vector(14, 8),
5802 => conv_std_logic_vector(14, 8),
5803 => conv_std_logic_vector(14, 8),
5804 => conv_std_logic_vector(14, 8),
5805 => conv_std_logic_vector(14, 8),
5806 => conv_std_logic_vector(14, 8),
5807 => conv_std_logic_vector(15, 8),
5808 => conv_std_logic_vector(15, 8),
5809 => conv_std_logic_vector(15, 8),
5810 => conv_std_logic_vector(15, 8),
5811 => conv_std_logic_vector(15, 8),
5812 => conv_std_logic_vector(15, 8),
5813 => conv_std_logic_vector(15, 8),
5814 => conv_std_logic_vector(15, 8),
5815 => conv_std_logic_vector(15, 8),
5816 => conv_std_logic_vector(15, 8),
5817 => conv_std_logic_vector(15, 8),
5818 => conv_std_logic_vector(15, 8),
5819 => conv_std_logic_vector(16, 8),
5820 => conv_std_logic_vector(16, 8),
5821 => conv_std_logic_vector(16, 8),
5822 => conv_std_logic_vector(16, 8),
5823 => conv_std_logic_vector(16, 8),
5824 => conv_std_logic_vector(16, 8),
5825 => conv_std_logic_vector(16, 8),
5826 => conv_std_logic_vector(16, 8),
5827 => conv_std_logic_vector(16, 8),
5828 => conv_std_logic_vector(16, 8),
5829 => conv_std_logic_vector(16, 8),
5830 => conv_std_logic_vector(17, 8),
5831 => conv_std_logic_vector(17, 8),
5832 => conv_std_logic_vector(17, 8),
5833 => conv_std_logic_vector(17, 8),
5834 => conv_std_logic_vector(17, 8),
5835 => conv_std_logic_vector(17, 8),
5836 => conv_std_logic_vector(17, 8),
5837 => conv_std_logic_vector(17, 8),
5838 => conv_std_logic_vector(17, 8),
5839 => conv_std_logic_vector(17, 8),
5840 => conv_std_logic_vector(17, 8),
5841 => conv_std_logic_vector(17, 8),
5842 => conv_std_logic_vector(18, 8),
5843 => conv_std_logic_vector(18, 8),
5844 => conv_std_logic_vector(18, 8),
5845 => conv_std_logic_vector(18, 8),
5846 => conv_std_logic_vector(18, 8),
5847 => conv_std_logic_vector(18, 8),
5848 => conv_std_logic_vector(18, 8),
5849 => conv_std_logic_vector(18, 8),
5850 => conv_std_logic_vector(18, 8),
5851 => conv_std_logic_vector(18, 8),
5852 => conv_std_logic_vector(18, 8),
5853 => conv_std_logic_vector(18, 8),
5854 => conv_std_logic_vector(19, 8),
5855 => conv_std_logic_vector(19, 8),
5856 => conv_std_logic_vector(19, 8),
5857 => conv_std_logic_vector(19, 8),
5858 => conv_std_logic_vector(19, 8),
5859 => conv_std_logic_vector(19, 8),
5860 => conv_std_logic_vector(19, 8),
5861 => conv_std_logic_vector(19, 8),
5862 => conv_std_logic_vector(19, 8),
5863 => conv_std_logic_vector(19, 8),
5864 => conv_std_logic_vector(19, 8),
5865 => conv_std_logic_vector(20, 8),
5866 => conv_std_logic_vector(20, 8),
5867 => conv_std_logic_vector(20, 8),
5868 => conv_std_logic_vector(20, 8),
5869 => conv_std_logic_vector(20, 8),
5870 => conv_std_logic_vector(20, 8),
5871 => conv_std_logic_vector(20, 8),
5872 => conv_std_logic_vector(20, 8),
5873 => conv_std_logic_vector(20, 8),
5874 => conv_std_logic_vector(20, 8),
5875 => conv_std_logic_vector(20, 8),
5876 => conv_std_logic_vector(20, 8),
5877 => conv_std_logic_vector(21, 8),
5878 => conv_std_logic_vector(21, 8),
5879 => conv_std_logic_vector(21, 8),
5880 => conv_std_logic_vector(21, 8),
5881 => conv_std_logic_vector(21, 8),
5882 => conv_std_logic_vector(21, 8),
5883 => conv_std_logic_vector(21, 8),
5884 => conv_std_logic_vector(21, 8),
5885 => conv_std_logic_vector(21, 8),
5886 => conv_std_logic_vector(21, 8),
5887 => conv_std_logic_vector(21, 8),
5888 => conv_std_logic_vector(0, 8),
5889 => conv_std_logic_vector(0, 8),
5890 => conv_std_logic_vector(0, 8),
5891 => conv_std_logic_vector(0, 8),
5892 => conv_std_logic_vector(0, 8),
5893 => conv_std_logic_vector(0, 8),
5894 => conv_std_logic_vector(0, 8),
5895 => conv_std_logic_vector(0, 8),
5896 => conv_std_logic_vector(0, 8),
5897 => conv_std_logic_vector(0, 8),
5898 => conv_std_logic_vector(0, 8),
5899 => conv_std_logic_vector(0, 8),
5900 => conv_std_logic_vector(1, 8),
5901 => conv_std_logic_vector(1, 8),
5902 => conv_std_logic_vector(1, 8),
5903 => conv_std_logic_vector(1, 8),
5904 => conv_std_logic_vector(1, 8),
5905 => conv_std_logic_vector(1, 8),
5906 => conv_std_logic_vector(1, 8),
5907 => conv_std_logic_vector(1, 8),
5908 => conv_std_logic_vector(1, 8),
5909 => conv_std_logic_vector(1, 8),
5910 => conv_std_logic_vector(1, 8),
5911 => conv_std_logic_vector(2, 8),
5912 => conv_std_logic_vector(2, 8),
5913 => conv_std_logic_vector(2, 8),
5914 => conv_std_logic_vector(2, 8),
5915 => conv_std_logic_vector(2, 8),
5916 => conv_std_logic_vector(2, 8),
5917 => conv_std_logic_vector(2, 8),
5918 => conv_std_logic_vector(2, 8),
5919 => conv_std_logic_vector(2, 8),
5920 => conv_std_logic_vector(2, 8),
5921 => conv_std_logic_vector(2, 8),
5922 => conv_std_logic_vector(3, 8),
5923 => conv_std_logic_vector(3, 8),
5924 => conv_std_logic_vector(3, 8),
5925 => conv_std_logic_vector(3, 8),
5926 => conv_std_logic_vector(3, 8),
5927 => conv_std_logic_vector(3, 8),
5928 => conv_std_logic_vector(3, 8),
5929 => conv_std_logic_vector(3, 8),
5930 => conv_std_logic_vector(3, 8),
5931 => conv_std_logic_vector(3, 8),
5932 => conv_std_logic_vector(3, 8),
5933 => conv_std_logic_vector(4, 8),
5934 => conv_std_logic_vector(4, 8),
5935 => conv_std_logic_vector(4, 8),
5936 => conv_std_logic_vector(4, 8),
5937 => conv_std_logic_vector(4, 8),
5938 => conv_std_logic_vector(4, 8),
5939 => conv_std_logic_vector(4, 8),
5940 => conv_std_logic_vector(4, 8),
5941 => conv_std_logic_vector(4, 8),
5942 => conv_std_logic_vector(4, 8),
5943 => conv_std_logic_vector(4, 8),
5944 => conv_std_logic_vector(5, 8),
5945 => conv_std_logic_vector(5, 8),
5946 => conv_std_logic_vector(5, 8),
5947 => conv_std_logic_vector(5, 8),
5948 => conv_std_logic_vector(5, 8),
5949 => conv_std_logic_vector(5, 8),
5950 => conv_std_logic_vector(5, 8),
5951 => conv_std_logic_vector(5, 8),
5952 => conv_std_logic_vector(5, 8),
5953 => conv_std_logic_vector(5, 8),
5954 => conv_std_logic_vector(5, 8),
5955 => conv_std_logic_vector(6, 8),
5956 => conv_std_logic_vector(6, 8),
5957 => conv_std_logic_vector(6, 8),
5958 => conv_std_logic_vector(6, 8),
5959 => conv_std_logic_vector(6, 8),
5960 => conv_std_logic_vector(6, 8),
5961 => conv_std_logic_vector(6, 8),
5962 => conv_std_logic_vector(6, 8),
5963 => conv_std_logic_vector(6, 8),
5964 => conv_std_logic_vector(6, 8),
5965 => conv_std_logic_vector(6, 8),
5966 => conv_std_logic_vector(7, 8),
5967 => conv_std_logic_vector(7, 8),
5968 => conv_std_logic_vector(7, 8),
5969 => conv_std_logic_vector(7, 8),
5970 => conv_std_logic_vector(7, 8),
5971 => conv_std_logic_vector(7, 8),
5972 => conv_std_logic_vector(7, 8),
5973 => conv_std_logic_vector(7, 8),
5974 => conv_std_logic_vector(7, 8),
5975 => conv_std_logic_vector(7, 8),
5976 => conv_std_logic_vector(7, 8),
5977 => conv_std_logic_vector(7, 8),
5978 => conv_std_logic_vector(8, 8),
5979 => conv_std_logic_vector(8, 8),
5980 => conv_std_logic_vector(8, 8),
5981 => conv_std_logic_vector(8, 8),
5982 => conv_std_logic_vector(8, 8),
5983 => conv_std_logic_vector(8, 8),
5984 => conv_std_logic_vector(8, 8),
5985 => conv_std_logic_vector(8, 8),
5986 => conv_std_logic_vector(8, 8),
5987 => conv_std_logic_vector(8, 8),
5988 => conv_std_logic_vector(8, 8),
5989 => conv_std_logic_vector(9, 8),
5990 => conv_std_logic_vector(9, 8),
5991 => conv_std_logic_vector(9, 8),
5992 => conv_std_logic_vector(9, 8),
5993 => conv_std_logic_vector(9, 8),
5994 => conv_std_logic_vector(9, 8),
5995 => conv_std_logic_vector(9, 8),
5996 => conv_std_logic_vector(9, 8),
5997 => conv_std_logic_vector(9, 8),
5998 => conv_std_logic_vector(9, 8),
5999 => conv_std_logic_vector(9, 8),
6000 => conv_std_logic_vector(10, 8),
6001 => conv_std_logic_vector(10, 8),
6002 => conv_std_logic_vector(10, 8),
6003 => conv_std_logic_vector(10, 8),
6004 => conv_std_logic_vector(10, 8),
6005 => conv_std_logic_vector(10, 8),
6006 => conv_std_logic_vector(10, 8),
6007 => conv_std_logic_vector(10, 8),
6008 => conv_std_logic_vector(10, 8),
6009 => conv_std_logic_vector(10, 8),
6010 => conv_std_logic_vector(10, 8),
6011 => conv_std_logic_vector(11, 8),
6012 => conv_std_logic_vector(11, 8),
6013 => conv_std_logic_vector(11, 8),
6014 => conv_std_logic_vector(11, 8),
6015 => conv_std_logic_vector(11, 8),
6016 => conv_std_logic_vector(11, 8),
6017 => conv_std_logic_vector(11, 8),
6018 => conv_std_logic_vector(11, 8),
6019 => conv_std_logic_vector(11, 8),
6020 => conv_std_logic_vector(11, 8),
6021 => conv_std_logic_vector(11, 8),
6022 => conv_std_logic_vector(12, 8),
6023 => conv_std_logic_vector(12, 8),
6024 => conv_std_logic_vector(12, 8),
6025 => conv_std_logic_vector(12, 8),
6026 => conv_std_logic_vector(12, 8),
6027 => conv_std_logic_vector(12, 8),
6028 => conv_std_logic_vector(12, 8),
6029 => conv_std_logic_vector(12, 8),
6030 => conv_std_logic_vector(12, 8),
6031 => conv_std_logic_vector(12, 8),
6032 => conv_std_logic_vector(12, 8),
6033 => conv_std_logic_vector(13, 8),
6034 => conv_std_logic_vector(13, 8),
6035 => conv_std_logic_vector(13, 8),
6036 => conv_std_logic_vector(13, 8),
6037 => conv_std_logic_vector(13, 8),
6038 => conv_std_logic_vector(13, 8),
6039 => conv_std_logic_vector(13, 8),
6040 => conv_std_logic_vector(13, 8),
6041 => conv_std_logic_vector(13, 8),
6042 => conv_std_logic_vector(13, 8),
6043 => conv_std_logic_vector(13, 8),
6044 => conv_std_logic_vector(14, 8),
6045 => conv_std_logic_vector(14, 8),
6046 => conv_std_logic_vector(14, 8),
6047 => conv_std_logic_vector(14, 8),
6048 => conv_std_logic_vector(14, 8),
6049 => conv_std_logic_vector(14, 8),
6050 => conv_std_logic_vector(14, 8),
6051 => conv_std_logic_vector(14, 8),
6052 => conv_std_logic_vector(14, 8),
6053 => conv_std_logic_vector(14, 8),
6054 => conv_std_logic_vector(14, 8),
6055 => conv_std_logic_vector(15, 8),
6056 => conv_std_logic_vector(15, 8),
6057 => conv_std_logic_vector(15, 8),
6058 => conv_std_logic_vector(15, 8),
6059 => conv_std_logic_vector(15, 8),
6060 => conv_std_logic_vector(15, 8),
6061 => conv_std_logic_vector(15, 8),
6062 => conv_std_logic_vector(15, 8),
6063 => conv_std_logic_vector(15, 8),
6064 => conv_std_logic_vector(15, 8),
6065 => conv_std_logic_vector(15, 8),
6066 => conv_std_logic_vector(15, 8),
6067 => conv_std_logic_vector(16, 8),
6068 => conv_std_logic_vector(16, 8),
6069 => conv_std_logic_vector(16, 8),
6070 => conv_std_logic_vector(16, 8),
6071 => conv_std_logic_vector(16, 8),
6072 => conv_std_logic_vector(16, 8),
6073 => conv_std_logic_vector(16, 8),
6074 => conv_std_logic_vector(16, 8),
6075 => conv_std_logic_vector(16, 8),
6076 => conv_std_logic_vector(16, 8),
6077 => conv_std_logic_vector(16, 8),
6078 => conv_std_logic_vector(17, 8),
6079 => conv_std_logic_vector(17, 8),
6080 => conv_std_logic_vector(17, 8),
6081 => conv_std_logic_vector(17, 8),
6082 => conv_std_logic_vector(17, 8),
6083 => conv_std_logic_vector(17, 8),
6084 => conv_std_logic_vector(17, 8),
6085 => conv_std_logic_vector(17, 8),
6086 => conv_std_logic_vector(17, 8),
6087 => conv_std_logic_vector(17, 8),
6088 => conv_std_logic_vector(17, 8),
6089 => conv_std_logic_vector(18, 8),
6090 => conv_std_logic_vector(18, 8),
6091 => conv_std_logic_vector(18, 8),
6092 => conv_std_logic_vector(18, 8),
6093 => conv_std_logic_vector(18, 8),
6094 => conv_std_logic_vector(18, 8),
6095 => conv_std_logic_vector(18, 8),
6096 => conv_std_logic_vector(18, 8),
6097 => conv_std_logic_vector(18, 8),
6098 => conv_std_logic_vector(18, 8),
6099 => conv_std_logic_vector(18, 8),
6100 => conv_std_logic_vector(19, 8),
6101 => conv_std_logic_vector(19, 8),
6102 => conv_std_logic_vector(19, 8),
6103 => conv_std_logic_vector(19, 8),
6104 => conv_std_logic_vector(19, 8),
6105 => conv_std_logic_vector(19, 8),
6106 => conv_std_logic_vector(19, 8),
6107 => conv_std_logic_vector(19, 8),
6108 => conv_std_logic_vector(19, 8),
6109 => conv_std_logic_vector(19, 8),
6110 => conv_std_logic_vector(19, 8),
6111 => conv_std_logic_vector(20, 8),
6112 => conv_std_logic_vector(20, 8),
6113 => conv_std_logic_vector(20, 8),
6114 => conv_std_logic_vector(20, 8),
6115 => conv_std_logic_vector(20, 8),
6116 => conv_std_logic_vector(20, 8),
6117 => conv_std_logic_vector(20, 8),
6118 => conv_std_logic_vector(20, 8),
6119 => conv_std_logic_vector(20, 8),
6120 => conv_std_logic_vector(20, 8),
6121 => conv_std_logic_vector(20, 8),
6122 => conv_std_logic_vector(21, 8),
6123 => conv_std_logic_vector(21, 8),
6124 => conv_std_logic_vector(21, 8),
6125 => conv_std_logic_vector(21, 8),
6126 => conv_std_logic_vector(21, 8),
6127 => conv_std_logic_vector(21, 8),
6128 => conv_std_logic_vector(21, 8),
6129 => conv_std_logic_vector(21, 8),
6130 => conv_std_logic_vector(21, 8),
6131 => conv_std_logic_vector(21, 8),
6132 => conv_std_logic_vector(21, 8),
6133 => conv_std_logic_vector(22, 8),
6134 => conv_std_logic_vector(22, 8),
6135 => conv_std_logic_vector(22, 8),
6136 => conv_std_logic_vector(22, 8),
6137 => conv_std_logic_vector(22, 8),
6138 => conv_std_logic_vector(22, 8),
6139 => conv_std_logic_vector(22, 8),
6140 => conv_std_logic_vector(22, 8),
6141 => conv_std_logic_vector(22, 8),
6142 => conv_std_logic_vector(22, 8),
6143 => conv_std_logic_vector(22, 8),
6144 => conv_std_logic_vector(0, 8),
6145 => conv_std_logic_vector(0, 8),
6146 => conv_std_logic_vector(0, 8),
6147 => conv_std_logic_vector(0, 8),
6148 => conv_std_logic_vector(0, 8),
6149 => conv_std_logic_vector(0, 8),
6150 => conv_std_logic_vector(0, 8),
6151 => conv_std_logic_vector(0, 8),
6152 => conv_std_logic_vector(0, 8),
6153 => conv_std_logic_vector(0, 8),
6154 => conv_std_logic_vector(0, 8),
6155 => conv_std_logic_vector(1, 8),
6156 => conv_std_logic_vector(1, 8),
6157 => conv_std_logic_vector(1, 8),
6158 => conv_std_logic_vector(1, 8),
6159 => conv_std_logic_vector(1, 8),
6160 => conv_std_logic_vector(1, 8),
6161 => conv_std_logic_vector(1, 8),
6162 => conv_std_logic_vector(1, 8),
6163 => conv_std_logic_vector(1, 8),
6164 => conv_std_logic_vector(1, 8),
6165 => conv_std_logic_vector(1, 8),
6166 => conv_std_logic_vector(2, 8),
6167 => conv_std_logic_vector(2, 8),
6168 => conv_std_logic_vector(2, 8),
6169 => conv_std_logic_vector(2, 8),
6170 => conv_std_logic_vector(2, 8),
6171 => conv_std_logic_vector(2, 8),
6172 => conv_std_logic_vector(2, 8),
6173 => conv_std_logic_vector(2, 8),
6174 => conv_std_logic_vector(2, 8),
6175 => conv_std_logic_vector(2, 8),
6176 => conv_std_logic_vector(3, 8),
6177 => conv_std_logic_vector(3, 8),
6178 => conv_std_logic_vector(3, 8),
6179 => conv_std_logic_vector(3, 8),
6180 => conv_std_logic_vector(3, 8),
6181 => conv_std_logic_vector(3, 8),
6182 => conv_std_logic_vector(3, 8),
6183 => conv_std_logic_vector(3, 8),
6184 => conv_std_logic_vector(3, 8),
6185 => conv_std_logic_vector(3, 8),
6186 => conv_std_logic_vector(3, 8),
6187 => conv_std_logic_vector(4, 8),
6188 => conv_std_logic_vector(4, 8),
6189 => conv_std_logic_vector(4, 8),
6190 => conv_std_logic_vector(4, 8),
6191 => conv_std_logic_vector(4, 8),
6192 => conv_std_logic_vector(4, 8),
6193 => conv_std_logic_vector(4, 8),
6194 => conv_std_logic_vector(4, 8),
6195 => conv_std_logic_vector(4, 8),
6196 => conv_std_logic_vector(4, 8),
6197 => conv_std_logic_vector(4, 8),
6198 => conv_std_logic_vector(5, 8),
6199 => conv_std_logic_vector(5, 8),
6200 => conv_std_logic_vector(5, 8),
6201 => conv_std_logic_vector(5, 8),
6202 => conv_std_logic_vector(5, 8),
6203 => conv_std_logic_vector(5, 8),
6204 => conv_std_logic_vector(5, 8),
6205 => conv_std_logic_vector(5, 8),
6206 => conv_std_logic_vector(5, 8),
6207 => conv_std_logic_vector(5, 8),
6208 => conv_std_logic_vector(6, 8),
6209 => conv_std_logic_vector(6, 8),
6210 => conv_std_logic_vector(6, 8),
6211 => conv_std_logic_vector(6, 8),
6212 => conv_std_logic_vector(6, 8),
6213 => conv_std_logic_vector(6, 8),
6214 => conv_std_logic_vector(6, 8),
6215 => conv_std_logic_vector(6, 8),
6216 => conv_std_logic_vector(6, 8),
6217 => conv_std_logic_vector(6, 8),
6218 => conv_std_logic_vector(6, 8),
6219 => conv_std_logic_vector(7, 8),
6220 => conv_std_logic_vector(7, 8),
6221 => conv_std_logic_vector(7, 8),
6222 => conv_std_logic_vector(7, 8),
6223 => conv_std_logic_vector(7, 8),
6224 => conv_std_logic_vector(7, 8),
6225 => conv_std_logic_vector(7, 8),
6226 => conv_std_logic_vector(7, 8),
6227 => conv_std_logic_vector(7, 8),
6228 => conv_std_logic_vector(7, 8),
6229 => conv_std_logic_vector(7, 8),
6230 => conv_std_logic_vector(8, 8),
6231 => conv_std_logic_vector(8, 8),
6232 => conv_std_logic_vector(8, 8),
6233 => conv_std_logic_vector(8, 8),
6234 => conv_std_logic_vector(8, 8),
6235 => conv_std_logic_vector(8, 8),
6236 => conv_std_logic_vector(8, 8),
6237 => conv_std_logic_vector(8, 8),
6238 => conv_std_logic_vector(8, 8),
6239 => conv_std_logic_vector(8, 8),
6240 => conv_std_logic_vector(9, 8),
6241 => conv_std_logic_vector(9, 8),
6242 => conv_std_logic_vector(9, 8),
6243 => conv_std_logic_vector(9, 8),
6244 => conv_std_logic_vector(9, 8),
6245 => conv_std_logic_vector(9, 8),
6246 => conv_std_logic_vector(9, 8),
6247 => conv_std_logic_vector(9, 8),
6248 => conv_std_logic_vector(9, 8),
6249 => conv_std_logic_vector(9, 8),
6250 => conv_std_logic_vector(9, 8),
6251 => conv_std_logic_vector(10, 8),
6252 => conv_std_logic_vector(10, 8),
6253 => conv_std_logic_vector(10, 8),
6254 => conv_std_logic_vector(10, 8),
6255 => conv_std_logic_vector(10, 8),
6256 => conv_std_logic_vector(10, 8),
6257 => conv_std_logic_vector(10, 8),
6258 => conv_std_logic_vector(10, 8),
6259 => conv_std_logic_vector(10, 8),
6260 => conv_std_logic_vector(10, 8),
6261 => conv_std_logic_vector(10, 8),
6262 => conv_std_logic_vector(11, 8),
6263 => conv_std_logic_vector(11, 8),
6264 => conv_std_logic_vector(11, 8),
6265 => conv_std_logic_vector(11, 8),
6266 => conv_std_logic_vector(11, 8),
6267 => conv_std_logic_vector(11, 8),
6268 => conv_std_logic_vector(11, 8),
6269 => conv_std_logic_vector(11, 8),
6270 => conv_std_logic_vector(11, 8),
6271 => conv_std_logic_vector(11, 8),
6272 => conv_std_logic_vector(12, 8),
6273 => conv_std_logic_vector(12, 8),
6274 => conv_std_logic_vector(12, 8),
6275 => conv_std_logic_vector(12, 8),
6276 => conv_std_logic_vector(12, 8),
6277 => conv_std_logic_vector(12, 8),
6278 => conv_std_logic_vector(12, 8),
6279 => conv_std_logic_vector(12, 8),
6280 => conv_std_logic_vector(12, 8),
6281 => conv_std_logic_vector(12, 8),
6282 => conv_std_logic_vector(12, 8),
6283 => conv_std_logic_vector(13, 8),
6284 => conv_std_logic_vector(13, 8),
6285 => conv_std_logic_vector(13, 8),
6286 => conv_std_logic_vector(13, 8),
6287 => conv_std_logic_vector(13, 8),
6288 => conv_std_logic_vector(13, 8),
6289 => conv_std_logic_vector(13, 8),
6290 => conv_std_logic_vector(13, 8),
6291 => conv_std_logic_vector(13, 8),
6292 => conv_std_logic_vector(13, 8),
6293 => conv_std_logic_vector(13, 8),
6294 => conv_std_logic_vector(14, 8),
6295 => conv_std_logic_vector(14, 8),
6296 => conv_std_logic_vector(14, 8),
6297 => conv_std_logic_vector(14, 8),
6298 => conv_std_logic_vector(14, 8),
6299 => conv_std_logic_vector(14, 8),
6300 => conv_std_logic_vector(14, 8),
6301 => conv_std_logic_vector(14, 8),
6302 => conv_std_logic_vector(14, 8),
6303 => conv_std_logic_vector(14, 8),
6304 => conv_std_logic_vector(15, 8),
6305 => conv_std_logic_vector(15, 8),
6306 => conv_std_logic_vector(15, 8),
6307 => conv_std_logic_vector(15, 8),
6308 => conv_std_logic_vector(15, 8),
6309 => conv_std_logic_vector(15, 8),
6310 => conv_std_logic_vector(15, 8),
6311 => conv_std_logic_vector(15, 8),
6312 => conv_std_logic_vector(15, 8),
6313 => conv_std_logic_vector(15, 8),
6314 => conv_std_logic_vector(15, 8),
6315 => conv_std_logic_vector(16, 8),
6316 => conv_std_logic_vector(16, 8),
6317 => conv_std_logic_vector(16, 8),
6318 => conv_std_logic_vector(16, 8),
6319 => conv_std_logic_vector(16, 8),
6320 => conv_std_logic_vector(16, 8),
6321 => conv_std_logic_vector(16, 8),
6322 => conv_std_logic_vector(16, 8),
6323 => conv_std_logic_vector(16, 8),
6324 => conv_std_logic_vector(16, 8),
6325 => conv_std_logic_vector(16, 8),
6326 => conv_std_logic_vector(17, 8),
6327 => conv_std_logic_vector(17, 8),
6328 => conv_std_logic_vector(17, 8),
6329 => conv_std_logic_vector(17, 8),
6330 => conv_std_logic_vector(17, 8),
6331 => conv_std_logic_vector(17, 8),
6332 => conv_std_logic_vector(17, 8),
6333 => conv_std_logic_vector(17, 8),
6334 => conv_std_logic_vector(17, 8),
6335 => conv_std_logic_vector(17, 8),
6336 => conv_std_logic_vector(18, 8),
6337 => conv_std_logic_vector(18, 8),
6338 => conv_std_logic_vector(18, 8),
6339 => conv_std_logic_vector(18, 8),
6340 => conv_std_logic_vector(18, 8),
6341 => conv_std_logic_vector(18, 8),
6342 => conv_std_logic_vector(18, 8),
6343 => conv_std_logic_vector(18, 8),
6344 => conv_std_logic_vector(18, 8),
6345 => conv_std_logic_vector(18, 8),
6346 => conv_std_logic_vector(18, 8),
6347 => conv_std_logic_vector(19, 8),
6348 => conv_std_logic_vector(19, 8),
6349 => conv_std_logic_vector(19, 8),
6350 => conv_std_logic_vector(19, 8),
6351 => conv_std_logic_vector(19, 8),
6352 => conv_std_logic_vector(19, 8),
6353 => conv_std_logic_vector(19, 8),
6354 => conv_std_logic_vector(19, 8),
6355 => conv_std_logic_vector(19, 8),
6356 => conv_std_logic_vector(19, 8),
6357 => conv_std_logic_vector(19, 8),
6358 => conv_std_logic_vector(20, 8),
6359 => conv_std_logic_vector(20, 8),
6360 => conv_std_logic_vector(20, 8),
6361 => conv_std_logic_vector(20, 8),
6362 => conv_std_logic_vector(20, 8),
6363 => conv_std_logic_vector(20, 8),
6364 => conv_std_logic_vector(20, 8),
6365 => conv_std_logic_vector(20, 8),
6366 => conv_std_logic_vector(20, 8),
6367 => conv_std_logic_vector(20, 8),
6368 => conv_std_logic_vector(21, 8),
6369 => conv_std_logic_vector(21, 8),
6370 => conv_std_logic_vector(21, 8),
6371 => conv_std_logic_vector(21, 8),
6372 => conv_std_logic_vector(21, 8),
6373 => conv_std_logic_vector(21, 8),
6374 => conv_std_logic_vector(21, 8),
6375 => conv_std_logic_vector(21, 8),
6376 => conv_std_logic_vector(21, 8),
6377 => conv_std_logic_vector(21, 8),
6378 => conv_std_logic_vector(21, 8),
6379 => conv_std_logic_vector(22, 8),
6380 => conv_std_logic_vector(22, 8),
6381 => conv_std_logic_vector(22, 8),
6382 => conv_std_logic_vector(22, 8),
6383 => conv_std_logic_vector(22, 8),
6384 => conv_std_logic_vector(22, 8),
6385 => conv_std_logic_vector(22, 8),
6386 => conv_std_logic_vector(22, 8),
6387 => conv_std_logic_vector(22, 8),
6388 => conv_std_logic_vector(22, 8),
6389 => conv_std_logic_vector(22, 8),
6390 => conv_std_logic_vector(23, 8),
6391 => conv_std_logic_vector(23, 8),
6392 => conv_std_logic_vector(23, 8),
6393 => conv_std_logic_vector(23, 8),
6394 => conv_std_logic_vector(23, 8),
6395 => conv_std_logic_vector(23, 8),
6396 => conv_std_logic_vector(23, 8),
6397 => conv_std_logic_vector(23, 8),
6398 => conv_std_logic_vector(23, 8),
6399 => conv_std_logic_vector(23, 8),
6400 => conv_std_logic_vector(0, 8),
6401 => conv_std_logic_vector(0, 8),
6402 => conv_std_logic_vector(0, 8),
6403 => conv_std_logic_vector(0, 8),
6404 => conv_std_logic_vector(0, 8),
6405 => conv_std_logic_vector(0, 8),
6406 => conv_std_logic_vector(0, 8),
6407 => conv_std_logic_vector(0, 8),
6408 => conv_std_logic_vector(0, 8),
6409 => conv_std_logic_vector(0, 8),
6410 => conv_std_logic_vector(0, 8),
6411 => conv_std_logic_vector(1, 8),
6412 => conv_std_logic_vector(1, 8),
6413 => conv_std_logic_vector(1, 8),
6414 => conv_std_logic_vector(1, 8),
6415 => conv_std_logic_vector(1, 8),
6416 => conv_std_logic_vector(1, 8),
6417 => conv_std_logic_vector(1, 8),
6418 => conv_std_logic_vector(1, 8),
6419 => conv_std_logic_vector(1, 8),
6420 => conv_std_logic_vector(1, 8),
6421 => conv_std_logic_vector(2, 8),
6422 => conv_std_logic_vector(2, 8),
6423 => conv_std_logic_vector(2, 8),
6424 => conv_std_logic_vector(2, 8),
6425 => conv_std_logic_vector(2, 8),
6426 => conv_std_logic_vector(2, 8),
6427 => conv_std_logic_vector(2, 8),
6428 => conv_std_logic_vector(2, 8),
6429 => conv_std_logic_vector(2, 8),
6430 => conv_std_logic_vector(2, 8),
6431 => conv_std_logic_vector(3, 8),
6432 => conv_std_logic_vector(3, 8),
6433 => conv_std_logic_vector(3, 8),
6434 => conv_std_logic_vector(3, 8),
6435 => conv_std_logic_vector(3, 8),
6436 => conv_std_logic_vector(3, 8),
6437 => conv_std_logic_vector(3, 8),
6438 => conv_std_logic_vector(3, 8),
6439 => conv_std_logic_vector(3, 8),
6440 => conv_std_logic_vector(3, 8),
6441 => conv_std_logic_vector(4, 8),
6442 => conv_std_logic_vector(4, 8),
6443 => conv_std_logic_vector(4, 8),
6444 => conv_std_logic_vector(4, 8),
6445 => conv_std_logic_vector(4, 8),
6446 => conv_std_logic_vector(4, 8),
6447 => conv_std_logic_vector(4, 8),
6448 => conv_std_logic_vector(4, 8),
6449 => conv_std_logic_vector(4, 8),
6450 => conv_std_logic_vector(4, 8),
6451 => conv_std_logic_vector(4, 8),
6452 => conv_std_logic_vector(5, 8),
6453 => conv_std_logic_vector(5, 8),
6454 => conv_std_logic_vector(5, 8),
6455 => conv_std_logic_vector(5, 8),
6456 => conv_std_logic_vector(5, 8),
6457 => conv_std_logic_vector(5, 8),
6458 => conv_std_logic_vector(5, 8),
6459 => conv_std_logic_vector(5, 8),
6460 => conv_std_logic_vector(5, 8),
6461 => conv_std_logic_vector(5, 8),
6462 => conv_std_logic_vector(6, 8),
6463 => conv_std_logic_vector(6, 8),
6464 => conv_std_logic_vector(6, 8),
6465 => conv_std_logic_vector(6, 8),
6466 => conv_std_logic_vector(6, 8),
6467 => conv_std_logic_vector(6, 8),
6468 => conv_std_logic_vector(6, 8),
6469 => conv_std_logic_vector(6, 8),
6470 => conv_std_logic_vector(6, 8),
6471 => conv_std_logic_vector(6, 8),
6472 => conv_std_logic_vector(7, 8),
6473 => conv_std_logic_vector(7, 8),
6474 => conv_std_logic_vector(7, 8),
6475 => conv_std_logic_vector(7, 8),
6476 => conv_std_logic_vector(7, 8),
6477 => conv_std_logic_vector(7, 8),
6478 => conv_std_logic_vector(7, 8),
6479 => conv_std_logic_vector(7, 8),
6480 => conv_std_logic_vector(7, 8),
6481 => conv_std_logic_vector(7, 8),
6482 => conv_std_logic_vector(8, 8),
6483 => conv_std_logic_vector(8, 8),
6484 => conv_std_logic_vector(8, 8),
6485 => conv_std_logic_vector(8, 8),
6486 => conv_std_logic_vector(8, 8),
6487 => conv_std_logic_vector(8, 8),
6488 => conv_std_logic_vector(8, 8),
6489 => conv_std_logic_vector(8, 8),
6490 => conv_std_logic_vector(8, 8),
6491 => conv_std_logic_vector(8, 8),
6492 => conv_std_logic_vector(8, 8),
6493 => conv_std_logic_vector(9, 8),
6494 => conv_std_logic_vector(9, 8),
6495 => conv_std_logic_vector(9, 8),
6496 => conv_std_logic_vector(9, 8),
6497 => conv_std_logic_vector(9, 8),
6498 => conv_std_logic_vector(9, 8),
6499 => conv_std_logic_vector(9, 8),
6500 => conv_std_logic_vector(9, 8),
6501 => conv_std_logic_vector(9, 8),
6502 => conv_std_logic_vector(9, 8),
6503 => conv_std_logic_vector(10, 8),
6504 => conv_std_logic_vector(10, 8),
6505 => conv_std_logic_vector(10, 8),
6506 => conv_std_logic_vector(10, 8),
6507 => conv_std_logic_vector(10, 8),
6508 => conv_std_logic_vector(10, 8),
6509 => conv_std_logic_vector(10, 8),
6510 => conv_std_logic_vector(10, 8),
6511 => conv_std_logic_vector(10, 8),
6512 => conv_std_logic_vector(10, 8),
6513 => conv_std_logic_vector(11, 8),
6514 => conv_std_logic_vector(11, 8),
6515 => conv_std_logic_vector(11, 8),
6516 => conv_std_logic_vector(11, 8),
6517 => conv_std_logic_vector(11, 8),
6518 => conv_std_logic_vector(11, 8),
6519 => conv_std_logic_vector(11, 8),
6520 => conv_std_logic_vector(11, 8),
6521 => conv_std_logic_vector(11, 8),
6522 => conv_std_logic_vector(11, 8),
6523 => conv_std_logic_vector(12, 8),
6524 => conv_std_logic_vector(12, 8),
6525 => conv_std_logic_vector(12, 8),
6526 => conv_std_logic_vector(12, 8),
6527 => conv_std_logic_vector(12, 8),
6528 => conv_std_logic_vector(12, 8),
6529 => conv_std_logic_vector(12, 8),
6530 => conv_std_logic_vector(12, 8),
6531 => conv_std_logic_vector(12, 8),
6532 => conv_std_logic_vector(12, 8),
6533 => conv_std_logic_vector(12, 8),
6534 => conv_std_logic_vector(13, 8),
6535 => conv_std_logic_vector(13, 8),
6536 => conv_std_logic_vector(13, 8),
6537 => conv_std_logic_vector(13, 8),
6538 => conv_std_logic_vector(13, 8),
6539 => conv_std_logic_vector(13, 8),
6540 => conv_std_logic_vector(13, 8),
6541 => conv_std_logic_vector(13, 8),
6542 => conv_std_logic_vector(13, 8),
6543 => conv_std_logic_vector(13, 8),
6544 => conv_std_logic_vector(14, 8),
6545 => conv_std_logic_vector(14, 8),
6546 => conv_std_logic_vector(14, 8),
6547 => conv_std_logic_vector(14, 8),
6548 => conv_std_logic_vector(14, 8),
6549 => conv_std_logic_vector(14, 8),
6550 => conv_std_logic_vector(14, 8),
6551 => conv_std_logic_vector(14, 8),
6552 => conv_std_logic_vector(14, 8),
6553 => conv_std_logic_vector(14, 8),
6554 => conv_std_logic_vector(15, 8),
6555 => conv_std_logic_vector(15, 8),
6556 => conv_std_logic_vector(15, 8),
6557 => conv_std_logic_vector(15, 8),
6558 => conv_std_logic_vector(15, 8),
6559 => conv_std_logic_vector(15, 8),
6560 => conv_std_logic_vector(15, 8),
6561 => conv_std_logic_vector(15, 8),
6562 => conv_std_logic_vector(15, 8),
6563 => conv_std_logic_vector(15, 8),
6564 => conv_std_logic_vector(16, 8),
6565 => conv_std_logic_vector(16, 8),
6566 => conv_std_logic_vector(16, 8),
6567 => conv_std_logic_vector(16, 8),
6568 => conv_std_logic_vector(16, 8),
6569 => conv_std_logic_vector(16, 8),
6570 => conv_std_logic_vector(16, 8),
6571 => conv_std_logic_vector(16, 8),
6572 => conv_std_logic_vector(16, 8),
6573 => conv_std_logic_vector(16, 8),
6574 => conv_std_logic_vector(16, 8),
6575 => conv_std_logic_vector(17, 8),
6576 => conv_std_logic_vector(17, 8),
6577 => conv_std_logic_vector(17, 8),
6578 => conv_std_logic_vector(17, 8),
6579 => conv_std_logic_vector(17, 8),
6580 => conv_std_logic_vector(17, 8),
6581 => conv_std_logic_vector(17, 8),
6582 => conv_std_logic_vector(17, 8),
6583 => conv_std_logic_vector(17, 8),
6584 => conv_std_logic_vector(17, 8),
6585 => conv_std_logic_vector(18, 8),
6586 => conv_std_logic_vector(18, 8),
6587 => conv_std_logic_vector(18, 8),
6588 => conv_std_logic_vector(18, 8),
6589 => conv_std_logic_vector(18, 8),
6590 => conv_std_logic_vector(18, 8),
6591 => conv_std_logic_vector(18, 8),
6592 => conv_std_logic_vector(18, 8),
6593 => conv_std_logic_vector(18, 8),
6594 => conv_std_logic_vector(18, 8),
6595 => conv_std_logic_vector(19, 8),
6596 => conv_std_logic_vector(19, 8),
6597 => conv_std_logic_vector(19, 8),
6598 => conv_std_logic_vector(19, 8),
6599 => conv_std_logic_vector(19, 8),
6600 => conv_std_logic_vector(19, 8),
6601 => conv_std_logic_vector(19, 8),
6602 => conv_std_logic_vector(19, 8),
6603 => conv_std_logic_vector(19, 8),
6604 => conv_std_logic_vector(19, 8),
6605 => conv_std_logic_vector(20, 8),
6606 => conv_std_logic_vector(20, 8),
6607 => conv_std_logic_vector(20, 8),
6608 => conv_std_logic_vector(20, 8),
6609 => conv_std_logic_vector(20, 8),
6610 => conv_std_logic_vector(20, 8),
6611 => conv_std_logic_vector(20, 8),
6612 => conv_std_logic_vector(20, 8),
6613 => conv_std_logic_vector(20, 8),
6614 => conv_std_logic_vector(20, 8),
6615 => conv_std_logic_vector(20, 8),
6616 => conv_std_logic_vector(21, 8),
6617 => conv_std_logic_vector(21, 8),
6618 => conv_std_logic_vector(21, 8),
6619 => conv_std_logic_vector(21, 8),
6620 => conv_std_logic_vector(21, 8),
6621 => conv_std_logic_vector(21, 8),
6622 => conv_std_logic_vector(21, 8),
6623 => conv_std_logic_vector(21, 8),
6624 => conv_std_logic_vector(21, 8),
6625 => conv_std_logic_vector(21, 8),
6626 => conv_std_logic_vector(22, 8),
6627 => conv_std_logic_vector(22, 8),
6628 => conv_std_logic_vector(22, 8),
6629 => conv_std_logic_vector(22, 8),
6630 => conv_std_logic_vector(22, 8),
6631 => conv_std_logic_vector(22, 8),
6632 => conv_std_logic_vector(22, 8),
6633 => conv_std_logic_vector(22, 8),
6634 => conv_std_logic_vector(22, 8),
6635 => conv_std_logic_vector(22, 8),
6636 => conv_std_logic_vector(23, 8),
6637 => conv_std_logic_vector(23, 8),
6638 => conv_std_logic_vector(23, 8),
6639 => conv_std_logic_vector(23, 8),
6640 => conv_std_logic_vector(23, 8),
6641 => conv_std_logic_vector(23, 8),
6642 => conv_std_logic_vector(23, 8),
6643 => conv_std_logic_vector(23, 8),
6644 => conv_std_logic_vector(23, 8),
6645 => conv_std_logic_vector(23, 8),
6646 => conv_std_logic_vector(24, 8),
6647 => conv_std_logic_vector(24, 8),
6648 => conv_std_logic_vector(24, 8),
6649 => conv_std_logic_vector(24, 8),
6650 => conv_std_logic_vector(24, 8),
6651 => conv_std_logic_vector(24, 8),
6652 => conv_std_logic_vector(24, 8),
6653 => conv_std_logic_vector(24, 8),
6654 => conv_std_logic_vector(24, 8),
6655 => conv_std_logic_vector(24, 8),
6656 => conv_std_logic_vector(0, 8),
6657 => conv_std_logic_vector(0, 8),
6658 => conv_std_logic_vector(0, 8),
6659 => conv_std_logic_vector(0, 8),
6660 => conv_std_logic_vector(0, 8),
6661 => conv_std_logic_vector(0, 8),
6662 => conv_std_logic_vector(0, 8),
6663 => conv_std_logic_vector(0, 8),
6664 => conv_std_logic_vector(0, 8),
6665 => conv_std_logic_vector(0, 8),
6666 => conv_std_logic_vector(1, 8),
6667 => conv_std_logic_vector(1, 8),
6668 => conv_std_logic_vector(1, 8),
6669 => conv_std_logic_vector(1, 8),
6670 => conv_std_logic_vector(1, 8),
6671 => conv_std_logic_vector(1, 8),
6672 => conv_std_logic_vector(1, 8),
6673 => conv_std_logic_vector(1, 8),
6674 => conv_std_logic_vector(1, 8),
6675 => conv_std_logic_vector(1, 8),
6676 => conv_std_logic_vector(2, 8),
6677 => conv_std_logic_vector(2, 8),
6678 => conv_std_logic_vector(2, 8),
6679 => conv_std_logic_vector(2, 8),
6680 => conv_std_logic_vector(2, 8),
6681 => conv_std_logic_vector(2, 8),
6682 => conv_std_logic_vector(2, 8),
6683 => conv_std_logic_vector(2, 8),
6684 => conv_std_logic_vector(2, 8),
6685 => conv_std_logic_vector(2, 8),
6686 => conv_std_logic_vector(3, 8),
6687 => conv_std_logic_vector(3, 8),
6688 => conv_std_logic_vector(3, 8),
6689 => conv_std_logic_vector(3, 8),
6690 => conv_std_logic_vector(3, 8),
6691 => conv_std_logic_vector(3, 8),
6692 => conv_std_logic_vector(3, 8),
6693 => conv_std_logic_vector(3, 8),
6694 => conv_std_logic_vector(3, 8),
6695 => conv_std_logic_vector(3, 8),
6696 => conv_std_logic_vector(4, 8),
6697 => conv_std_logic_vector(4, 8),
6698 => conv_std_logic_vector(4, 8),
6699 => conv_std_logic_vector(4, 8),
6700 => conv_std_logic_vector(4, 8),
6701 => conv_std_logic_vector(4, 8),
6702 => conv_std_logic_vector(4, 8),
6703 => conv_std_logic_vector(4, 8),
6704 => conv_std_logic_vector(4, 8),
6705 => conv_std_logic_vector(4, 8),
6706 => conv_std_logic_vector(5, 8),
6707 => conv_std_logic_vector(5, 8),
6708 => conv_std_logic_vector(5, 8),
6709 => conv_std_logic_vector(5, 8),
6710 => conv_std_logic_vector(5, 8),
6711 => conv_std_logic_vector(5, 8),
6712 => conv_std_logic_vector(5, 8),
6713 => conv_std_logic_vector(5, 8),
6714 => conv_std_logic_vector(5, 8),
6715 => conv_std_logic_vector(5, 8),
6716 => conv_std_logic_vector(6, 8),
6717 => conv_std_logic_vector(6, 8),
6718 => conv_std_logic_vector(6, 8),
6719 => conv_std_logic_vector(6, 8),
6720 => conv_std_logic_vector(6, 8),
6721 => conv_std_logic_vector(6, 8),
6722 => conv_std_logic_vector(6, 8),
6723 => conv_std_logic_vector(6, 8),
6724 => conv_std_logic_vector(6, 8),
6725 => conv_std_logic_vector(7, 8),
6726 => conv_std_logic_vector(7, 8),
6727 => conv_std_logic_vector(7, 8),
6728 => conv_std_logic_vector(7, 8),
6729 => conv_std_logic_vector(7, 8),
6730 => conv_std_logic_vector(7, 8),
6731 => conv_std_logic_vector(7, 8),
6732 => conv_std_logic_vector(7, 8),
6733 => conv_std_logic_vector(7, 8),
6734 => conv_std_logic_vector(7, 8),
6735 => conv_std_logic_vector(8, 8),
6736 => conv_std_logic_vector(8, 8),
6737 => conv_std_logic_vector(8, 8),
6738 => conv_std_logic_vector(8, 8),
6739 => conv_std_logic_vector(8, 8),
6740 => conv_std_logic_vector(8, 8),
6741 => conv_std_logic_vector(8, 8),
6742 => conv_std_logic_vector(8, 8),
6743 => conv_std_logic_vector(8, 8),
6744 => conv_std_logic_vector(8, 8),
6745 => conv_std_logic_vector(9, 8),
6746 => conv_std_logic_vector(9, 8),
6747 => conv_std_logic_vector(9, 8),
6748 => conv_std_logic_vector(9, 8),
6749 => conv_std_logic_vector(9, 8),
6750 => conv_std_logic_vector(9, 8),
6751 => conv_std_logic_vector(9, 8),
6752 => conv_std_logic_vector(9, 8),
6753 => conv_std_logic_vector(9, 8),
6754 => conv_std_logic_vector(9, 8),
6755 => conv_std_logic_vector(10, 8),
6756 => conv_std_logic_vector(10, 8),
6757 => conv_std_logic_vector(10, 8),
6758 => conv_std_logic_vector(10, 8),
6759 => conv_std_logic_vector(10, 8),
6760 => conv_std_logic_vector(10, 8),
6761 => conv_std_logic_vector(10, 8),
6762 => conv_std_logic_vector(10, 8),
6763 => conv_std_logic_vector(10, 8),
6764 => conv_std_logic_vector(10, 8),
6765 => conv_std_logic_vector(11, 8),
6766 => conv_std_logic_vector(11, 8),
6767 => conv_std_logic_vector(11, 8),
6768 => conv_std_logic_vector(11, 8),
6769 => conv_std_logic_vector(11, 8),
6770 => conv_std_logic_vector(11, 8),
6771 => conv_std_logic_vector(11, 8),
6772 => conv_std_logic_vector(11, 8),
6773 => conv_std_logic_vector(11, 8),
6774 => conv_std_logic_vector(11, 8),
6775 => conv_std_logic_vector(12, 8),
6776 => conv_std_logic_vector(12, 8),
6777 => conv_std_logic_vector(12, 8),
6778 => conv_std_logic_vector(12, 8),
6779 => conv_std_logic_vector(12, 8),
6780 => conv_std_logic_vector(12, 8),
6781 => conv_std_logic_vector(12, 8),
6782 => conv_std_logic_vector(12, 8),
6783 => conv_std_logic_vector(12, 8),
6784 => conv_std_logic_vector(13, 8),
6785 => conv_std_logic_vector(13, 8),
6786 => conv_std_logic_vector(13, 8),
6787 => conv_std_logic_vector(13, 8),
6788 => conv_std_logic_vector(13, 8),
6789 => conv_std_logic_vector(13, 8),
6790 => conv_std_logic_vector(13, 8),
6791 => conv_std_logic_vector(13, 8),
6792 => conv_std_logic_vector(13, 8),
6793 => conv_std_logic_vector(13, 8),
6794 => conv_std_logic_vector(14, 8),
6795 => conv_std_logic_vector(14, 8),
6796 => conv_std_logic_vector(14, 8),
6797 => conv_std_logic_vector(14, 8),
6798 => conv_std_logic_vector(14, 8),
6799 => conv_std_logic_vector(14, 8),
6800 => conv_std_logic_vector(14, 8),
6801 => conv_std_logic_vector(14, 8),
6802 => conv_std_logic_vector(14, 8),
6803 => conv_std_logic_vector(14, 8),
6804 => conv_std_logic_vector(15, 8),
6805 => conv_std_logic_vector(15, 8),
6806 => conv_std_logic_vector(15, 8),
6807 => conv_std_logic_vector(15, 8),
6808 => conv_std_logic_vector(15, 8),
6809 => conv_std_logic_vector(15, 8),
6810 => conv_std_logic_vector(15, 8),
6811 => conv_std_logic_vector(15, 8),
6812 => conv_std_logic_vector(15, 8),
6813 => conv_std_logic_vector(15, 8),
6814 => conv_std_logic_vector(16, 8),
6815 => conv_std_logic_vector(16, 8),
6816 => conv_std_logic_vector(16, 8),
6817 => conv_std_logic_vector(16, 8),
6818 => conv_std_logic_vector(16, 8),
6819 => conv_std_logic_vector(16, 8),
6820 => conv_std_logic_vector(16, 8),
6821 => conv_std_logic_vector(16, 8),
6822 => conv_std_logic_vector(16, 8),
6823 => conv_std_logic_vector(16, 8),
6824 => conv_std_logic_vector(17, 8),
6825 => conv_std_logic_vector(17, 8),
6826 => conv_std_logic_vector(17, 8),
6827 => conv_std_logic_vector(17, 8),
6828 => conv_std_logic_vector(17, 8),
6829 => conv_std_logic_vector(17, 8),
6830 => conv_std_logic_vector(17, 8),
6831 => conv_std_logic_vector(17, 8),
6832 => conv_std_logic_vector(17, 8),
6833 => conv_std_logic_vector(17, 8),
6834 => conv_std_logic_vector(18, 8),
6835 => conv_std_logic_vector(18, 8),
6836 => conv_std_logic_vector(18, 8),
6837 => conv_std_logic_vector(18, 8),
6838 => conv_std_logic_vector(18, 8),
6839 => conv_std_logic_vector(18, 8),
6840 => conv_std_logic_vector(18, 8),
6841 => conv_std_logic_vector(18, 8),
6842 => conv_std_logic_vector(18, 8),
6843 => conv_std_logic_vector(18, 8),
6844 => conv_std_logic_vector(19, 8),
6845 => conv_std_logic_vector(19, 8),
6846 => conv_std_logic_vector(19, 8),
6847 => conv_std_logic_vector(19, 8),
6848 => conv_std_logic_vector(19, 8),
6849 => conv_std_logic_vector(19, 8),
6850 => conv_std_logic_vector(19, 8),
6851 => conv_std_logic_vector(19, 8),
6852 => conv_std_logic_vector(19, 8),
6853 => conv_std_logic_vector(20, 8),
6854 => conv_std_logic_vector(20, 8),
6855 => conv_std_logic_vector(20, 8),
6856 => conv_std_logic_vector(20, 8),
6857 => conv_std_logic_vector(20, 8),
6858 => conv_std_logic_vector(20, 8),
6859 => conv_std_logic_vector(20, 8),
6860 => conv_std_logic_vector(20, 8),
6861 => conv_std_logic_vector(20, 8),
6862 => conv_std_logic_vector(20, 8),
6863 => conv_std_logic_vector(21, 8),
6864 => conv_std_logic_vector(21, 8),
6865 => conv_std_logic_vector(21, 8),
6866 => conv_std_logic_vector(21, 8),
6867 => conv_std_logic_vector(21, 8),
6868 => conv_std_logic_vector(21, 8),
6869 => conv_std_logic_vector(21, 8),
6870 => conv_std_logic_vector(21, 8),
6871 => conv_std_logic_vector(21, 8),
6872 => conv_std_logic_vector(21, 8),
6873 => conv_std_logic_vector(22, 8),
6874 => conv_std_logic_vector(22, 8),
6875 => conv_std_logic_vector(22, 8),
6876 => conv_std_logic_vector(22, 8),
6877 => conv_std_logic_vector(22, 8),
6878 => conv_std_logic_vector(22, 8),
6879 => conv_std_logic_vector(22, 8),
6880 => conv_std_logic_vector(22, 8),
6881 => conv_std_logic_vector(22, 8),
6882 => conv_std_logic_vector(22, 8),
6883 => conv_std_logic_vector(23, 8),
6884 => conv_std_logic_vector(23, 8),
6885 => conv_std_logic_vector(23, 8),
6886 => conv_std_logic_vector(23, 8),
6887 => conv_std_logic_vector(23, 8),
6888 => conv_std_logic_vector(23, 8),
6889 => conv_std_logic_vector(23, 8),
6890 => conv_std_logic_vector(23, 8),
6891 => conv_std_logic_vector(23, 8),
6892 => conv_std_logic_vector(23, 8),
6893 => conv_std_logic_vector(24, 8),
6894 => conv_std_logic_vector(24, 8),
6895 => conv_std_logic_vector(24, 8),
6896 => conv_std_logic_vector(24, 8),
6897 => conv_std_logic_vector(24, 8),
6898 => conv_std_logic_vector(24, 8),
6899 => conv_std_logic_vector(24, 8),
6900 => conv_std_logic_vector(24, 8),
6901 => conv_std_logic_vector(24, 8),
6902 => conv_std_logic_vector(24, 8),
6903 => conv_std_logic_vector(25, 8),
6904 => conv_std_logic_vector(25, 8),
6905 => conv_std_logic_vector(25, 8),
6906 => conv_std_logic_vector(25, 8),
6907 => conv_std_logic_vector(25, 8),
6908 => conv_std_logic_vector(25, 8),
6909 => conv_std_logic_vector(25, 8),
6910 => conv_std_logic_vector(25, 8),
6911 => conv_std_logic_vector(25, 8),
6912 => conv_std_logic_vector(0, 8),
6913 => conv_std_logic_vector(0, 8),
6914 => conv_std_logic_vector(0, 8),
6915 => conv_std_logic_vector(0, 8),
6916 => conv_std_logic_vector(0, 8),
6917 => conv_std_logic_vector(0, 8),
6918 => conv_std_logic_vector(0, 8),
6919 => conv_std_logic_vector(0, 8),
6920 => conv_std_logic_vector(0, 8),
6921 => conv_std_logic_vector(0, 8),
6922 => conv_std_logic_vector(1, 8),
6923 => conv_std_logic_vector(1, 8),
6924 => conv_std_logic_vector(1, 8),
6925 => conv_std_logic_vector(1, 8),
6926 => conv_std_logic_vector(1, 8),
6927 => conv_std_logic_vector(1, 8),
6928 => conv_std_logic_vector(1, 8),
6929 => conv_std_logic_vector(1, 8),
6930 => conv_std_logic_vector(1, 8),
6931 => conv_std_logic_vector(2, 8),
6932 => conv_std_logic_vector(2, 8),
6933 => conv_std_logic_vector(2, 8),
6934 => conv_std_logic_vector(2, 8),
6935 => conv_std_logic_vector(2, 8),
6936 => conv_std_logic_vector(2, 8),
6937 => conv_std_logic_vector(2, 8),
6938 => conv_std_logic_vector(2, 8),
6939 => conv_std_logic_vector(2, 8),
6940 => conv_std_logic_vector(2, 8),
6941 => conv_std_logic_vector(3, 8),
6942 => conv_std_logic_vector(3, 8),
6943 => conv_std_logic_vector(3, 8),
6944 => conv_std_logic_vector(3, 8),
6945 => conv_std_logic_vector(3, 8),
6946 => conv_std_logic_vector(3, 8),
6947 => conv_std_logic_vector(3, 8),
6948 => conv_std_logic_vector(3, 8),
6949 => conv_std_logic_vector(3, 8),
6950 => conv_std_logic_vector(4, 8),
6951 => conv_std_logic_vector(4, 8),
6952 => conv_std_logic_vector(4, 8),
6953 => conv_std_logic_vector(4, 8),
6954 => conv_std_logic_vector(4, 8),
6955 => conv_std_logic_vector(4, 8),
6956 => conv_std_logic_vector(4, 8),
6957 => conv_std_logic_vector(4, 8),
6958 => conv_std_logic_vector(4, 8),
6959 => conv_std_logic_vector(4, 8),
6960 => conv_std_logic_vector(5, 8),
6961 => conv_std_logic_vector(5, 8),
6962 => conv_std_logic_vector(5, 8),
6963 => conv_std_logic_vector(5, 8),
6964 => conv_std_logic_vector(5, 8),
6965 => conv_std_logic_vector(5, 8),
6966 => conv_std_logic_vector(5, 8),
6967 => conv_std_logic_vector(5, 8),
6968 => conv_std_logic_vector(5, 8),
6969 => conv_std_logic_vector(6, 8),
6970 => conv_std_logic_vector(6, 8),
6971 => conv_std_logic_vector(6, 8),
6972 => conv_std_logic_vector(6, 8),
6973 => conv_std_logic_vector(6, 8),
6974 => conv_std_logic_vector(6, 8),
6975 => conv_std_logic_vector(6, 8),
6976 => conv_std_logic_vector(6, 8),
6977 => conv_std_logic_vector(6, 8),
6978 => conv_std_logic_vector(6, 8),
6979 => conv_std_logic_vector(7, 8),
6980 => conv_std_logic_vector(7, 8),
6981 => conv_std_logic_vector(7, 8),
6982 => conv_std_logic_vector(7, 8),
6983 => conv_std_logic_vector(7, 8),
6984 => conv_std_logic_vector(7, 8),
6985 => conv_std_logic_vector(7, 8),
6986 => conv_std_logic_vector(7, 8),
6987 => conv_std_logic_vector(7, 8),
6988 => conv_std_logic_vector(8, 8),
6989 => conv_std_logic_vector(8, 8),
6990 => conv_std_logic_vector(8, 8),
6991 => conv_std_logic_vector(8, 8),
6992 => conv_std_logic_vector(8, 8),
6993 => conv_std_logic_vector(8, 8),
6994 => conv_std_logic_vector(8, 8),
6995 => conv_std_logic_vector(8, 8),
6996 => conv_std_logic_vector(8, 8),
6997 => conv_std_logic_vector(8, 8),
6998 => conv_std_logic_vector(9, 8),
6999 => conv_std_logic_vector(9, 8),
7000 => conv_std_logic_vector(9, 8),
7001 => conv_std_logic_vector(9, 8),
7002 => conv_std_logic_vector(9, 8),
7003 => conv_std_logic_vector(9, 8),
7004 => conv_std_logic_vector(9, 8),
7005 => conv_std_logic_vector(9, 8),
7006 => conv_std_logic_vector(9, 8),
7007 => conv_std_logic_vector(10, 8),
7008 => conv_std_logic_vector(10, 8),
7009 => conv_std_logic_vector(10, 8),
7010 => conv_std_logic_vector(10, 8),
7011 => conv_std_logic_vector(10, 8),
7012 => conv_std_logic_vector(10, 8),
7013 => conv_std_logic_vector(10, 8),
7014 => conv_std_logic_vector(10, 8),
7015 => conv_std_logic_vector(10, 8),
7016 => conv_std_logic_vector(10, 8),
7017 => conv_std_logic_vector(11, 8),
7018 => conv_std_logic_vector(11, 8),
7019 => conv_std_logic_vector(11, 8),
7020 => conv_std_logic_vector(11, 8),
7021 => conv_std_logic_vector(11, 8),
7022 => conv_std_logic_vector(11, 8),
7023 => conv_std_logic_vector(11, 8),
7024 => conv_std_logic_vector(11, 8),
7025 => conv_std_logic_vector(11, 8),
7026 => conv_std_logic_vector(12, 8),
7027 => conv_std_logic_vector(12, 8),
7028 => conv_std_logic_vector(12, 8),
7029 => conv_std_logic_vector(12, 8),
7030 => conv_std_logic_vector(12, 8),
7031 => conv_std_logic_vector(12, 8),
7032 => conv_std_logic_vector(12, 8),
7033 => conv_std_logic_vector(12, 8),
7034 => conv_std_logic_vector(12, 8),
7035 => conv_std_logic_vector(12, 8),
7036 => conv_std_logic_vector(13, 8),
7037 => conv_std_logic_vector(13, 8),
7038 => conv_std_logic_vector(13, 8),
7039 => conv_std_logic_vector(13, 8),
7040 => conv_std_logic_vector(13, 8),
7041 => conv_std_logic_vector(13, 8),
7042 => conv_std_logic_vector(13, 8),
7043 => conv_std_logic_vector(13, 8),
7044 => conv_std_logic_vector(13, 8),
7045 => conv_std_logic_vector(14, 8),
7046 => conv_std_logic_vector(14, 8),
7047 => conv_std_logic_vector(14, 8),
7048 => conv_std_logic_vector(14, 8),
7049 => conv_std_logic_vector(14, 8),
7050 => conv_std_logic_vector(14, 8),
7051 => conv_std_logic_vector(14, 8),
7052 => conv_std_logic_vector(14, 8),
7053 => conv_std_logic_vector(14, 8),
7054 => conv_std_logic_vector(14, 8),
7055 => conv_std_logic_vector(15, 8),
7056 => conv_std_logic_vector(15, 8),
7057 => conv_std_logic_vector(15, 8),
7058 => conv_std_logic_vector(15, 8),
7059 => conv_std_logic_vector(15, 8),
7060 => conv_std_logic_vector(15, 8),
7061 => conv_std_logic_vector(15, 8),
7062 => conv_std_logic_vector(15, 8),
7063 => conv_std_logic_vector(15, 8),
7064 => conv_std_logic_vector(16, 8),
7065 => conv_std_logic_vector(16, 8),
7066 => conv_std_logic_vector(16, 8),
7067 => conv_std_logic_vector(16, 8),
7068 => conv_std_logic_vector(16, 8),
7069 => conv_std_logic_vector(16, 8),
7070 => conv_std_logic_vector(16, 8),
7071 => conv_std_logic_vector(16, 8),
7072 => conv_std_logic_vector(16, 8),
7073 => conv_std_logic_vector(16, 8),
7074 => conv_std_logic_vector(17, 8),
7075 => conv_std_logic_vector(17, 8),
7076 => conv_std_logic_vector(17, 8),
7077 => conv_std_logic_vector(17, 8),
7078 => conv_std_logic_vector(17, 8),
7079 => conv_std_logic_vector(17, 8),
7080 => conv_std_logic_vector(17, 8),
7081 => conv_std_logic_vector(17, 8),
7082 => conv_std_logic_vector(17, 8),
7083 => conv_std_logic_vector(18, 8),
7084 => conv_std_logic_vector(18, 8),
7085 => conv_std_logic_vector(18, 8),
7086 => conv_std_logic_vector(18, 8),
7087 => conv_std_logic_vector(18, 8),
7088 => conv_std_logic_vector(18, 8),
7089 => conv_std_logic_vector(18, 8),
7090 => conv_std_logic_vector(18, 8),
7091 => conv_std_logic_vector(18, 8),
7092 => conv_std_logic_vector(18, 8),
7093 => conv_std_logic_vector(19, 8),
7094 => conv_std_logic_vector(19, 8),
7095 => conv_std_logic_vector(19, 8),
7096 => conv_std_logic_vector(19, 8),
7097 => conv_std_logic_vector(19, 8),
7098 => conv_std_logic_vector(19, 8),
7099 => conv_std_logic_vector(19, 8),
7100 => conv_std_logic_vector(19, 8),
7101 => conv_std_logic_vector(19, 8),
7102 => conv_std_logic_vector(20, 8),
7103 => conv_std_logic_vector(20, 8),
7104 => conv_std_logic_vector(20, 8),
7105 => conv_std_logic_vector(20, 8),
7106 => conv_std_logic_vector(20, 8),
7107 => conv_std_logic_vector(20, 8),
7108 => conv_std_logic_vector(20, 8),
7109 => conv_std_logic_vector(20, 8),
7110 => conv_std_logic_vector(20, 8),
7111 => conv_std_logic_vector(20, 8),
7112 => conv_std_logic_vector(21, 8),
7113 => conv_std_logic_vector(21, 8),
7114 => conv_std_logic_vector(21, 8),
7115 => conv_std_logic_vector(21, 8),
7116 => conv_std_logic_vector(21, 8),
7117 => conv_std_logic_vector(21, 8),
7118 => conv_std_logic_vector(21, 8),
7119 => conv_std_logic_vector(21, 8),
7120 => conv_std_logic_vector(21, 8),
7121 => conv_std_logic_vector(22, 8),
7122 => conv_std_logic_vector(22, 8),
7123 => conv_std_logic_vector(22, 8),
7124 => conv_std_logic_vector(22, 8),
7125 => conv_std_logic_vector(22, 8),
7126 => conv_std_logic_vector(22, 8),
7127 => conv_std_logic_vector(22, 8),
7128 => conv_std_logic_vector(22, 8),
7129 => conv_std_logic_vector(22, 8),
7130 => conv_std_logic_vector(22, 8),
7131 => conv_std_logic_vector(23, 8),
7132 => conv_std_logic_vector(23, 8),
7133 => conv_std_logic_vector(23, 8),
7134 => conv_std_logic_vector(23, 8),
7135 => conv_std_logic_vector(23, 8),
7136 => conv_std_logic_vector(23, 8),
7137 => conv_std_logic_vector(23, 8),
7138 => conv_std_logic_vector(23, 8),
7139 => conv_std_logic_vector(23, 8),
7140 => conv_std_logic_vector(24, 8),
7141 => conv_std_logic_vector(24, 8),
7142 => conv_std_logic_vector(24, 8),
7143 => conv_std_logic_vector(24, 8),
7144 => conv_std_logic_vector(24, 8),
7145 => conv_std_logic_vector(24, 8),
7146 => conv_std_logic_vector(24, 8),
7147 => conv_std_logic_vector(24, 8),
7148 => conv_std_logic_vector(24, 8),
7149 => conv_std_logic_vector(24, 8),
7150 => conv_std_logic_vector(25, 8),
7151 => conv_std_logic_vector(25, 8),
7152 => conv_std_logic_vector(25, 8),
7153 => conv_std_logic_vector(25, 8),
7154 => conv_std_logic_vector(25, 8),
7155 => conv_std_logic_vector(25, 8),
7156 => conv_std_logic_vector(25, 8),
7157 => conv_std_logic_vector(25, 8),
7158 => conv_std_logic_vector(25, 8),
7159 => conv_std_logic_vector(26, 8),
7160 => conv_std_logic_vector(26, 8),
7161 => conv_std_logic_vector(26, 8),
7162 => conv_std_logic_vector(26, 8),
7163 => conv_std_logic_vector(26, 8),
7164 => conv_std_logic_vector(26, 8),
7165 => conv_std_logic_vector(26, 8),
7166 => conv_std_logic_vector(26, 8),
7167 => conv_std_logic_vector(26, 8),
7168 => conv_std_logic_vector(0, 8),
7169 => conv_std_logic_vector(0, 8),
7170 => conv_std_logic_vector(0, 8),
7171 => conv_std_logic_vector(0, 8),
7172 => conv_std_logic_vector(0, 8),
7173 => conv_std_logic_vector(0, 8),
7174 => conv_std_logic_vector(0, 8),
7175 => conv_std_logic_vector(0, 8),
7176 => conv_std_logic_vector(0, 8),
7177 => conv_std_logic_vector(0, 8),
7178 => conv_std_logic_vector(1, 8),
7179 => conv_std_logic_vector(1, 8),
7180 => conv_std_logic_vector(1, 8),
7181 => conv_std_logic_vector(1, 8),
7182 => conv_std_logic_vector(1, 8),
7183 => conv_std_logic_vector(1, 8),
7184 => conv_std_logic_vector(1, 8),
7185 => conv_std_logic_vector(1, 8),
7186 => conv_std_logic_vector(1, 8),
7187 => conv_std_logic_vector(2, 8),
7188 => conv_std_logic_vector(2, 8),
7189 => conv_std_logic_vector(2, 8),
7190 => conv_std_logic_vector(2, 8),
7191 => conv_std_logic_vector(2, 8),
7192 => conv_std_logic_vector(2, 8),
7193 => conv_std_logic_vector(2, 8),
7194 => conv_std_logic_vector(2, 8),
7195 => conv_std_logic_vector(2, 8),
7196 => conv_std_logic_vector(3, 8),
7197 => conv_std_logic_vector(3, 8),
7198 => conv_std_logic_vector(3, 8),
7199 => conv_std_logic_vector(3, 8),
7200 => conv_std_logic_vector(3, 8),
7201 => conv_std_logic_vector(3, 8),
7202 => conv_std_logic_vector(3, 8),
7203 => conv_std_logic_vector(3, 8),
7204 => conv_std_logic_vector(3, 8),
7205 => conv_std_logic_vector(4, 8),
7206 => conv_std_logic_vector(4, 8),
7207 => conv_std_logic_vector(4, 8),
7208 => conv_std_logic_vector(4, 8),
7209 => conv_std_logic_vector(4, 8),
7210 => conv_std_logic_vector(4, 8),
7211 => conv_std_logic_vector(4, 8),
7212 => conv_std_logic_vector(4, 8),
7213 => conv_std_logic_vector(4, 8),
7214 => conv_std_logic_vector(5, 8),
7215 => conv_std_logic_vector(5, 8),
7216 => conv_std_logic_vector(5, 8),
7217 => conv_std_logic_vector(5, 8),
7218 => conv_std_logic_vector(5, 8),
7219 => conv_std_logic_vector(5, 8),
7220 => conv_std_logic_vector(5, 8),
7221 => conv_std_logic_vector(5, 8),
7222 => conv_std_logic_vector(5, 8),
7223 => conv_std_logic_vector(6, 8),
7224 => conv_std_logic_vector(6, 8),
7225 => conv_std_logic_vector(6, 8),
7226 => conv_std_logic_vector(6, 8),
7227 => conv_std_logic_vector(6, 8),
7228 => conv_std_logic_vector(6, 8),
7229 => conv_std_logic_vector(6, 8),
7230 => conv_std_logic_vector(6, 8),
7231 => conv_std_logic_vector(6, 8),
7232 => conv_std_logic_vector(7, 8),
7233 => conv_std_logic_vector(7, 8),
7234 => conv_std_logic_vector(7, 8),
7235 => conv_std_logic_vector(7, 8),
7236 => conv_std_logic_vector(7, 8),
7237 => conv_std_logic_vector(7, 8),
7238 => conv_std_logic_vector(7, 8),
7239 => conv_std_logic_vector(7, 8),
7240 => conv_std_logic_vector(7, 8),
7241 => conv_std_logic_vector(7, 8),
7242 => conv_std_logic_vector(8, 8),
7243 => conv_std_logic_vector(8, 8),
7244 => conv_std_logic_vector(8, 8),
7245 => conv_std_logic_vector(8, 8),
7246 => conv_std_logic_vector(8, 8),
7247 => conv_std_logic_vector(8, 8),
7248 => conv_std_logic_vector(8, 8),
7249 => conv_std_logic_vector(8, 8),
7250 => conv_std_logic_vector(8, 8),
7251 => conv_std_logic_vector(9, 8),
7252 => conv_std_logic_vector(9, 8),
7253 => conv_std_logic_vector(9, 8),
7254 => conv_std_logic_vector(9, 8),
7255 => conv_std_logic_vector(9, 8),
7256 => conv_std_logic_vector(9, 8),
7257 => conv_std_logic_vector(9, 8),
7258 => conv_std_logic_vector(9, 8),
7259 => conv_std_logic_vector(9, 8),
7260 => conv_std_logic_vector(10, 8),
7261 => conv_std_logic_vector(10, 8),
7262 => conv_std_logic_vector(10, 8),
7263 => conv_std_logic_vector(10, 8),
7264 => conv_std_logic_vector(10, 8),
7265 => conv_std_logic_vector(10, 8),
7266 => conv_std_logic_vector(10, 8),
7267 => conv_std_logic_vector(10, 8),
7268 => conv_std_logic_vector(10, 8),
7269 => conv_std_logic_vector(11, 8),
7270 => conv_std_logic_vector(11, 8),
7271 => conv_std_logic_vector(11, 8),
7272 => conv_std_logic_vector(11, 8),
7273 => conv_std_logic_vector(11, 8),
7274 => conv_std_logic_vector(11, 8),
7275 => conv_std_logic_vector(11, 8),
7276 => conv_std_logic_vector(11, 8),
7277 => conv_std_logic_vector(11, 8),
7278 => conv_std_logic_vector(12, 8),
7279 => conv_std_logic_vector(12, 8),
7280 => conv_std_logic_vector(12, 8),
7281 => conv_std_logic_vector(12, 8),
7282 => conv_std_logic_vector(12, 8),
7283 => conv_std_logic_vector(12, 8),
7284 => conv_std_logic_vector(12, 8),
7285 => conv_std_logic_vector(12, 8),
7286 => conv_std_logic_vector(12, 8),
7287 => conv_std_logic_vector(13, 8),
7288 => conv_std_logic_vector(13, 8),
7289 => conv_std_logic_vector(13, 8),
7290 => conv_std_logic_vector(13, 8),
7291 => conv_std_logic_vector(13, 8),
7292 => conv_std_logic_vector(13, 8),
7293 => conv_std_logic_vector(13, 8),
7294 => conv_std_logic_vector(13, 8),
7295 => conv_std_logic_vector(13, 8),
7296 => conv_std_logic_vector(14, 8),
7297 => conv_std_logic_vector(14, 8),
7298 => conv_std_logic_vector(14, 8),
7299 => conv_std_logic_vector(14, 8),
7300 => conv_std_logic_vector(14, 8),
7301 => conv_std_logic_vector(14, 8),
7302 => conv_std_logic_vector(14, 8),
7303 => conv_std_logic_vector(14, 8),
7304 => conv_std_logic_vector(14, 8),
7305 => conv_std_logic_vector(14, 8),
7306 => conv_std_logic_vector(15, 8),
7307 => conv_std_logic_vector(15, 8),
7308 => conv_std_logic_vector(15, 8),
7309 => conv_std_logic_vector(15, 8),
7310 => conv_std_logic_vector(15, 8),
7311 => conv_std_logic_vector(15, 8),
7312 => conv_std_logic_vector(15, 8),
7313 => conv_std_logic_vector(15, 8),
7314 => conv_std_logic_vector(15, 8),
7315 => conv_std_logic_vector(16, 8),
7316 => conv_std_logic_vector(16, 8),
7317 => conv_std_logic_vector(16, 8),
7318 => conv_std_logic_vector(16, 8),
7319 => conv_std_logic_vector(16, 8),
7320 => conv_std_logic_vector(16, 8),
7321 => conv_std_logic_vector(16, 8),
7322 => conv_std_logic_vector(16, 8),
7323 => conv_std_logic_vector(16, 8),
7324 => conv_std_logic_vector(17, 8),
7325 => conv_std_logic_vector(17, 8),
7326 => conv_std_logic_vector(17, 8),
7327 => conv_std_logic_vector(17, 8),
7328 => conv_std_logic_vector(17, 8),
7329 => conv_std_logic_vector(17, 8),
7330 => conv_std_logic_vector(17, 8),
7331 => conv_std_logic_vector(17, 8),
7332 => conv_std_logic_vector(17, 8),
7333 => conv_std_logic_vector(18, 8),
7334 => conv_std_logic_vector(18, 8),
7335 => conv_std_logic_vector(18, 8),
7336 => conv_std_logic_vector(18, 8),
7337 => conv_std_logic_vector(18, 8),
7338 => conv_std_logic_vector(18, 8),
7339 => conv_std_logic_vector(18, 8),
7340 => conv_std_logic_vector(18, 8),
7341 => conv_std_logic_vector(18, 8),
7342 => conv_std_logic_vector(19, 8),
7343 => conv_std_logic_vector(19, 8),
7344 => conv_std_logic_vector(19, 8),
7345 => conv_std_logic_vector(19, 8),
7346 => conv_std_logic_vector(19, 8),
7347 => conv_std_logic_vector(19, 8),
7348 => conv_std_logic_vector(19, 8),
7349 => conv_std_logic_vector(19, 8),
7350 => conv_std_logic_vector(19, 8),
7351 => conv_std_logic_vector(20, 8),
7352 => conv_std_logic_vector(20, 8),
7353 => conv_std_logic_vector(20, 8),
7354 => conv_std_logic_vector(20, 8),
7355 => conv_std_logic_vector(20, 8),
7356 => conv_std_logic_vector(20, 8),
7357 => conv_std_logic_vector(20, 8),
7358 => conv_std_logic_vector(20, 8),
7359 => conv_std_logic_vector(20, 8),
7360 => conv_std_logic_vector(21, 8),
7361 => conv_std_logic_vector(21, 8),
7362 => conv_std_logic_vector(21, 8),
7363 => conv_std_logic_vector(21, 8),
7364 => conv_std_logic_vector(21, 8),
7365 => conv_std_logic_vector(21, 8),
7366 => conv_std_logic_vector(21, 8),
7367 => conv_std_logic_vector(21, 8),
7368 => conv_std_logic_vector(21, 8),
7369 => conv_std_logic_vector(21, 8),
7370 => conv_std_logic_vector(22, 8),
7371 => conv_std_logic_vector(22, 8),
7372 => conv_std_logic_vector(22, 8),
7373 => conv_std_logic_vector(22, 8),
7374 => conv_std_logic_vector(22, 8),
7375 => conv_std_logic_vector(22, 8),
7376 => conv_std_logic_vector(22, 8),
7377 => conv_std_logic_vector(22, 8),
7378 => conv_std_logic_vector(22, 8),
7379 => conv_std_logic_vector(23, 8),
7380 => conv_std_logic_vector(23, 8),
7381 => conv_std_logic_vector(23, 8),
7382 => conv_std_logic_vector(23, 8),
7383 => conv_std_logic_vector(23, 8),
7384 => conv_std_logic_vector(23, 8),
7385 => conv_std_logic_vector(23, 8),
7386 => conv_std_logic_vector(23, 8),
7387 => conv_std_logic_vector(23, 8),
7388 => conv_std_logic_vector(24, 8),
7389 => conv_std_logic_vector(24, 8),
7390 => conv_std_logic_vector(24, 8),
7391 => conv_std_logic_vector(24, 8),
7392 => conv_std_logic_vector(24, 8),
7393 => conv_std_logic_vector(24, 8),
7394 => conv_std_logic_vector(24, 8),
7395 => conv_std_logic_vector(24, 8),
7396 => conv_std_logic_vector(24, 8),
7397 => conv_std_logic_vector(25, 8),
7398 => conv_std_logic_vector(25, 8),
7399 => conv_std_logic_vector(25, 8),
7400 => conv_std_logic_vector(25, 8),
7401 => conv_std_logic_vector(25, 8),
7402 => conv_std_logic_vector(25, 8),
7403 => conv_std_logic_vector(25, 8),
7404 => conv_std_logic_vector(25, 8),
7405 => conv_std_logic_vector(25, 8),
7406 => conv_std_logic_vector(26, 8),
7407 => conv_std_logic_vector(26, 8),
7408 => conv_std_logic_vector(26, 8),
7409 => conv_std_logic_vector(26, 8),
7410 => conv_std_logic_vector(26, 8),
7411 => conv_std_logic_vector(26, 8),
7412 => conv_std_logic_vector(26, 8),
7413 => conv_std_logic_vector(26, 8),
7414 => conv_std_logic_vector(26, 8),
7415 => conv_std_logic_vector(27, 8),
7416 => conv_std_logic_vector(27, 8),
7417 => conv_std_logic_vector(27, 8),
7418 => conv_std_logic_vector(27, 8),
7419 => conv_std_logic_vector(27, 8),
7420 => conv_std_logic_vector(27, 8),
7421 => conv_std_logic_vector(27, 8),
7422 => conv_std_logic_vector(27, 8),
7423 => conv_std_logic_vector(27, 8),
7424 => conv_std_logic_vector(0, 8),
7425 => conv_std_logic_vector(0, 8),
7426 => conv_std_logic_vector(0, 8),
7427 => conv_std_logic_vector(0, 8),
7428 => conv_std_logic_vector(0, 8),
7429 => conv_std_logic_vector(0, 8),
7430 => conv_std_logic_vector(0, 8),
7431 => conv_std_logic_vector(0, 8),
7432 => conv_std_logic_vector(0, 8),
7433 => conv_std_logic_vector(1, 8),
7434 => conv_std_logic_vector(1, 8),
7435 => conv_std_logic_vector(1, 8),
7436 => conv_std_logic_vector(1, 8),
7437 => conv_std_logic_vector(1, 8),
7438 => conv_std_logic_vector(1, 8),
7439 => conv_std_logic_vector(1, 8),
7440 => conv_std_logic_vector(1, 8),
7441 => conv_std_logic_vector(1, 8),
7442 => conv_std_logic_vector(2, 8),
7443 => conv_std_logic_vector(2, 8),
7444 => conv_std_logic_vector(2, 8),
7445 => conv_std_logic_vector(2, 8),
7446 => conv_std_logic_vector(2, 8),
7447 => conv_std_logic_vector(2, 8),
7448 => conv_std_logic_vector(2, 8),
7449 => conv_std_logic_vector(2, 8),
7450 => conv_std_logic_vector(2, 8),
7451 => conv_std_logic_vector(3, 8),
7452 => conv_std_logic_vector(3, 8),
7453 => conv_std_logic_vector(3, 8),
7454 => conv_std_logic_vector(3, 8),
7455 => conv_std_logic_vector(3, 8),
7456 => conv_std_logic_vector(3, 8),
7457 => conv_std_logic_vector(3, 8),
7458 => conv_std_logic_vector(3, 8),
7459 => conv_std_logic_vector(3, 8),
7460 => conv_std_logic_vector(4, 8),
7461 => conv_std_logic_vector(4, 8),
7462 => conv_std_logic_vector(4, 8),
7463 => conv_std_logic_vector(4, 8),
7464 => conv_std_logic_vector(4, 8),
7465 => conv_std_logic_vector(4, 8),
7466 => conv_std_logic_vector(4, 8),
7467 => conv_std_logic_vector(4, 8),
7468 => conv_std_logic_vector(4, 8),
7469 => conv_std_logic_vector(5, 8),
7470 => conv_std_logic_vector(5, 8),
7471 => conv_std_logic_vector(5, 8),
7472 => conv_std_logic_vector(5, 8),
7473 => conv_std_logic_vector(5, 8),
7474 => conv_std_logic_vector(5, 8),
7475 => conv_std_logic_vector(5, 8),
7476 => conv_std_logic_vector(5, 8),
7477 => conv_std_logic_vector(6, 8),
7478 => conv_std_logic_vector(6, 8),
7479 => conv_std_logic_vector(6, 8),
7480 => conv_std_logic_vector(6, 8),
7481 => conv_std_logic_vector(6, 8),
7482 => conv_std_logic_vector(6, 8),
7483 => conv_std_logic_vector(6, 8),
7484 => conv_std_logic_vector(6, 8),
7485 => conv_std_logic_vector(6, 8),
7486 => conv_std_logic_vector(7, 8),
7487 => conv_std_logic_vector(7, 8),
7488 => conv_std_logic_vector(7, 8),
7489 => conv_std_logic_vector(7, 8),
7490 => conv_std_logic_vector(7, 8),
7491 => conv_std_logic_vector(7, 8),
7492 => conv_std_logic_vector(7, 8),
7493 => conv_std_logic_vector(7, 8),
7494 => conv_std_logic_vector(7, 8),
7495 => conv_std_logic_vector(8, 8),
7496 => conv_std_logic_vector(8, 8),
7497 => conv_std_logic_vector(8, 8),
7498 => conv_std_logic_vector(8, 8),
7499 => conv_std_logic_vector(8, 8),
7500 => conv_std_logic_vector(8, 8),
7501 => conv_std_logic_vector(8, 8),
7502 => conv_std_logic_vector(8, 8),
7503 => conv_std_logic_vector(8, 8),
7504 => conv_std_logic_vector(9, 8),
7505 => conv_std_logic_vector(9, 8),
7506 => conv_std_logic_vector(9, 8),
7507 => conv_std_logic_vector(9, 8),
7508 => conv_std_logic_vector(9, 8),
7509 => conv_std_logic_vector(9, 8),
7510 => conv_std_logic_vector(9, 8),
7511 => conv_std_logic_vector(9, 8),
7512 => conv_std_logic_vector(9, 8),
7513 => conv_std_logic_vector(10, 8),
7514 => conv_std_logic_vector(10, 8),
7515 => conv_std_logic_vector(10, 8),
7516 => conv_std_logic_vector(10, 8),
7517 => conv_std_logic_vector(10, 8),
7518 => conv_std_logic_vector(10, 8),
7519 => conv_std_logic_vector(10, 8),
7520 => conv_std_logic_vector(10, 8),
7521 => conv_std_logic_vector(10, 8),
7522 => conv_std_logic_vector(11, 8),
7523 => conv_std_logic_vector(11, 8),
7524 => conv_std_logic_vector(11, 8),
7525 => conv_std_logic_vector(11, 8),
7526 => conv_std_logic_vector(11, 8),
7527 => conv_std_logic_vector(11, 8),
7528 => conv_std_logic_vector(11, 8),
7529 => conv_std_logic_vector(11, 8),
7530 => conv_std_logic_vector(12, 8),
7531 => conv_std_logic_vector(12, 8),
7532 => conv_std_logic_vector(12, 8),
7533 => conv_std_logic_vector(12, 8),
7534 => conv_std_logic_vector(12, 8),
7535 => conv_std_logic_vector(12, 8),
7536 => conv_std_logic_vector(12, 8),
7537 => conv_std_logic_vector(12, 8),
7538 => conv_std_logic_vector(12, 8),
7539 => conv_std_logic_vector(13, 8),
7540 => conv_std_logic_vector(13, 8),
7541 => conv_std_logic_vector(13, 8),
7542 => conv_std_logic_vector(13, 8),
7543 => conv_std_logic_vector(13, 8),
7544 => conv_std_logic_vector(13, 8),
7545 => conv_std_logic_vector(13, 8),
7546 => conv_std_logic_vector(13, 8),
7547 => conv_std_logic_vector(13, 8),
7548 => conv_std_logic_vector(14, 8),
7549 => conv_std_logic_vector(14, 8),
7550 => conv_std_logic_vector(14, 8),
7551 => conv_std_logic_vector(14, 8),
7552 => conv_std_logic_vector(14, 8),
7553 => conv_std_logic_vector(14, 8),
7554 => conv_std_logic_vector(14, 8),
7555 => conv_std_logic_vector(14, 8),
7556 => conv_std_logic_vector(14, 8),
7557 => conv_std_logic_vector(15, 8),
7558 => conv_std_logic_vector(15, 8),
7559 => conv_std_logic_vector(15, 8),
7560 => conv_std_logic_vector(15, 8),
7561 => conv_std_logic_vector(15, 8),
7562 => conv_std_logic_vector(15, 8),
7563 => conv_std_logic_vector(15, 8),
7564 => conv_std_logic_vector(15, 8),
7565 => conv_std_logic_vector(15, 8),
7566 => conv_std_logic_vector(16, 8),
7567 => conv_std_logic_vector(16, 8),
7568 => conv_std_logic_vector(16, 8),
7569 => conv_std_logic_vector(16, 8),
7570 => conv_std_logic_vector(16, 8),
7571 => conv_std_logic_vector(16, 8),
7572 => conv_std_logic_vector(16, 8),
7573 => conv_std_logic_vector(16, 8),
7574 => conv_std_logic_vector(16, 8),
7575 => conv_std_logic_vector(17, 8),
7576 => conv_std_logic_vector(17, 8),
7577 => conv_std_logic_vector(17, 8),
7578 => conv_std_logic_vector(17, 8),
7579 => conv_std_logic_vector(17, 8),
7580 => conv_std_logic_vector(17, 8),
7581 => conv_std_logic_vector(17, 8),
7582 => conv_std_logic_vector(17, 8),
7583 => conv_std_logic_vector(18, 8),
7584 => conv_std_logic_vector(18, 8),
7585 => conv_std_logic_vector(18, 8),
7586 => conv_std_logic_vector(18, 8),
7587 => conv_std_logic_vector(18, 8),
7588 => conv_std_logic_vector(18, 8),
7589 => conv_std_logic_vector(18, 8),
7590 => conv_std_logic_vector(18, 8),
7591 => conv_std_logic_vector(18, 8),
7592 => conv_std_logic_vector(19, 8),
7593 => conv_std_logic_vector(19, 8),
7594 => conv_std_logic_vector(19, 8),
7595 => conv_std_logic_vector(19, 8),
7596 => conv_std_logic_vector(19, 8),
7597 => conv_std_logic_vector(19, 8),
7598 => conv_std_logic_vector(19, 8),
7599 => conv_std_logic_vector(19, 8),
7600 => conv_std_logic_vector(19, 8),
7601 => conv_std_logic_vector(20, 8),
7602 => conv_std_logic_vector(20, 8),
7603 => conv_std_logic_vector(20, 8),
7604 => conv_std_logic_vector(20, 8),
7605 => conv_std_logic_vector(20, 8),
7606 => conv_std_logic_vector(20, 8),
7607 => conv_std_logic_vector(20, 8),
7608 => conv_std_logic_vector(20, 8),
7609 => conv_std_logic_vector(20, 8),
7610 => conv_std_logic_vector(21, 8),
7611 => conv_std_logic_vector(21, 8),
7612 => conv_std_logic_vector(21, 8),
7613 => conv_std_logic_vector(21, 8),
7614 => conv_std_logic_vector(21, 8),
7615 => conv_std_logic_vector(21, 8),
7616 => conv_std_logic_vector(21, 8),
7617 => conv_std_logic_vector(21, 8),
7618 => conv_std_logic_vector(21, 8),
7619 => conv_std_logic_vector(22, 8),
7620 => conv_std_logic_vector(22, 8),
7621 => conv_std_logic_vector(22, 8),
7622 => conv_std_logic_vector(22, 8),
7623 => conv_std_logic_vector(22, 8),
7624 => conv_std_logic_vector(22, 8),
7625 => conv_std_logic_vector(22, 8),
7626 => conv_std_logic_vector(22, 8),
7627 => conv_std_logic_vector(22, 8),
7628 => conv_std_logic_vector(23, 8),
7629 => conv_std_logic_vector(23, 8),
7630 => conv_std_logic_vector(23, 8),
7631 => conv_std_logic_vector(23, 8),
7632 => conv_std_logic_vector(23, 8),
7633 => conv_std_logic_vector(23, 8),
7634 => conv_std_logic_vector(23, 8),
7635 => conv_std_logic_vector(23, 8),
7636 => conv_std_logic_vector(24, 8),
7637 => conv_std_logic_vector(24, 8),
7638 => conv_std_logic_vector(24, 8),
7639 => conv_std_logic_vector(24, 8),
7640 => conv_std_logic_vector(24, 8),
7641 => conv_std_logic_vector(24, 8),
7642 => conv_std_logic_vector(24, 8),
7643 => conv_std_logic_vector(24, 8),
7644 => conv_std_logic_vector(24, 8),
7645 => conv_std_logic_vector(25, 8),
7646 => conv_std_logic_vector(25, 8),
7647 => conv_std_logic_vector(25, 8),
7648 => conv_std_logic_vector(25, 8),
7649 => conv_std_logic_vector(25, 8),
7650 => conv_std_logic_vector(25, 8),
7651 => conv_std_logic_vector(25, 8),
7652 => conv_std_logic_vector(25, 8),
7653 => conv_std_logic_vector(25, 8),
7654 => conv_std_logic_vector(26, 8),
7655 => conv_std_logic_vector(26, 8),
7656 => conv_std_logic_vector(26, 8),
7657 => conv_std_logic_vector(26, 8),
7658 => conv_std_logic_vector(26, 8),
7659 => conv_std_logic_vector(26, 8),
7660 => conv_std_logic_vector(26, 8),
7661 => conv_std_logic_vector(26, 8),
7662 => conv_std_logic_vector(26, 8),
7663 => conv_std_logic_vector(27, 8),
7664 => conv_std_logic_vector(27, 8),
7665 => conv_std_logic_vector(27, 8),
7666 => conv_std_logic_vector(27, 8),
7667 => conv_std_logic_vector(27, 8),
7668 => conv_std_logic_vector(27, 8),
7669 => conv_std_logic_vector(27, 8),
7670 => conv_std_logic_vector(27, 8),
7671 => conv_std_logic_vector(27, 8),
7672 => conv_std_logic_vector(28, 8),
7673 => conv_std_logic_vector(28, 8),
7674 => conv_std_logic_vector(28, 8),
7675 => conv_std_logic_vector(28, 8),
7676 => conv_std_logic_vector(28, 8),
7677 => conv_std_logic_vector(28, 8),
7678 => conv_std_logic_vector(28, 8),
7679 => conv_std_logic_vector(28, 8),
7680 => conv_std_logic_vector(0, 8),
7681 => conv_std_logic_vector(0, 8),
7682 => conv_std_logic_vector(0, 8),
7683 => conv_std_logic_vector(0, 8),
7684 => conv_std_logic_vector(0, 8),
7685 => conv_std_logic_vector(0, 8),
7686 => conv_std_logic_vector(0, 8),
7687 => conv_std_logic_vector(0, 8),
7688 => conv_std_logic_vector(0, 8),
7689 => conv_std_logic_vector(1, 8),
7690 => conv_std_logic_vector(1, 8),
7691 => conv_std_logic_vector(1, 8),
7692 => conv_std_logic_vector(1, 8),
7693 => conv_std_logic_vector(1, 8),
7694 => conv_std_logic_vector(1, 8),
7695 => conv_std_logic_vector(1, 8),
7696 => conv_std_logic_vector(1, 8),
7697 => conv_std_logic_vector(1, 8),
7698 => conv_std_logic_vector(2, 8),
7699 => conv_std_logic_vector(2, 8),
7700 => conv_std_logic_vector(2, 8),
7701 => conv_std_logic_vector(2, 8),
7702 => conv_std_logic_vector(2, 8),
7703 => conv_std_logic_vector(2, 8),
7704 => conv_std_logic_vector(2, 8),
7705 => conv_std_logic_vector(2, 8),
7706 => conv_std_logic_vector(3, 8),
7707 => conv_std_logic_vector(3, 8),
7708 => conv_std_logic_vector(3, 8),
7709 => conv_std_logic_vector(3, 8),
7710 => conv_std_logic_vector(3, 8),
7711 => conv_std_logic_vector(3, 8),
7712 => conv_std_logic_vector(3, 8),
7713 => conv_std_logic_vector(3, 8),
7714 => conv_std_logic_vector(3, 8),
7715 => conv_std_logic_vector(4, 8),
7716 => conv_std_logic_vector(4, 8),
7717 => conv_std_logic_vector(4, 8),
7718 => conv_std_logic_vector(4, 8),
7719 => conv_std_logic_vector(4, 8),
7720 => conv_std_logic_vector(4, 8),
7721 => conv_std_logic_vector(4, 8),
7722 => conv_std_logic_vector(4, 8),
7723 => conv_std_logic_vector(5, 8),
7724 => conv_std_logic_vector(5, 8),
7725 => conv_std_logic_vector(5, 8),
7726 => conv_std_logic_vector(5, 8),
7727 => conv_std_logic_vector(5, 8),
7728 => conv_std_logic_vector(5, 8),
7729 => conv_std_logic_vector(5, 8),
7730 => conv_std_logic_vector(5, 8),
7731 => conv_std_logic_vector(5, 8),
7732 => conv_std_logic_vector(6, 8),
7733 => conv_std_logic_vector(6, 8),
7734 => conv_std_logic_vector(6, 8),
7735 => conv_std_logic_vector(6, 8),
7736 => conv_std_logic_vector(6, 8),
7737 => conv_std_logic_vector(6, 8),
7738 => conv_std_logic_vector(6, 8),
7739 => conv_std_logic_vector(6, 8),
7740 => conv_std_logic_vector(7, 8),
7741 => conv_std_logic_vector(7, 8),
7742 => conv_std_logic_vector(7, 8),
7743 => conv_std_logic_vector(7, 8),
7744 => conv_std_logic_vector(7, 8),
7745 => conv_std_logic_vector(7, 8),
7746 => conv_std_logic_vector(7, 8),
7747 => conv_std_logic_vector(7, 8),
7748 => conv_std_logic_vector(7, 8),
7749 => conv_std_logic_vector(8, 8),
7750 => conv_std_logic_vector(8, 8),
7751 => conv_std_logic_vector(8, 8),
7752 => conv_std_logic_vector(8, 8),
7753 => conv_std_logic_vector(8, 8),
7754 => conv_std_logic_vector(8, 8),
7755 => conv_std_logic_vector(8, 8),
7756 => conv_std_logic_vector(8, 8),
7757 => conv_std_logic_vector(9, 8),
7758 => conv_std_logic_vector(9, 8),
7759 => conv_std_logic_vector(9, 8),
7760 => conv_std_logic_vector(9, 8),
7761 => conv_std_logic_vector(9, 8),
7762 => conv_std_logic_vector(9, 8),
7763 => conv_std_logic_vector(9, 8),
7764 => conv_std_logic_vector(9, 8),
7765 => conv_std_logic_vector(9, 8),
7766 => conv_std_logic_vector(10, 8),
7767 => conv_std_logic_vector(10, 8),
7768 => conv_std_logic_vector(10, 8),
7769 => conv_std_logic_vector(10, 8),
7770 => conv_std_logic_vector(10, 8),
7771 => conv_std_logic_vector(10, 8),
7772 => conv_std_logic_vector(10, 8),
7773 => conv_std_logic_vector(10, 8),
7774 => conv_std_logic_vector(11, 8),
7775 => conv_std_logic_vector(11, 8),
7776 => conv_std_logic_vector(11, 8),
7777 => conv_std_logic_vector(11, 8),
7778 => conv_std_logic_vector(11, 8),
7779 => conv_std_logic_vector(11, 8),
7780 => conv_std_logic_vector(11, 8),
7781 => conv_std_logic_vector(11, 8),
7782 => conv_std_logic_vector(11, 8),
7783 => conv_std_logic_vector(12, 8),
7784 => conv_std_logic_vector(12, 8),
7785 => conv_std_logic_vector(12, 8),
7786 => conv_std_logic_vector(12, 8),
7787 => conv_std_logic_vector(12, 8),
7788 => conv_std_logic_vector(12, 8),
7789 => conv_std_logic_vector(12, 8),
7790 => conv_std_logic_vector(12, 8),
7791 => conv_std_logic_vector(13, 8),
7792 => conv_std_logic_vector(13, 8),
7793 => conv_std_logic_vector(13, 8),
7794 => conv_std_logic_vector(13, 8),
7795 => conv_std_logic_vector(13, 8),
7796 => conv_std_logic_vector(13, 8),
7797 => conv_std_logic_vector(13, 8),
7798 => conv_std_logic_vector(13, 8),
7799 => conv_std_logic_vector(13, 8),
7800 => conv_std_logic_vector(14, 8),
7801 => conv_std_logic_vector(14, 8),
7802 => conv_std_logic_vector(14, 8),
7803 => conv_std_logic_vector(14, 8),
7804 => conv_std_logic_vector(14, 8),
7805 => conv_std_logic_vector(14, 8),
7806 => conv_std_logic_vector(14, 8),
7807 => conv_std_logic_vector(14, 8),
7808 => conv_std_logic_vector(15, 8),
7809 => conv_std_logic_vector(15, 8),
7810 => conv_std_logic_vector(15, 8),
7811 => conv_std_logic_vector(15, 8),
7812 => conv_std_logic_vector(15, 8),
7813 => conv_std_logic_vector(15, 8),
7814 => conv_std_logic_vector(15, 8),
7815 => conv_std_logic_vector(15, 8),
7816 => conv_std_logic_vector(15, 8),
7817 => conv_std_logic_vector(16, 8),
7818 => conv_std_logic_vector(16, 8),
7819 => conv_std_logic_vector(16, 8),
7820 => conv_std_logic_vector(16, 8),
7821 => conv_std_logic_vector(16, 8),
7822 => conv_std_logic_vector(16, 8),
7823 => conv_std_logic_vector(16, 8),
7824 => conv_std_logic_vector(16, 8),
7825 => conv_std_logic_vector(16, 8),
7826 => conv_std_logic_vector(17, 8),
7827 => conv_std_logic_vector(17, 8),
7828 => conv_std_logic_vector(17, 8),
7829 => conv_std_logic_vector(17, 8),
7830 => conv_std_logic_vector(17, 8),
7831 => conv_std_logic_vector(17, 8),
7832 => conv_std_logic_vector(17, 8),
7833 => conv_std_logic_vector(17, 8),
7834 => conv_std_logic_vector(18, 8),
7835 => conv_std_logic_vector(18, 8),
7836 => conv_std_logic_vector(18, 8),
7837 => conv_std_logic_vector(18, 8),
7838 => conv_std_logic_vector(18, 8),
7839 => conv_std_logic_vector(18, 8),
7840 => conv_std_logic_vector(18, 8),
7841 => conv_std_logic_vector(18, 8),
7842 => conv_std_logic_vector(18, 8),
7843 => conv_std_logic_vector(19, 8),
7844 => conv_std_logic_vector(19, 8),
7845 => conv_std_logic_vector(19, 8),
7846 => conv_std_logic_vector(19, 8),
7847 => conv_std_logic_vector(19, 8),
7848 => conv_std_logic_vector(19, 8),
7849 => conv_std_logic_vector(19, 8),
7850 => conv_std_logic_vector(19, 8),
7851 => conv_std_logic_vector(20, 8),
7852 => conv_std_logic_vector(20, 8),
7853 => conv_std_logic_vector(20, 8),
7854 => conv_std_logic_vector(20, 8),
7855 => conv_std_logic_vector(20, 8),
7856 => conv_std_logic_vector(20, 8),
7857 => conv_std_logic_vector(20, 8),
7858 => conv_std_logic_vector(20, 8),
7859 => conv_std_logic_vector(20, 8),
7860 => conv_std_logic_vector(21, 8),
7861 => conv_std_logic_vector(21, 8),
7862 => conv_std_logic_vector(21, 8),
7863 => conv_std_logic_vector(21, 8),
7864 => conv_std_logic_vector(21, 8),
7865 => conv_std_logic_vector(21, 8),
7866 => conv_std_logic_vector(21, 8),
7867 => conv_std_logic_vector(21, 8),
7868 => conv_std_logic_vector(22, 8),
7869 => conv_std_logic_vector(22, 8),
7870 => conv_std_logic_vector(22, 8),
7871 => conv_std_logic_vector(22, 8),
7872 => conv_std_logic_vector(22, 8),
7873 => conv_std_logic_vector(22, 8),
7874 => conv_std_logic_vector(22, 8),
7875 => conv_std_logic_vector(22, 8),
7876 => conv_std_logic_vector(22, 8),
7877 => conv_std_logic_vector(23, 8),
7878 => conv_std_logic_vector(23, 8),
7879 => conv_std_logic_vector(23, 8),
7880 => conv_std_logic_vector(23, 8),
7881 => conv_std_logic_vector(23, 8),
7882 => conv_std_logic_vector(23, 8),
7883 => conv_std_logic_vector(23, 8),
7884 => conv_std_logic_vector(23, 8),
7885 => conv_std_logic_vector(24, 8),
7886 => conv_std_logic_vector(24, 8),
7887 => conv_std_logic_vector(24, 8),
7888 => conv_std_logic_vector(24, 8),
7889 => conv_std_logic_vector(24, 8),
7890 => conv_std_logic_vector(24, 8),
7891 => conv_std_logic_vector(24, 8),
7892 => conv_std_logic_vector(24, 8),
7893 => conv_std_logic_vector(24, 8),
7894 => conv_std_logic_vector(25, 8),
7895 => conv_std_logic_vector(25, 8),
7896 => conv_std_logic_vector(25, 8),
7897 => conv_std_logic_vector(25, 8),
7898 => conv_std_logic_vector(25, 8),
7899 => conv_std_logic_vector(25, 8),
7900 => conv_std_logic_vector(25, 8),
7901 => conv_std_logic_vector(25, 8),
7902 => conv_std_logic_vector(26, 8),
7903 => conv_std_logic_vector(26, 8),
7904 => conv_std_logic_vector(26, 8),
7905 => conv_std_logic_vector(26, 8),
7906 => conv_std_logic_vector(26, 8),
7907 => conv_std_logic_vector(26, 8),
7908 => conv_std_logic_vector(26, 8),
7909 => conv_std_logic_vector(26, 8),
7910 => conv_std_logic_vector(26, 8),
7911 => conv_std_logic_vector(27, 8),
7912 => conv_std_logic_vector(27, 8),
7913 => conv_std_logic_vector(27, 8),
7914 => conv_std_logic_vector(27, 8),
7915 => conv_std_logic_vector(27, 8),
7916 => conv_std_logic_vector(27, 8),
7917 => conv_std_logic_vector(27, 8),
7918 => conv_std_logic_vector(27, 8),
7919 => conv_std_logic_vector(28, 8),
7920 => conv_std_logic_vector(28, 8),
7921 => conv_std_logic_vector(28, 8),
7922 => conv_std_logic_vector(28, 8),
7923 => conv_std_logic_vector(28, 8),
7924 => conv_std_logic_vector(28, 8),
7925 => conv_std_logic_vector(28, 8),
7926 => conv_std_logic_vector(28, 8),
7927 => conv_std_logic_vector(28, 8),
7928 => conv_std_logic_vector(29, 8),
7929 => conv_std_logic_vector(29, 8),
7930 => conv_std_logic_vector(29, 8),
7931 => conv_std_logic_vector(29, 8),
7932 => conv_std_logic_vector(29, 8),
7933 => conv_std_logic_vector(29, 8),
7934 => conv_std_logic_vector(29, 8),
7935 => conv_std_logic_vector(29, 8),
7936 => conv_std_logic_vector(0, 8),
7937 => conv_std_logic_vector(0, 8),
7938 => conv_std_logic_vector(0, 8),
7939 => conv_std_logic_vector(0, 8),
7940 => conv_std_logic_vector(0, 8),
7941 => conv_std_logic_vector(0, 8),
7942 => conv_std_logic_vector(0, 8),
7943 => conv_std_logic_vector(0, 8),
7944 => conv_std_logic_vector(0, 8),
7945 => conv_std_logic_vector(1, 8),
7946 => conv_std_logic_vector(1, 8),
7947 => conv_std_logic_vector(1, 8),
7948 => conv_std_logic_vector(1, 8),
7949 => conv_std_logic_vector(1, 8),
7950 => conv_std_logic_vector(1, 8),
7951 => conv_std_logic_vector(1, 8),
7952 => conv_std_logic_vector(1, 8),
7953 => conv_std_logic_vector(2, 8),
7954 => conv_std_logic_vector(2, 8),
7955 => conv_std_logic_vector(2, 8),
7956 => conv_std_logic_vector(2, 8),
7957 => conv_std_logic_vector(2, 8),
7958 => conv_std_logic_vector(2, 8),
7959 => conv_std_logic_vector(2, 8),
7960 => conv_std_logic_vector(2, 8),
7961 => conv_std_logic_vector(3, 8),
7962 => conv_std_logic_vector(3, 8),
7963 => conv_std_logic_vector(3, 8),
7964 => conv_std_logic_vector(3, 8),
7965 => conv_std_logic_vector(3, 8),
7966 => conv_std_logic_vector(3, 8),
7967 => conv_std_logic_vector(3, 8),
7968 => conv_std_logic_vector(3, 8),
7969 => conv_std_logic_vector(3, 8),
7970 => conv_std_logic_vector(4, 8),
7971 => conv_std_logic_vector(4, 8),
7972 => conv_std_logic_vector(4, 8),
7973 => conv_std_logic_vector(4, 8),
7974 => conv_std_logic_vector(4, 8),
7975 => conv_std_logic_vector(4, 8),
7976 => conv_std_logic_vector(4, 8),
7977 => conv_std_logic_vector(4, 8),
7978 => conv_std_logic_vector(5, 8),
7979 => conv_std_logic_vector(5, 8),
7980 => conv_std_logic_vector(5, 8),
7981 => conv_std_logic_vector(5, 8),
7982 => conv_std_logic_vector(5, 8),
7983 => conv_std_logic_vector(5, 8),
7984 => conv_std_logic_vector(5, 8),
7985 => conv_std_logic_vector(5, 8),
7986 => conv_std_logic_vector(6, 8),
7987 => conv_std_logic_vector(6, 8),
7988 => conv_std_logic_vector(6, 8),
7989 => conv_std_logic_vector(6, 8),
7990 => conv_std_logic_vector(6, 8),
7991 => conv_std_logic_vector(6, 8),
7992 => conv_std_logic_vector(6, 8),
7993 => conv_std_logic_vector(6, 8),
7994 => conv_std_logic_vector(7, 8),
7995 => conv_std_logic_vector(7, 8),
7996 => conv_std_logic_vector(7, 8),
7997 => conv_std_logic_vector(7, 8),
7998 => conv_std_logic_vector(7, 8),
7999 => conv_std_logic_vector(7, 8),
8000 => conv_std_logic_vector(7, 8),
8001 => conv_std_logic_vector(7, 8),
8002 => conv_std_logic_vector(7, 8),
8003 => conv_std_logic_vector(8, 8),
8004 => conv_std_logic_vector(8, 8),
8005 => conv_std_logic_vector(8, 8),
8006 => conv_std_logic_vector(8, 8),
8007 => conv_std_logic_vector(8, 8),
8008 => conv_std_logic_vector(8, 8),
8009 => conv_std_logic_vector(8, 8),
8010 => conv_std_logic_vector(8, 8),
8011 => conv_std_logic_vector(9, 8),
8012 => conv_std_logic_vector(9, 8),
8013 => conv_std_logic_vector(9, 8),
8014 => conv_std_logic_vector(9, 8),
8015 => conv_std_logic_vector(9, 8),
8016 => conv_std_logic_vector(9, 8),
8017 => conv_std_logic_vector(9, 8),
8018 => conv_std_logic_vector(9, 8),
8019 => conv_std_logic_vector(10, 8),
8020 => conv_std_logic_vector(10, 8),
8021 => conv_std_logic_vector(10, 8),
8022 => conv_std_logic_vector(10, 8),
8023 => conv_std_logic_vector(10, 8),
8024 => conv_std_logic_vector(10, 8),
8025 => conv_std_logic_vector(10, 8),
8026 => conv_std_logic_vector(10, 8),
8027 => conv_std_logic_vector(11, 8),
8028 => conv_std_logic_vector(11, 8),
8029 => conv_std_logic_vector(11, 8),
8030 => conv_std_logic_vector(11, 8),
8031 => conv_std_logic_vector(11, 8),
8032 => conv_std_logic_vector(11, 8),
8033 => conv_std_logic_vector(11, 8),
8034 => conv_std_logic_vector(11, 8),
8035 => conv_std_logic_vector(11, 8),
8036 => conv_std_logic_vector(12, 8),
8037 => conv_std_logic_vector(12, 8),
8038 => conv_std_logic_vector(12, 8),
8039 => conv_std_logic_vector(12, 8),
8040 => conv_std_logic_vector(12, 8),
8041 => conv_std_logic_vector(12, 8),
8042 => conv_std_logic_vector(12, 8),
8043 => conv_std_logic_vector(12, 8),
8044 => conv_std_logic_vector(13, 8),
8045 => conv_std_logic_vector(13, 8),
8046 => conv_std_logic_vector(13, 8),
8047 => conv_std_logic_vector(13, 8),
8048 => conv_std_logic_vector(13, 8),
8049 => conv_std_logic_vector(13, 8),
8050 => conv_std_logic_vector(13, 8),
8051 => conv_std_logic_vector(13, 8),
8052 => conv_std_logic_vector(14, 8),
8053 => conv_std_logic_vector(14, 8),
8054 => conv_std_logic_vector(14, 8),
8055 => conv_std_logic_vector(14, 8),
8056 => conv_std_logic_vector(14, 8),
8057 => conv_std_logic_vector(14, 8),
8058 => conv_std_logic_vector(14, 8),
8059 => conv_std_logic_vector(14, 8),
8060 => conv_std_logic_vector(15, 8),
8061 => conv_std_logic_vector(15, 8),
8062 => conv_std_logic_vector(15, 8),
8063 => conv_std_logic_vector(15, 8),
8064 => conv_std_logic_vector(15, 8),
8065 => conv_std_logic_vector(15, 8),
8066 => conv_std_logic_vector(15, 8),
8067 => conv_std_logic_vector(15, 8),
8068 => conv_std_logic_vector(15, 8),
8069 => conv_std_logic_vector(16, 8),
8070 => conv_std_logic_vector(16, 8),
8071 => conv_std_logic_vector(16, 8),
8072 => conv_std_logic_vector(16, 8),
8073 => conv_std_logic_vector(16, 8),
8074 => conv_std_logic_vector(16, 8),
8075 => conv_std_logic_vector(16, 8),
8076 => conv_std_logic_vector(16, 8),
8077 => conv_std_logic_vector(17, 8),
8078 => conv_std_logic_vector(17, 8),
8079 => conv_std_logic_vector(17, 8),
8080 => conv_std_logic_vector(17, 8),
8081 => conv_std_logic_vector(17, 8),
8082 => conv_std_logic_vector(17, 8),
8083 => conv_std_logic_vector(17, 8),
8084 => conv_std_logic_vector(17, 8),
8085 => conv_std_logic_vector(18, 8),
8086 => conv_std_logic_vector(18, 8),
8087 => conv_std_logic_vector(18, 8),
8088 => conv_std_logic_vector(18, 8),
8089 => conv_std_logic_vector(18, 8),
8090 => conv_std_logic_vector(18, 8),
8091 => conv_std_logic_vector(18, 8),
8092 => conv_std_logic_vector(18, 8),
8093 => conv_std_logic_vector(19, 8),
8094 => conv_std_logic_vector(19, 8),
8095 => conv_std_logic_vector(19, 8),
8096 => conv_std_logic_vector(19, 8),
8097 => conv_std_logic_vector(19, 8),
8098 => conv_std_logic_vector(19, 8),
8099 => conv_std_logic_vector(19, 8),
8100 => conv_std_logic_vector(19, 8),
8101 => conv_std_logic_vector(19, 8),
8102 => conv_std_logic_vector(20, 8),
8103 => conv_std_logic_vector(20, 8),
8104 => conv_std_logic_vector(20, 8),
8105 => conv_std_logic_vector(20, 8),
8106 => conv_std_logic_vector(20, 8),
8107 => conv_std_logic_vector(20, 8),
8108 => conv_std_logic_vector(20, 8),
8109 => conv_std_logic_vector(20, 8),
8110 => conv_std_logic_vector(21, 8),
8111 => conv_std_logic_vector(21, 8),
8112 => conv_std_logic_vector(21, 8),
8113 => conv_std_logic_vector(21, 8),
8114 => conv_std_logic_vector(21, 8),
8115 => conv_std_logic_vector(21, 8),
8116 => conv_std_logic_vector(21, 8),
8117 => conv_std_logic_vector(21, 8),
8118 => conv_std_logic_vector(22, 8),
8119 => conv_std_logic_vector(22, 8),
8120 => conv_std_logic_vector(22, 8),
8121 => conv_std_logic_vector(22, 8),
8122 => conv_std_logic_vector(22, 8),
8123 => conv_std_logic_vector(22, 8),
8124 => conv_std_logic_vector(22, 8),
8125 => conv_std_logic_vector(22, 8),
8126 => conv_std_logic_vector(23, 8),
8127 => conv_std_logic_vector(23, 8),
8128 => conv_std_logic_vector(23, 8),
8129 => conv_std_logic_vector(23, 8),
8130 => conv_std_logic_vector(23, 8),
8131 => conv_std_logic_vector(23, 8),
8132 => conv_std_logic_vector(23, 8),
8133 => conv_std_logic_vector(23, 8),
8134 => conv_std_logic_vector(23, 8),
8135 => conv_std_logic_vector(24, 8),
8136 => conv_std_logic_vector(24, 8),
8137 => conv_std_logic_vector(24, 8),
8138 => conv_std_logic_vector(24, 8),
8139 => conv_std_logic_vector(24, 8),
8140 => conv_std_logic_vector(24, 8),
8141 => conv_std_logic_vector(24, 8),
8142 => conv_std_logic_vector(24, 8),
8143 => conv_std_logic_vector(25, 8),
8144 => conv_std_logic_vector(25, 8),
8145 => conv_std_logic_vector(25, 8),
8146 => conv_std_logic_vector(25, 8),
8147 => conv_std_logic_vector(25, 8),
8148 => conv_std_logic_vector(25, 8),
8149 => conv_std_logic_vector(25, 8),
8150 => conv_std_logic_vector(25, 8),
8151 => conv_std_logic_vector(26, 8),
8152 => conv_std_logic_vector(26, 8),
8153 => conv_std_logic_vector(26, 8),
8154 => conv_std_logic_vector(26, 8),
8155 => conv_std_logic_vector(26, 8),
8156 => conv_std_logic_vector(26, 8),
8157 => conv_std_logic_vector(26, 8),
8158 => conv_std_logic_vector(26, 8),
8159 => conv_std_logic_vector(27, 8),
8160 => conv_std_logic_vector(27, 8),
8161 => conv_std_logic_vector(27, 8),
8162 => conv_std_logic_vector(27, 8),
8163 => conv_std_logic_vector(27, 8),
8164 => conv_std_logic_vector(27, 8),
8165 => conv_std_logic_vector(27, 8),
8166 => conv_std_logic_vector(27, 8),
8167 => conv_std_logic_vector(27, 8),
8168 => conv_std_logic_vector(28, 8),
8169 => conv_std_logic_vector(28, 8),
8170 => conv_std_logic_vector(28, 8),
8171 => conv_std_logic_vector(28, 8),
8172 => conv_std_logic_vector(28, 8),
8173 => conv_std_logic_vector(28, 8),
8174 => conv_std_logic_vector(28, 8),
8175 => conv_std_logic_vector(28, 8),
8176 => conv_std_logic_vector(29, 8),
8177 => conv_std_logic_vector(29, 8),
8178 => conv_std_logic_vector(29, 8),
8179 => conv_std_logic_vector(29, 8),
8180 => conv_std_logic_vector(29, 8),
8181 => conv_std_logic_vector(29, 8),
8182 => conv_std_logic_vector(29, 8),
8183 => conv_std_logic_vector(29, 8),
8184 => conv_std_logic_vector(30, 8),
8185 => conv_std_logic_vector(30, 8),
8186 => conv_std_logic_vector(30, 8),
8187 => conv_std_logic_vector(30, 8),
8188 => conv_std_logic_vector(30, 8),
8189 => conv_std_logic_vector(30, 8),
8190 => conv_std_logic_vector(30, 8),
8191 => conv_std_logic_vector(30, 8),
8192 => conv_std_logic_vector(0, 8),
8193 => conv_std_logic_vector(0, 8),
8194 => conv_std_logic_vector(0, 8),
8195 => conv_std_logic_vector(0, 8),
8196 => conv_std_logic_vector(0, 8),
8197 => conv_std_logic_vector(0, 8),
8198 => conv_std_logic_vector(0, 8),
8199 => conv_std_logic_vector(0, 8),
8200 => conv_std_logic_vector(1, 8),
8201 => conv_std_logic_vector(1, 8),
8202 => conv_std_logic_vector(1, 8),
8203 => conv_std_logic_vector(1, 8),
8204 => conv_std_logic_vector(1, 8),
8205 => conv_std_logic_vector(1, 8),
8206 => conv_std_logic_vector(1, 8),
8207 => conv_std_logic_vector(1, 8),
8208 => conv_std_logic_vector(2, 8),
8209 => conv_std_logic_vector(2, 8),
8210 => conv_std_logic_vector(2, 8),
8211 => conv_std_logic_vector(2, 8),
8212 => conv_std_logic_vector(2, 8),
8213 => conv_std_logic_vector(2, 8),
8214 => conv_std_logic_vector(2, 8),
8215 => conv_std_logic_vector(2, 8),
8216 => conv_std_logic_vector(3, 8),
8217 => conv_std_logic_vector(3, 8),
8218 => conv_std_logic_vector(3, 8),
8219 => conv_std_logic_vector(3, 8),
8220 => conv_std_logic_vector(3, 8),
8221 => conv_std_logic_vector(3, 8),
8222 => conv_std_logic_vector(3, 8),
8223 => conv_std_logic_vector(3, 8),
8224 => conv_std_logic_vector(4, 8),
8225 => conv_std_logic_vector(4, 8),
8226 => conv_std_logic_vector(4, 8),
8227 => conv_std_logic_vector(4, 8),
8228 => conv_std_logic_vector(4, 8),
8229 => conv_std_logic_vector(4, 8),
8230 => conv_std_logic_vector(4, 8),
8231 => conv_std_logic_vector(4, 8),
8232 => conv_std_logic_vector(5, 8),
8233 => conv_std_logic_vector(5, 8),
8234 => conv_std_logic_vector(5, 8),
8235 => conv_std_logic_vector(5, 8),
8236 => conv_std_logic_vector(5, 8),
8237 => conv_std_logic_vector(5, 8),
8238 => conv_std_logic_vector(5, 8),
8239 => conv_std_logic_vector(5, 8),
8240 => conv_std_logic_vector(6, 8),
8241 => conv_std_logic_vector(6, 8),
8242 => conv_std_logic_vector(6, 8),
8243 => conv_std_logic_vector(6, 8),
8244 => conv_std_logic_vector(6, 8),
8245 => conv_std_logic_vector(6, 8),
8246 => conv_std_logic_vector(6, 8),
8247 => conv_std_logic_vector(6, 8),
8248 => conv_std_logic_vector(7, 8),
8249 => conv_std_logic_vector(7, 8),
8250 => conv_std_logic_vector(7, 8),
8251 => conv_std_logic_vector(7, 8),
8252 => conv_std_logic_vector(7, 8),
8253 => conv_std_logic_vector(7, 8),
8254 => conv_std_logic_vector(7, 8),
8255 => conv_std_logic_vector(7, 8),
8256 => conv_std_logic_vector(8, 8),
8257 => conv_std_logic_vector(8, 8),
8258 => conv_std_logic_vector(8, 8),
8259 => conv_std_logic_vector(8, 8),
8260 => conv_std_logic_vector(8, 8),
8261 => conv_std_logic_vector(8, 8),
8262 => conv_std_logic_vector(8, 8),
8263 => conv_std_logic_vector(8, 8),
8264 => conv_std_logic_vector(9, 8),
8265 => conv_std_logic_vector(9, 8),
8266 => conv_std_logic_vector(9, 8),
8267 => conv_std_logic_vector(9, 8),
8268 => conv_std_logic_vector(9, 8),
8269 => conv_std_logic_vector(9, 8),
8270 => conv_std_logic_vector(9, 8),
8271 => conv_std_logic_vector(9, 8),
8272 => conv_std_logic_vector(10, 8),
8273 => conv_std_logic_vector(10, 8),
8274 => conv_std_logic_vector(10, 8),
8275 => conv_std_logic_vector(10, 8),
8276 => conv_std_logic_vector(10, 8),
8277 => conv_std_logic_vector(10, 8),
8278 => conv_std_logic_vector(10, 8),
8279 => conv_std_logic_vector(10, 8),
8280 => conv_std_logic_vector(11, 8),
8281 => conv_std_logic_vector(11, 8),
8282 => conv_std_logic_vector(11, 8),
8283 => conv_std_logic_vector(11, 8),
8284 => conv_std_logic_vector(11, 8),
8285 => conv_std_logic_vector(11, 8),
8286 => conv_std_logic_vector(11, 8),
8287 => conv_std_logic_vector(11, 8),
8288 => conv_std_logic_vector(12, 8),
8289 => conv_std_logic_vector(12, 8),
8290 => conv_std_logic_vector(12, 8),
8291 => conv_std_logic_vector(12, 8),
8292 => conv_std_logic_vector(12, 8),
8293 => conv_std_logic_vector(12, 8),
8294 => conv_std_logic_vector(12, 8),
8295 => conv_std_logic_vector(12, 8),
8296 => conv_std_logic_vector(13, 8),
8297 => conv_std_logic_vector(13, 8),
8298 => conv_std_logic_vector(13, 8),
8299 => conv_std_logic_vector(13, 8),
8300 => conv_std_logic_vector(13, 8),
8301 => conv_std_logic_vector(13, 8),
8302 => conv_std_logic_vector(13, 8),
8303 => conv_std_logic_vector(13, 8),
8304 => conv_std_logic_vector(14, 8),
8305 => conv_std_logic_vector(14, 8),
8306 => conv_std_logic_vector(14, 8),
8307 => conv_std_logic_vector(14, 8),
8308 => conv_std_logic_vector(14, 8),
8309 => conv_std_logic_vector(14, 8),
8310 => conv_std_logic_vector(14, 8),
8311 => conv_std_logic_vector(14, 8),
8312 => conv_std_logic_vector(15, 8),
8313 => conv_std_logic_vector(15, 8),
8314 => conv_std_logic_vector(15, 8),
8315 => conv_std_logic_vector(15, 8),
8316 => conv_std_logic_vector(15, 8),
8317 => conv_std_logic_vector(15, 8),
8318 => conv_std_logic_vector(15, 8),
8319 => conv_std_logic_vector(15, 8),
8320 => conv_std_logic_vector(16, 8),
8321 => conv_std_logic_vector(16, 8),
8322 => conv_std_logic_vector(16, 8),
8323 => conv_std_logic_vector(16, 8),
8324 => conv_std_logic_vector(16, 8),
8325 => conv_std_logic_vector(16, 8),
8326 => conv_std_logic_vector(16, 8),
8327 => conv_std_logic_vector(16, 8),
8328 => conv_std_logic_vector(17, 8),
8329 => conv_std_logic_vector(17, 8),
8330 => conv_std_logic_vector(17, 8),
8331 => conv_std_logic_vector(17, 8),
8332 => conv_std_logic_vector(17, 8),
8333 => conv_std_logic_vector(17, 8),
8334 => conv_std_logic_vector(17, 8),
8335 => conv_std_logic_vector(17, 8),
8336 => conv_std_logic_vector(18, 8),
8337 => conv_std_logic_vector(18, 8),
8338 => conv_std_logic_vector(18, 8),
8339 => conv_std_logic_vector(18, 8),
8340 => conv_std_logic_vector(18, 8),
8341 => conv_std_logic_vector(18, 8),
8342 => conv_std_logic_vector(18, 8),
8343 => conv_std_logic_vector(18, 8),
8344 => conv_std_logic_vector(19, 8),
8345 => conv_std_logic_vector(19, 8),
8346 => conv_std_logic_vector(19, 8),
8347 => conv_std_logic_vector(19, 8),
8348 => conv_std_logic_vector(19, 8),
8349 => conv_std_logic_vector(19, 8),
8350 => conv_std_logic_vector(19, 8),
8351 => conv_std_logic_vector(19, 8),
8352 => conv_std_logic_vector(20, 8),
8353 => conv_std_logic_vector(20, 8),
8354 => conv_std_logic_vector(20, 8),
8355 => conv_std_logic_vector(20, 8),
8356 => conv_std_logic_vector(20, 8),
8357 => conv_std_logic_vector(20, 8),
8358 => conv_std_logic_vector(20, 8),
8359 => conv_std_logic_vector(20, 8),
8360 => conv_std_logic_vector(21, 8),
8361 => conv_std_logic_vector(21, 8),
8362 => conv_std_logic_vector(21, 8),
8363 => conv_std_logic_vector(21, 8),
8364 => conv_std_logic_vector(21, 8),
8365 => conv_std_logic_vector(21, 8),
8366 => conv_std_logic_vector(21, 8),
8367 => conv_std_logic_vector(21, 8),
8368 => conv_std_logic_vector(22, 8),
8369 => conv_std_logic_vector(22, 8),
8370 => conv_std_logic_vector(22, 8),
8371 => conv_std_logic_vector(22, 8),
8372 => conv_std_logic_vector(22, 8),
8373 => conv_std_logic_vector(22, 8),
8374 => conv_std_logic_vector(22, 8),
8375 => conv_std_logic_vector(22, 8),
8376 => conv_std_logic_vector(23, 8),
8377 => conv_std_logic_vector(23, 8),
8378 => conv_std_logic_vector(23, 8),
8379 => conv_std_logic_vector(23, 8),
8380 => conv_std_logic_vector(23, 8),
8381 => conv_std_logic_vector(23, 8),
8382 => conv_std_logic_vector(23, 8),
8383 => conv_std_logic_vector(23, 8),
8384 => conv_std_logic_vector(24, 8),
8385 => conv_std_logic_vector(24, 8),
8386 => conv_std_logic_vector(24, 8),
8387 => conv_std_logic_vector(24, 8),
8388 => conv_std_logic_vector(24, 8),
8389 => conv_std_logic_vector(24, 8),
8390 => conv_std_logic_vector(24, 8),
8391 => conv_std_logic_vector(24, 8),
8392 => conv_std_logic_vector(25, 8),
8393 => conv_std_logic_vector(25, 8),
8394 => conv_std_logic_vector(25, 8),
8395 => conv_std_logic_vector(25, 8),
8396 => conv_std_logic_vector(25, 8),
8397 => conv_std_logic_vector(25, 8),
8398 => conv_std_logic_vector(25, 8),
8399 => conv_std_logic_vector(25, 8),
8400 => conv_std_logic_vector(26, 8),
8401 => conv_std_logic_vector(26, 8),
8402 => conv_std_logic_vector(26, 8),
8403 => conv_std_logic_vector(26, 8),
8404 => conv_std_logic_vector(26, 8),
8405 => conv_std_logic_vector(26, 8),
8406 => conv_std_logic_vector(26, 8),
8407 => conv_std_logic_vector(26, 8),
8408 => conv_std_logic_vector(27, 8),
8409 => conv_std_logic_vector(27, 8),
8410 => conv_std_logic_vector(27, 8),
8411 => conv_std_logic_vector(27, 8),
8412 => conv_std_logic_vector(27, 8),
8413 => conv_std_logic_vector(27, 8),
8414 => conv_std_logic_vector(27, 8),
8415 => conv_std_logic_vector(27, 8),
8416 => conv_std_logic_vector(28, 8),
8417 => conv_std_logic_vector(28, 8),
8418 => conv_std_logic_vector(28, 8),
8419 => conv_std_logic_vector(28, 8),
8420 => conv_std_logic_vector(28, 8),
8421 => conv_std_logic_vector(28, 8),
8422 => conv_std_logic_vector(28, 8),
8423 => conv_std_logic_vector(28, 8),
8424 => conv_std_logic_vector(29, 8),
8425 => conv_std_logic_vector(29, 8),
8426 => conv_std_logic_vector(29, 8),
8427 => conv_std_logic_vector(29, 8),
8428 => conv_std_logic_vector(29, 8),
8429 => conv_std_logic_vector(29, 8),
8430 => conv_std_logic_vector(29, 8),
8431 => conv_std_logic_vector(29, 8),
8432 => conv_std_logic_vector(30, 8),
8433 => conv_std_logic_vector(30, 8),
8434 => conv_std_logic_vector(30, 8),
8435 => conv_std_logic_vector(30, 8),
8436 => conv_std_logic_vector(30, 8),
8437 => conv_std_logic_vector(30, 8),
8438 => conv_std_logic_vector(30, 8),
8439 => conv_std_logic_vector(30, 8),
8440 => conv_std_logic_vector(31, 8),
8441 => conv_std_logic_vector(31, 8),
8442 => conv_std_logic_vector(31, 8),
8443 => conv_std_logic_vector(31, 8),
8444 => conv_std_logic_vector(31, 8),
8445 => conv_std_logic_vector(31, 8),
8446 => conv_std_logic_vector(31, 8),
8447 => conv_std_logic_vector(31, 8),
8448 => conv_std_logic_vector(0, 8),
8449 => conv_std_logic_vector(0, 8),
8450 => conv_std_logic_vector(0, 8),
8451 => conv_std_logic_vector(0, 8),
8452 => conv_std_logic_vector(0, 8),
8453 => conv_std_logic_vector(0, 8),
8454 => conv_std_logic_vector(0, 8),
8455 => conv_std_logic_vector(0, 8),
8456 => conv_std_logic_vector(1, 8),
8457 => conv_std_logic_vector(1, 8),
8458 => conv_std_logic_vector(1, 8),
8459 => conv_std_logic_vector(1, 8),
8460 => conv_std_logic_vector(1, 8),
8461 => conv_std_logic_vector(1, 8),
8462 => conv_std_logic_vector(1, 8),
8463 => conv_std_logic_vector(1, 8),
8464 => conv_std_logic_vector(2, 8),
8465 => conv_std_logic_vector(2, 8),
8466 => conv_std_logic_vector(2, 8),
8467 => conv_std_logic_vector(2, 8),
8468 => conv_std_logic_vector(2, 8),
8469 => conv_std_logic_vector(2, 8),
8470 => conv_std_logic_vector(2, 8),
8471 => conv_std_logic_vector(2, 8),
8472 => conv_std_logic_vector(3, 8),
8473 => conv_std_logic_vector(3, 8),
8474 => conv_std_logic_vector(3, 8),
8475 => conv_std_logic_vector(3, 8),
8476 => conv_std_logic_vector(3, 8),
8477 => conv_std_logic_vector(3, 8),
8478 => conv_std_logic_vector(3, 8),
8479 => conv_std_logic_vector(3, 8),
8480 => conv_std_logic_vector(4, 8),
8481 => conv_std_logic_vector(4, 8),
8482 => conv_std_logic_vector(4, 8),
8483 => conv_std_logic_vector(4, 8),
8484 => conv_std_logic_vector(4, 8),
8485 => conv_std_logic_vector(4, 8),
8486 => conv_std_logic_vector(4, 8),
8487 => conv_std_logic_vector(5, 8),
8488 => conv_std_logic_vector(5, 8),
8489 => conv_std_logic_vector(5, 8),
8490 => conv_std_logic_vector(5, 8),
8491 => conv_std_logic_vector(5, 8),
8492 => conv_std_logic_vector(5, 8),
8493 => conv_std_logic_vector(5, 8),
8494 => conv_std_logic_vector(5, 8),
8495 => conv_std_logic_vector(6, 8),
8496 => conv_std_logic_vector(6, 8),
8497 => conv_std_logic_vector(6, 8),
8498 => conv_std_logic_vector(6, 8),
8499 => conv_std_logic_vector(6, 8),
8500 => conv_std_logic_vector(6, 8),
8501 => conv_std_logic_vector(6, 8),
8502 => conv_std_logic_vector(6, 8),
8503 => conv_std_logic_vector(7, 8),
8504 => conv_std_logic_vector(7, 8),
8505 => conv_std_logic_vector(7, 8),
8506 => conv_std_logic_vector(7, 8),
8507 => conv_std_logic_vector(7, 8),
8508 => conv_std_logic_vector(7, 8),
8509 => conv_std_logic_vector(7, 8),
8510 => conv_std_logic_vector(7, 8),
8511 => conv_std_logic_vector(8, 8),
8512 => conv_std_logic_vector(8, 8),
8513 => conv_std_logic_vector(8, 8),
8514 => conv_std_logic_vector(8, 8),
8515 => conv_std_logic_vector(8, 8),
8516 => conv_std_logic_vector(8, 8),
8517 => conv_std_logic_vector(8, 8),
8518 => conv_std_logic_vector(9, 8),
8519 => conv_std_logic_vector(9, 8),
8520 => conv_std_logic_vector(9, 8),
8521 => conv_std_logic_vector(9, 8),
8522 => conv_std_logic_vector(9, 8),
8523 => conv_std_logic_vector(9, 8),
8524 => conv_std_logic_vector(9, 8),
8525 => conv_std_logic_vector(9, 8),
8526 => conv_std_logic_vector(10, 8),
8527 => conv_std_logic_vector(10, 8),
8528 => conv_std_logic_vector(10, 8),
8529 => conv_std_logic_vector(10, 8),
8530 => conv_std_logic_vector(10, 8),
8531 => conv_std_logic_vector(10, 8),
8532 => conv_std_logic_vector(10, 8),
8533 => conv_std_logic_vector(10, 8),
8534 => conv_std_logic_vector(11, 8),
8535 => conv_std_logic_vector(11, 8),
8536 => conv_std_logic_vector(11, 8),
8537 => conv_std_logic_vector(11, 8),
8538 => conv_std_logic_vector(11, 8),
8539 => conv_std_logic_vector(11, 8),
8540 => conv_std_logic_vector(11, 8),
8541 => conv_std_logic_vector(11, 8),
8542 => conv_std_logic_vector(12, 8),
8543 => conv_std_logic_vector(12, 8),
8544 => conv_std_logic_vector(12, 8),
8545 => conv_std_logic_vector(12, 8),
8546 => conv_std_logic_vector(12, 8),
8547 => conv_std_logic_vector(12, 8),
8548 => conv_std_logic_vector(12, 8),
8549 => conv_std_logic_vector(13, 8),
8550 => conv_std_logic_vector(13, 8),
8551 => conv_std_logic_vector(13, 8),
8552 => conv_std_logic_vector(13, 8),
8553 => conv_std_logic_vector(13, 8),
8554 => conv_std_logic_vector(13, 8),
8555 => conv_std_logic_vector(13, 8),
8556 => conv_std_logic_vector(13, 8),
8557 => conv_std_logic_vector(14, 8),
8558 => conv_std_logic_vector(14, 8),
8559 => conv_std_logic_vector(14, 8),
8560 => conv_std_logic_vector(14, 8),
8561 => conv_std_logic_vector(14, 8),
8562 => conv_std_logic_vector(14, 8),
8563 => conv_std_logic_vector(14, 8),
8564 => conv_std_logic_vector(14, 8),
8565 => conv_std_logic_vector(15, 8),
8566 => conv_std_logic_vector(15, 8),
8567 => conv_std_logic_vector(15, 8),
8568 => conv_std_logic_vector(15, 8),
8569 => conv_std_logic_vector(15, 8),
8570 => conv_std_logic_vector(15, 8),
8571 => conv_std_logic_vector(15, 8),
8572 => conv_std_logic_vector(15, 8),
8573 => conv_std_logic_vector(16, 8),
8574 => conv_std_logic_vector(16, 8),
8575 => conv_std_logic_vector(16, 8),
8576 => conv_std_logic_vector(16, 8),
8577 => conv_std_logic_vector(16, 8),
8578 => conv_std_logic_vector(16, 8),
8579 => conv_std_logic_vector(16, 8),
8580 => conv_std_logic_vector(17, 8),
8581 => conv_std_logic_vector(17, 8),
8582 => conv_std_logic_vector(17, 8),
8583 => conv_std_logic_vector(17, 8),
8584 => conv_std_logic_vector(17, 8),
8585 => conv_std_logic_vector(17, 8),
8586 => conv_std_logic_vector(17, 8),
8587 => conv_std_logic_vector(17, 8),
8588 => conv_std_logic_vector(18, 8),
8589 => conv_std_logic_vector(18, 8),
8590 => conv_std_logic_vector(18, 8),
8591 => conv_std_logic_vector(18, 8),
8592 => conv_std_logic_vector(18, 8),
8593 => conv_std_logic_vector(18, 8),
8594 => conv_std_logic_vector(18, 8),
8595 => conv_std_logic_vector(18, 8),
8596 => conv_std_logic_vector(19, 8),
8597 => conv_std_logic_vector(19, 8),
8598 => conv_std_logic_vector(19, 8),
8599 => conv_std_logic_vector(19, 8),
8600 => conv_std_logic_vector(19, 8),
8601 => conv_std_logic_vector(19, 8),
8602 => conv_std_logic_vector(19, 8),
8603 => conv_std_logic_vector(19, 8),
8604 => conv_std_logic_vector(20, 8),
8605 => conv_std_logic_vector(20, 8),
8606 => conv_std_logic_vector(20, 8),
8607 => conv_std_logic_vector(20, 8),
8608 => conv_std_logic_vector(20, 8),
8609 => conv_std_logic_vector(20, 8),
8610 => conv_std_logic_vector(20, 8),
8611 => conv_std_logic_vector(21, 8),
8612 => conv_std_logic_vector(21, 8),
8613 => conv_std_logic_vector(21, 8),
8614 => conv_std_logic_vector(21, 8),
8615 => conv_std_logic_vector(21, 8),
8616 => conv_std_logic_vector(21, 8),
8617 => conv_std_logic_vector(21, 8),
8618 => conv_std_logic_vector(21, 8),
8619 => conv_std_logic_vector(22, 8),
8620 => conv_std_logic_vector(22, 8),
8621 => conv_std_logic_vector(22, 8),
8622 => conv_std_logic_vector(22, 8),
8623 => conv_std_logic_vector(22, 8),
8624 => conv_std_logic_vector(22, 8),
8625 => conv_std_logic_vector(22, 8),
8626 => conv_std_logic_vector(22, 8),
8627 => conv_std_logic_vector(23, 8),
8628 => conv_std_logic_vector(23, 8),
8629 => conv_std_logic_vector(23, 8),
8630 => conv_std_logic_vector(23, 8),
8631 => conv_std_logic_vector(23, 8),
8632 => conv_std_logic_vector(23, 8),
8633 => conv_std_logic_vector(23, 8),
8634 => conv_std_logic_vector(23, 8),
8635 => conv_std_logic_vector(24, 8),
8636 => conv_std_logic_vector(24, 8),
8637 => conv_std_logic_vector(24, 8),
8638 => conv_std_logic_vector(24, 8),
8639 => conv_std_logic_vector(24, 8),
8640 => conv_std_logic_vector(24, 8),
8641 => conv_std_logic_vector(24, 8),
8642 => conv_std_logic_vector(25, 8),
8643 => conv_std_logic_vector(25, 8),
8644 => conv_std_logic_vector(25, 8),
8645 => conv_std_logic_vector(25, 8),
8646 => conv_std_logic_vector(25, 8),
8647 => conv_std_logic_vector(25, 8),
8648 => conv_std_logic_vector(25, 8),
8649 => conv_std_logic_vector(25, 8),
8650 => conv_std_logic_vector(26, 8),
8651 => conv_std_logic_vector(26, 8),
8652 => conv_std_logic_vector(26, 8),
8653 => conv_std_logic_vector(26, 8),
8654 => conv_std_logic_vector(26, 8),
8655 => conv_std_logic_vector(26, 8),
8656 => conv_std_logic_vector(26, 8),
8657 => conv_std_logic_vector(26, 8),
8658 => conv_std_logic_vector(27, 8),
8659 => conv_std_logic_vector(27, 8),
8660 => conv_std_logic_vector(27, 8),
8661 => conv_std_logic_vector(27, 8),
8662 => conv_std_logic_vector(27, 8),
8663 => conv_std_logic_vector(27, 8),
8664 => conv_std_logic_vector(27, 8),
8665 => conv_std_logic_vector(27, 8),
8666 => conv_std_logic_vector(28, 8),
8667 => conv_std_logic_vector(28, 8),
8668 => conv_std_logic_vector(28, 8),
8669 => conv_std_logic_vector(28, 8),
8670 => conv_std_logic_vector(28, 8),
8671 => conv_std_logic_vector(28, 8),
8672 => conv_std_logic_vector(28, 8),
8673 => conv_std_logic_vector(29, 8),
8674 => conv_std_logic_vector(29, 8),
8675 => conv_std_logic_vector(29, 8),
8676 => conv_std_logic_vector(29, 8),
8677 => conv_std_logic_vector(29, 8),
8678 => conv_std_logic_vector(29, 8),
8679 => conv_std_logic_vector(29, 8),
8680 => conv_std_logic_vector(29, 8),
8681 => conv_std_logic_vector(30, 8),
8682 => conv_std_logic_vector(30, 8),
8683 => conv_std_logic_vector(30, 8),
8684 => conv_std_logic_vector(30, 8),
8685 => conv_std_logic_vector(30, 8),
8686 => conv_std_logic_vector(30, 8),
8687 => conv_std_logic_vector(30, 8),
8688 => conv_std_logic_vector(30, 8),
8689 => conv_std_logic_vector(31, 8),
8690 => conv_std_logic_vector(31, 8),
8691 => conv_std_logic_vector(31, 8),
8692 => conv_std_logic_vector(31, 8),
8693 => conv_std_logic_vector(31, 8),
8694 => conv_std_logic_vector(31, 8),
8695 => conv_std_logic_vector(31, 8),
8696 => conv_std_logic_vector(31, 8),
8697 => conv_std_logic_vector(32, 8),
8698 => conv_std_logic_vector(32, 8),
8699 => conv_std_logic_vector(32, 8),
8700 => conv_std_logic_vector(32, 8),
8701 => conv_std_logic_vector(32, 8),
8702 => conv_std_logic_vector(32, 8),
8703 => conv_std_logic_vector(32, 8),
8704 => conv_std_logic_vector(0, 8),
8705 => conv_std_logic_vector(0, 8),
8706 => conv_std_logic_vector(0, 8),
8707 => conv_std_logic_vector(0, 8),
8708 => conv_std_logic_vector(0, 8),
8709 => conv_std_logic_vector(0, 8),
8710 => conv_std_logic_vector(0, 8),
8711 => conv_std_logic_vector(0, 8),
8712 => conv_std_logic_vector(1, 8),
8713 => conv_std_logic_vector(1, 8),
8714 => conv_std_logic_vector(1, 8),
8715 => conv_std_logic_vector(1, 8),
8716 => conv_std_logic_vector(1, 8),
8717 => conv_std_logic_vector(1, 8),
8718 => conv_std_logic_vector(1, 8),
8719 => conv_std_logic_vector(1, 8),
8720 => conv_std_logic_vector(2, 8),
8721 => conv_std_logic_vector(2, 8),
8722 => conv_std_logic_vector(2, 8),
8723 => conv_std_logic_vector(2, 8),
8724 => conv_std_logic_vector(2, 8),
8725 => conv_std_logic_vector(2, 8),
8726 => conv_std_logic_vector(2, 8),
8727 => conv_std_logic_vector(3, 8),
8728 => conv_std_logic_vector(3, 8),
8729 => conv_std_logic_vector(3, 8),
8730 => conv_std_logic_vector(3, 8),
8731 => conv_std_logic_vector(3, 8),
8732 => conv_std_logic_vector(3, 8),
8733 => conv_std_logic_vector(3, 8),
8734 => conv_std_logic_vector(3, 8),
8735 => conv_std_logic_vector(4, 8),
8736 => conv_std_logic_vector(4, 8),
8737 => conv_std_logic_vector(4, 8),
8738 => conv_std_logic_vector(4, 8),
8739 => conv_std_logic_vector(4, 8),
8740 => conv_std_logic_vector(4, 8),
8741 => conv_std_logic_vector(4, 8),
8742 => conv_std_logic_vector(5, 8),
8743 => conv_std_logic_vector(5, 8),
8744 => conv_std_logic_vector(5, 8),
8745 => conv_std_logic_vector(5, 8),
8746 => conv_std_logic_vector(5, 8),
8747 => conv_std_logic_vector(5, 8),
8748 => conv_std_logic_vector(5, 8),
8749 => conv_std_logic_vector(5, 8),
8750 => conv_std_logic_vector(6, 8),
8751 => conv_std_logic_vector(6, 8),
8752 => conv_std_logic_vector(6, 8),
8753 => conv_std_logic_vector(6, 8),
8754 => conv_std_logic_vector(6, 8),
8755 => conv_std_logic_vector(6, 8),
8756 => conv_std_logic_vector(6, 8),
8757 => conv_std_logic_vector(7, 8),
8758 => conv_std_logic_vector(7, 8),
8759 => conv_std_logic_vector(7, 8),
8760 => conv_std_logic_vector(7, 8),
8761 => conv_std_logic_vector(7, 8),
8762 => conv_std_logic_vector(7, 8),
8763 => conv_std_logic_vector(7, 8),
8764 => conv_std_logic_vector(7, 8),
8765 => conv_std_logic_vector(8, 8),
8766 => conv_std_logic_vector(8, 8),
8767 => conv_std_logic_vector(8, 8),
8768 => conv_std_logic_vector(8, 8),
8769 => conv_std_logic_vector(8, 8),
8770 => conv_std_logic_vector(8, 8),
8771 => conv_std_logic_vector(8, 8),
8772 => conv_std_logic_vector(9, 8),
8773 => conv_std_logic_vector(9, 8),
8774 => conv_std_logic_vector(9, 8),
8775 => conv_std_logic_vector(9, 8),
8776 => conv_std_logic_vector(9, 8),
8777 => conv_std_logic_vector(9, 8),
8778 => conv_std_logic_vector(9, 8),
8779 => conv_std_logic_vector(9, 8),
8780 => conv_std_logic_vector(10, 8),
8781 => conv_std_logic_vector(10, 8),
8782 => conv_std_logic_vector(10, 8),
8783 => conv_std_logic_vector(10, 8),
8784 => conv_std_logic_vector(10, 8),
8785 => conv_std_logic_vector(10, 8),
8786 => conv_std_logic_vector(10, 8),
8787 => conv_std_logic_vector(11, 8),
8788 => conv_std_logic_vector(11, 8),
8789 => conv_std_logic_vector(11, 8),
8790 => conv_std_logic_vector(11, 8),
8791 => conv_std_logic_vector(11, 8),
8792 => conv_std_logic_vector(11, 8),
8793 => conv_std_logic_vector(11, 8),
8794 => conv_std_logic_vector(11, 8),
8795 => conv_std_logic_vector(12, 8),
8796 => conv_std_logic_vector(12, 8),
8797 => conv_std_logic_vector(12, 8),
8798 => conv_std_logic_vector(12, 8),
8799 => conv_std_logic_vector(12, 8),
8800 => conv_std_logic_vector(12, 8),
8801 => conv_std_logic_vector(12, 8),
8802 => conv_std_logic_vector(13, 8),
8803 => conv_std_logic_vector(13, 8),
8804 => conv_std_logic_vector(13, 8),
8805 => conv_std_logic_vector(13, 8),
8806 => conv_std_logic_vector(13, 8),
8807 => conv_std_logic_vector(13, 8),
8808 => conv_std_logic_vector(13, 8),
8809 => conv_std_logic_vector(13, 8),
8810 => conv_std_logic_vector(14, 8),
8811 => conv_std_logic_vector(14, 8),
8812 => conv_std_logic_vector(14, 8),
8813 => conv_std_logic_vector(14, 8),
8814 => conv_std_logic_vector(14, 8),
8815 => conv_std_logic_vector(14, 8),
8816 => conv_std_logic_vector(14, 8),
8817 => conv_std_logic_vector(15, 8),
8818 => conv_std_logic_vector(15, 8),
8819 => conv_std_logic_vector(15, 8),
8820 => conv_std_logic_vector(15, 8),
8821 => conv_std_logic_vector(15, 8),
8822 => conv_std_logic_vector(15, 8),
8823 => conv_std_logic_vector(15, 8),
8824 => conv_std_logic_vector(15, 8),
8825 => conv_std_logic_vector(16, 8),
8826 => conv_std_logic_vector(16, 8),
8827 => conv_std_logic_vector(16, 8),
8828 => conv_std_logic_vector(16, 8),
8829 => conv_std_logic_vector(16, 8),
8830 => conv_std_logic_vector(16, 8),
8831 => conv_std_logic_vector(16, 8),
8832 => conv_std_logic_vector(17, 8),
8833 => conv_std_logic_vector(17, 8),
8834 => conv_std_logic_vector(17, 8),
8835 => conv_std_logic_vector(17, 8),
8836 => conv_std_logic_vector(17, 8),
8837 => conv_std_logic_vector(17, 8),
8838 => conv_std_logic_vector(17, 8),
8839 => conv_std_logic_vector(17, 8),
8840 => conv_std_logic_vector(18, 8),
8841 => conv_std_logic_vector(18, 8),
8842 => conv_std_logic_vector(18, 8),
8843 => conv_std_logic_vector(18, 8),
8844 => conv_std_logic_vector(18, 8),
8845 => conv_std_logic_vector(18, 8),
8846 => conv_std_logic_vector(18, 8),
8847 => conv_std_logic_vector(18, 8),
8848 => conv_std_logic_vector(19, 8),
8849 => conv_std_logic_vector(19, 8),
8850 => conv_std_logic_vector(19, 8),
8851 => conv_std_logic_vector(19, 8),
8852 => conv_std_logic_vector(19, 8),
8853 => conv_std_logic_vector(19, 8),
8854 => conv_std_logic_vector(19, 8),
8855 => conv_std_logic_vector(20, 8),
8856 => conv_std_logic_vector(20, 8),
8857 => conv_std_logic_vector(20, 8),
8858 => conv_std_logic_vector(20, 8),
8859 => conv_std_logic_vector(20, 8),
8860 => conv_std_logic_vector(20, 8),
8861 => conv_std_logic_vector(20, 8),
8862 => conv_std_logic_vector(20, 8),
8863 => conv_std_logic_vector(21, 8),
8864 => conv_std_logic_vector(21, 8),
8865 => conv_std_logic_vector(21, 8),
8866 => conv_std_logic_vector(21, 8),
8867 => conv_std_logic_vector(21, 8),
8868 => conv_std_logic_vector(21, 8),
8869 => conv_std_logic_vector(21, 8),
8870 => conv_std_logic_vector(22, 8),
8871 => conv_std_logic_vector(22, 8),
8872 => conv_std_logic_vector(22, 8),
8873 => conv_std_logic_vector(22, 8),
8874 => conv_std_logic_vector(22, 8),
8875 => conv_std_logic_vector(22, 8),
8876 => conv_std_logic_vector(22, 8),
8877 => conv_std_logic_vector(22, 8),
8878 => conv_std_logic_vector(23, 8),
8879 => conv_std_logic_vector(23, 8),
8880 => conv_std_logic_vector(23, 8),
8881 => conv_std_logic_vector(23, 8),
8882 => conv_std_logic_vector(23, 8),
8883 => conv_std_logic_vector(23, 8),
8884 => conv_std_logic_vector(23, 8),
8885 => conv_std_logic_vector(24, 8),
8886 => conv_std_logic_vector(24, 8),
8887 => conv_std_logic_vector(24, 8),
8888 => conv_std_logic_vector(24, 8),
8889 => conv_std_logic_vector(24, 8),
8890 => conv_std_logic_vector(24, 8),
8891 => conv_std_logic_vector(24, 8),
8892 => conv_std_logic_vector(24, 8),
8893 => conv_std_logic_vector(25, 8),
8894 => conv_std_logic_vector(25, 8),
8895 => conv_std_logic_vector(25, 8),
8896 => conv_std_logic_vector(25, 8),
8897 => conv_std_logic_vector(25, 8),
8898 => conv_std_logic_vector(25, 8),
8899 => conv_std_logic_vector(25, 8),
8900 => conv_std_logic_vector(26, 8),
8901 => conv_std_logic_vector(26, 8),
8902 => conv_std_logic_vector(26, 8),
8903 => conv_std_logic_vector(26, 8),
8904 => conv_std_logic_vector(26, 8),
8905 => conv_std_logic_vector(26, 8),
8906 => conv_std_logic_vector(26, 8),
8907 => conv_std_logic_vector(26, 8),
8908 => conv_std_logic_vector(27, 8),
8909 => conv_std_logic_vector(27, 8),
8910 => conv_std_logic_vector(27, 8),
8911 => conv_std_logic_vector(27, 8),
8912 => conv_std_logic_vector(27, 8),
8913 => conv_std_logic_vector(27, 8),
8914 => conv_std_logic_vector(27, 8),
8915 => conv_std_logic_vector(28, 8),
8916 => conv_std_logic_vector(28, 8),
8917 => conv_std_logic_vector(28, 8),
8918 => conv_std_logic_vector(28, 8),
8919 => conv_std_logic_vector(28, 8),
8920 => conv_std_logic_vector(28, 8),
8921 => conv_std_logic_vector(28, 8),
8922 => conv_std_logic_vector(28, 8),
8923 => conv_std_logic_vector(29, 8),
8924 => conv_std_logic_vector(29, 8),
8925 => conv_std_logic_vector(29, 8),
8926 => conv_std_logic_vector(29, 8),
8927 => conv_std_logic_vector(29, 8),
8928 => conv_std_logic_vector(29, 8),
8929 => conv_std_logic_vector(29, 8),
8930 => conv_std_logic_vector(30, 8),
8931 => conv_std_logic_vector(30, 8),
8932 => conv_std_logic_vector(30, 8),
8933 => conv_std_logic_vector(30, 8),
8934 => conv_std_logic_vector(30, 8),
8935 => conv_std_logic_vector(30, 8),
8936 => conv_std_logic_vector(30, 8),
8937 => conv_std_logic_vector(30, 8),
8938 => conv_std_logic_vector(31, 8),
8939 => conv_std_logic_vector(31, 8),
8940 => conv_std_logic_vector(31, 8),
8941 => conv_std_logic_vector(31, 8),
8942 => conv_std_logic_vector(31, 8),
8943 => conv_std_logic_vector(31, 8),
8944 => conv_std_logic_vector(31, 8),
8945 => conv_std_logic_vector(32, 8),
8946 => conv_std_logic_vector(32, 8),
8947 => conv_std_logic_vector(32, 8),
8948 => conv_std_logic_vector(32, 8),
8949 => conv_std_logic_vector(32, 8),
8950 => conv_std_logic_vector(32, 8),
8951 => conv_std_logic_vector(32, 8),
8952 => conv_std_logic_vector(32, 8),
8953 => conv_std_logic_vector(33, 8),
8954 => conv_std_logic_vector(33, 8),
8955 => conv_std_logic_vector(33, 8),
8956 => conv_std_logic_vector(33, 8),
8957 => conv_std_logic_vector(33, 8),
8958 => conv_std_logic_vector(33, 8),
8959 => conv_std_logic_vector(33, 8),
8960 => conv_std_logic_vector(0, 8),
8961 => conv_std_logic_vector(0, 8),
8962 => conv_std_logic_vector(0, 8),
8963 => conv_std_logic_vector(0, 8),
8964 => conv_std_logic_vector(0, 8),
8965 => conv_std_logic_vector(0, 8),
8966 => conv_std_logic_vector(0, 8),
8967 => conv_std_logic_vector(0, 8),
8968 => conv_std_logic_vector(1, 8),
8969 => conv_std_logic_vector(1, 8),
8970 => conv_std_logic_vector(1, 8),
8971 => conv_std_logic_vector(1, 8),
8972 => conv_std_logic_vector(1, 8),
8973 => conv_std_logic_vector(1, 8),
8974 => conv_std_logic_vector(1, 8),
8975 => conv_std_logic_vector(2, 8),
8976 => conv_std_logic_vector(2, 8),
8977 => conv_std_logic_vector(2, 8),
8978 => conv_std_logic_vector(2, 8),
8979 => conv_std_logic_vector(2, 8),
8980 => conv_std_logic_vector(2, 8),
8981 => conv_std_logic_vector(2, 8),
8982 => conv_std_logic_vector(3, 8),
8983 => conv_std_logic_vector(3, 8),
8984 => conv_std_logic_vector(3, 8),
8985 => conv_std_logic_vector(3, 8),
8986 => conv_std_logic_vector(3, 8),
8987 => conv_std_logic_vector(3, 8),
8988 => conv_std_logic_vector(3, 8),
8989 => conv_std_logic_vector(3, 8),
8990 => conv_std_logic_vector(4, 8),
8991 => conv_std_logic_vector(4, 8),
8992 => conv_std_logic_vector(4, 8),
8993 => conv_std_logic_vector(4, 8),
8994 => conv_std_logic_vector(4, 8),
8995 => conv_std_logic_vector(4, 8),
8996 => conv_std_logic_vector(4, 8),
8997 => conv_std_logic_vector(5, 8),
8998 => conv_std_logic_vector(5, 8),
8999 => conv_std_logic_vector(5, 8),
9000 => conv_std_logic_vector(5, 8),
9001 => conv_std_logic_vector(5, 8),
9002 => conv_std_logic_vector(5, 8),
9003 => conv_std_logic_vector(5, 8),
9004 => conv_std_logic_vector(6, 8),
9005 => conv_std_logic_vector(6, 8),
9006 => conv_std_logic_vector(6, 8),
9007 => conv_std_logic_vector(6, 8),
9008 => conv_std_logic_vector(6, 8),
9009 => conv_std_logic_vector(6, 8),
9010 => conv_std_logic_vector(6, 8),
9011 => conv_std_logic_vector(6, 8),
9012 => conv_std_logic_vector(7, 8),
9013 => conv_std_logic_vector(7, 8),
9014 => conv_std_logic_vector(7, 8),
9015 => conv_std_logic_vector(7, 8),
9016 => conv_std_logic_vector(7, 8),
9017 => conv_std_logic_vector(7, 8),
9018 => conv_std_logic_vector(7, 8),
9019 => conv_std_logic_vector(8, 8),
9020 => conv_std_logic_vector(8, 8),
9021 => conv_std_logic_vector(8, 8),
9022 => conv_std_logic_vector(8, 8),
9023 => conv_std_logic_vector(8, 8),
9024 => conv_std_logic_vector(8, 8),
9025 => conv_std_logic_vector(8, 8),
9026 => conv_std_logic_vector(9, 8),
9027 => conv_std_logic_vector(9, 8),
9028 => conv_std_logic_vector(9, 8),
9029 => conv_std_logic_vector(9, 8),
9030 => conv_std_logic_vector(9, 8),
9031 => conv_std_logic_vector(9, 8),
9032 => conv_std_logic_vector(9, 8),
9033 => conv_std_logic_vector(9, 8),
9034 => conv_std_logic_vector(10, 8),
9035 => conv_std_logic_vector(10, 8),
9036 => conv_std_logic_vector(10, 8),
9037 => conv_std_logic_vector(10, 8),
9038 => conv_std_logic_vector(10, 8),
9039 => conv_std_logic_vector(10, 8),
9040 => conv_std_logic_vector(10, 8),
9041 => conv_std_logic_vector(11, 8),
9042 => conv_std_logic_vector(11, 8),
9043 => conv_std_logic_vector(11, 8),
9044 => conv_std_logic_vector(11, 8),
9045 => conv_std_logic_vector(11, 8),
9046 => conv_std_logic_vector(11, 8),
9047 => conv_std_logic_vector(11, 8),
9048 => conv_std_logic_vector(12, 8),
9049 => conv_std_logic_vector(12, 8),
9050 => conv_std_logic_vector(12, 8),
9051 => conv_std_logic_vector(12, 8),
9052 => conv_std_logic_vector(12, 8),
9053 => conv_std_logic_vector(12, 8),
9054 => conv_std_logic_vector(12, 8),
9055 => conv_std_logic_vector(12, 8),
9056 => conv_std_logic_vector(13, 8),
9057 => conv_std_logic_vector(13, 8),
9058 => conv_std_logic_vector(13, 8),
9059 => conv_std_logic_vector(13, 8),
9060 => conv_std_logic_vector(13, 8),
9061 => conv_std_logic_vector(13, 8),
9062 => conv_std_logic_vector(13, 8),
9063 => conv_std_logic_vector(14, 8),
9064 => conv_std_logic_vector(14, 8),
9065 => conv_std_logic_vector(14, 8),
9066 => conv_std_logic_vector(14, 8),
9067 => conv_std_logic_vector(14, 8),
9068 => conv_std_logic_vector(14, 8),
9069 => conv_std_logic_vector(14, 8),
9070 => conv_std_logic_vector(15, 8),
9071 => conv_std_logic_vector(15, 8),
9072 => conv_std_logic_vector(15, 8),
9073 => conv_std_logic_vector(15, 8),
9074 => conv_std_logic_vector(15, 8),
9075 => conv_std_logic_vector(15, 8),
9076 => conv_std_logic_vector(15, 8),
9077 => conv_std_logic_vector(15, 8),
9078 => conv_std_logic_vector(16, 8),
9079 => conv_std_logic_vector(16, 8),
9080 => conv_std_logic_vector(16, 8),
9081 => conv_std_logic_vector(16, 8),
9082 => conv_std_logic_vector(16, 8),
9083 => conv_std_logic_vector(16, 8),
9084 => conv_std_logic_vector(16, 8),
9085 => conv_std_logic_vector(17, 8),
9086 => conv_std_logic_vector(17, 8),
9087 => conv_std_logic_vector(17, 8),
9088 => conv_std_logic_vector(17, 8),
9089 => conv_std_logic_vector(17, 8),
9090 => conv_std_logic_vector(17, 8),
9091 => conv_std_logic_vector(17, 8),
9092 => conv_std_logic_vector(18, 8),
9093 => conv_std_logic_vector(18, 8),
9094 => conv_std_logic_vector(18, 8),
9095 => conv_std_logic_vector(18, 8),
9096 => conv_std_logic_vector(18, 8),
9097 => conv_std_logic_vector(18, 8),
9098 => conv_std_logic_vector(18, 8),
9099 => conv_std_logic_vector(19, 8),
9100 => conv_std_logic_vector(19, 8),
9101 => conv_std_logic_vector(19, 8),
9102 => conv_std_logic_vector(19, 8),
9103 => conv_std_logic_vector(19, 8),
9104 => conv_std_logic_vector(19, 8),
9105 => conv_std_logic_vector(19, 8),
9106 => conv_std_logic_vector(19, 8),
9107 => conv_std_logic_vector(20, 8),
9108 => conv_std_logic_vector(20, 8),
9109 => conv_std_logic_vector(20, 8),
9110 => conv_std_logic_vector(20, 8),
9111 => conv_std_logic_vector(20, 8),
9112 => conv_std_logic_vector(20, 8),
9113 => conv_std_logic_vector(20, 8),
9114 => conv_std_logic_vector(21, 8),
9115 => conv_std_logic_vector(21, 8),
9116 => conv_std_logic_vector(21, 8),
9117 => conv_std_logic_vector(21, 8),
9118 => conv_std_logic_vector(21, 8),
9119 => conv_std_logic_vector(21, 8),
9120 => conv_std_logic_vector(21, 8),
9121 => conv_std_logic_vector(22, 8),
9122 => conv_std_logic_vector(22, 8),
9123 => conv_std_logic_vector(22, 8),
9124 => conv_std_logic_vector(22, 8),
9125 => conv_std_logic_vector(22, 8),
9126 => conv_std_logic_vector(22, 8),
9127 => conv_std_logic_vector(22, 8),
9128 => conv_std_logic_vector(22, 8),
9129 => conv_std_logic_vector(23, 8),
9130 => conv_std_logic_vector(23, 8),
9131 => conv_std_logic_vector(23, 8),
9132 => conv_std_logic_vector(23, 8),
9133 => conv_std_logic_vector(23, 8),
9134 => conv_std_logic_vector(23, 8),
9135 => conv_std_logic_vector(23, 8),
9136 => conv_std_logic_vector(24, 8),
9137 => conv_std_logic_vector(24, 8),
9138 => conv_std_logic_vector(24, 8),
9139 => conv_std_logic_vector(24, 8),
9140 => conv_std_logic_vector(24, 8),
9141 => conv_std_logic_vector(24, 8),
9142 => conv_std_logic_vector(24, 8),
9143 => conv_std_logic_vector(25, 8),
9144 => conv_std_logic_vector(25, 8),
9145 => conv_std_logic_vector(25, 8),
9146 => conv_std_logic_vector(25, 8),
9147 => conv_std_logic_vector(25, 8),
9148 => conv_std_logic_vector(25, 8),
9149 => conv_std_logic_vector(25, 8),
9150 => conv_std_logic_vector(25, 8),
9151 => conv_std_logic_vector(26, 8),
9152 => conv_std_logic_vector(26, 8),
9153 => conv_std_logic_vector(26, 8),
9154 => conv_std_logic_vector(26, 8),
9155 => conv_std_logic_vector(26, 8),
9156 => conv_std_logic_vector(26, 8),
9157 => conv_std_logic_vector(26, 8),
9158 => conv_std_logic_vector(27, 8),
9159 => conv_std_logic_vector(27, 8),
9160 => conv_std_logic_vector(27, 8),
9161 => conv_std_logic_vector(27, 8),
9162 => conv_std_logic_vector(27, 8),
9163 => conv_std_logic_vector(27, 8),
9164 => conv_std_logic_vector(27, 8),
9165 => conv_std_logic_vector(28, 8),
9166 => conv_std_logic_vector(28, 8),
9167 => conv_std_logic_vector(28, 8),
9168 => conv_std_logic_vector(28, 8),
9169 => conv_std_logic_vector(28, 8),
9170 => conv_std_logic_vector(28, 8),
9171 => conv_std_logic_vector(28, 8),
9172 => conv_std_logic_vector(28, 8),
9173 => conv_std_logic_vector(29, 8),
9174 => conv_std_logic_vector(29, 8),
9175 => conv_std_logic_vector(29, 8),
9176 => conv_std_logic_vector(29, 8),
9177 => conv_std_logic_vector(29, 8),
9178 => conv_std_logic_vector(29, 8),
9179 => conv_std_logic_vector(29, 8),
9180 => conv_std_logic_vector(30, 8),
9181 => conv_std_logic_vector(30, 8),
9182 => conv_std_logic_vector(30, 8),
9183 => conv_std_logic_vector(30, 8),
9184 => conv_std_logic_vector(30, 8),
9185 => conv_std_logic_vector(30, 8),
9186 => conv_std_logic_vector(30, 8),
9187 => conv_std_logic_vector(31, 8),
9188 => conv_std_logic_vector(31, 8),
9189 => conv_std_logic_vector(31, 8),
9190 => conv_std_logic_vector(31, 8),
9191 => conv_std_logic_vector(31, 8),
9192 => conv_std_logic_vector(31, 8),
9193 => conv_std_logic_vector(31, 8),
9194 => conv_std_logic_vector(31, 8),
9195 => conv_std_logic_vector(32, 8),
9196 => conv_std_logic_vector(32, 8),
9197 => conv_std_logic_vector(32, 8),
9198 => conv_std_logic_vector(32, 8),
9199 => conv_std_logic_vector(32, 8),
9200 => conv_std_logic_vector(32, 8),
9201 => conv_std_logic_vector(32, 8),
9202 => conv_std_logic_vector(33, 8),
9203 => conv_std_logic_vector(33, 8),
9204 => conv_std_logic_vector(33, 8),
9205 => conv_std_logic_vector(33, 8),
9206 => conv_std_logic_vector(33, 8),
9207 => conv_std_logic_vector(33, 8),
9208 => conv_std_logic_vector(33, 8),
9209 => conv_std_logic_vector(34, 8),
9210 => conv_std_logic_vector(34, 8),
9211 => conv_std_logic_vector(34, 8),
9212 => conv_std_logic_vector(34, 8),
9213 => conv_std_logic_vector(34, 8),
9214 => conv_std_logic_vector(34, 8),
9215 => conv_std_logic_vector(34, 8),
9216 => conv_std_logic_vector(0, 8),
9217 => conv_std_logic_vector(0, 8),
9218 => conv_std_logic_vector(0, 8),
9219 => conv_std_logic_vector(0, 8),
9220 => conv_std_logic_vector(0, 8),
9221 => conv_std_logic_vector(0, 8),
9222 => conv_std_logic_vector(0, 8),
9223 => conv_std_logic_vector(0, 8),
9224 => conv_std_logic_vector(1, 8),
9225 => conv_std_logic_vector(1, 8),
9226 => conv_std_logic_vector(1, 8),
9227 => conv_std_logic_vector(1, 8),
9228 => conv_std_logic_vector(1, 8),
9229 => conv_std_logic_vector(1, 8),
9230 => conv_std_logic_vector(1, 8),
9231 => conv_std_logic_vector(2, 8),
9232 => conv_std_logic_vector(2, 8),
9233 => conv_std_logic_vector(2, 8),
9234 => conv_std_logic_vector(2, 8),
9235 => conv_std_logic_vector(2, 8),
9236 => conv_std_logic_vector(2, 8),
9237 => conv_std_logic_vector(2, 8),
9238 => conv_std_logic_vector(3, 8),
9239 => conv_std_logic_vector(3, 8),
9240 => conv_std_logic_vector(3, 8),
9241 => conv_std_logic_vector(3, 8),
9242 => conv_std_logic_vector(3, 8),
9243 => conv_std_logic_vector(3, 8),
9244 => conv_std_logic_vector(3, 8),
9245 => conv_std_logic_vector(4, 8),
9246 => conv_std_logic_vector(4, 8),
9247 => conv_std_logic_vector(4, 8),
9248 => conv_std_logic_vector(4, 8),
9249 => conv_std_logic_vector(4, 8),
9250 => conv_std_logic_vector(4, 8),
9251 => conv_std_logic_vector(4, 8),
9252 => conv_std_logic_vector(5, 8),
9253 => conv_std_logic_vector(5, 8),
9254 => conv_std_logic_vector(5, 8),
9255 => conv_std_logic_vector(5, 8),
9256 => conv_std_logic_vector(5, 8),
9257 => conv_std_logic_vector(5, 8),
9258 => conv_std_logic_vector(5, 8),
9259 => conv_std_logic_vector(6, 8),
9260 => conv_std_logic_vector(6, 8),
9261 => conv_std_logic_vector(6, 8),
9262 => conv_std_logic_vector(6, 8),
9263 => conv_std_logic_vector(6, 8),
9264 => conv_std_logic_vector(6, 8),
9265 => conv_std_logic_vector(6, 8),
9266 => conv_std_logic_vector(7, 8),
9267 => conv_std_logic_vector(7, 8),
9268 => conv_std_logic_vector(7, 8),
9269 => conv_std_logic_vector(7, 8),
9270 => conv_std_logic_vector(7, 8),
9271 => conv_std_logic_vector(7, 8),
9272 => conv_std_logic_vector(7, 8),
9273 => conv_std_logic_vector(8, 8),
9274 => conv_std_logic_vector(8, 8),
9275 => conv_std_logic_vector(8, 8),
9276 => conv_std_logic_vector(8, 8),
9277 => conv_std_logic_vector(8, 8),
9278 => conv_std_logic_vector(8, 8),
9279 => conv_std_logic_vector(8, 8),
9280 => conv_std_logic_vector(9, 8),
9281 => conv_std_logic_vector(9, 8),
9282 => conv_std_logic_vector(9, 8),
9283 => conv_std_logic_vector(9, 8),
9284 => conv_std_logic_vector(9, 8),
9285 => conv_std_logic_vector(9, 8),
9286 => conv_std_logic_vector(9, 8),
9287 => conv_std_logic_vector(9, 8),
9288 => conv_std_logic_vector(10, 8),
9289 => conv_std_logic_vector(10, 8),
9290 => conv_std_logic_vector(10, 8),
9291 => conv_std_logic_vector(10, 8),
9292 => conv_std_logic_vector(10, 8),
9293 => conv_std_logic_vector(10, 8),
9294 => conv_std_logic_vector(10, 8),
9295 => conv_std_logic_vector(11, 8),
9296 => conv_std_logic_vector(11, 8),
9297 => conv_std_logic_vector(11, 8),
9298 => conv_std_logic_vector(11, 8),
9299 => conv_std_logic_vector(11, 8),
9300 => conv_std_logic_vector(11, 8),
9301 => conv_std_logic_vector(11, 8),
9302 => conv_std_logic_vector(12, 8),
9303 => conv_std_logic_vector(12, 8),
9304 => conv_std_logic_vector(12, 8),
9305 => conv_std_logic_vector(12, 8),
9306 => conv_std_logic_vector(12, 8),
9307 => conv_std_logic_vector(12, 8),
9308 => conv_std_logic_vector(12, 8),
9309 => conv_std_logic_vector(13, 8),
9310 => conv_std_logic_vector(13, 8),
9311 => conv_std_logic_vector(13, 8),
9312 => conv_std_logic_vector(13, 8),
9313 => conv_std_logic_vector(13, 8),
9314 => conv_std_logic_vector(13, 8),
9315 => conv_std_logic_vector(13, 8),
9316 => conv_std_logic_vector(14, 8),
9317 => conv_std_logic_vector(14, 8),
9318 => conv_std_logic_vector(14, 8),
9319 => conv_std_logic_vector(14, 8),
9320 => conv_std_logic_vector(14, 8),
9321 => conv_std_logic_vector(14, 8),
9322 => conv_std_logic_vector(14, 8),
9323 => conv_std_logic_vector(15, 8),
9324 => conv_std_logic_vector(15, 8),
9325 => conv_std_logic_vector(15, 8),
9326 => conv_std_logic_vector(15, 8),
9327 => conv_std_logic_vector(15, 8),
9328 => conv_std_logic_vector(15, 8),
9329 => conv_std_logic_vector(15, 8),
9330 => conv_std_logic_vector(16, 8),
9331 => conv_std_logic_vector(16, 8),
9332 => conv_std_logic_vector(16, 8),
9333 => conv_std_logic_vector(16, 8),
9334 => conv_std_logic_vector(16, 8),
9335 => conv_std_logic_vector(16, 8),
9336 => conv_std_logic_vector(16, 8),
9337 => conv_std_logic_vector(17, 8),
9338 => conv_std_logic_vector(17, 8),
9339 => conv_std_logic_vector(17, 8),
9340 => conv_std_logic_vector(17, 8),
9341 => conv_std_logic_vector(17, 8),
9342 => conv_std_logic_vector(17, 8),
9343 => conv_std_logic_vector(17, 8),
9344 => conv_std_logic_vector(18, 8),
9345 => conv_std_logic_vector(18, 8),
9346 => conv_std_logic_vector(18, 8),
9347 => conv_std_logic_vector(18, 8),
9348 => conv_std_logic_vector(18, 8),
9349 => conv_std_logic_vector(18, 8),
9350 => conv_std_logic_vector(18, 8),
9351 => conv_std_logic_vector(18, 8),
9352 => conv_std_logic_vector(19, 8),
9353 => conv_std_logic_vector(19, 8),
9354 => conv_std_logic_vector(19, 8),
9355 => conv_std_logic_vector(19, 8),
9356 => conv_std_logic_vector(19, 8),
9357 => conv_std_logic_vector(19, 8),
9358 => conv_std_logic_vector(19, 8),
9359 => conv_std_logic_vector(20, 8),
9360 => conv_std_logic_vector(20, 8),
9361 => conv_std_logic_vector(20, 8),
9362 => conv_std_logic_vector(20, 8),
9363 => conv_std_logic_vector(20, 8),
9364 => conv_std_logic_vector(20, 8),
9365 => conv_std_logic_vector(20, 8),
9366 => conv_std_logic_vector(21, 8),
9367 => conv_std_logic_vector(21, 8),
9368 => conv_std_logic_vector(21, 8),
9369 => conv_std_logic_vector(21, 8),
9370 => conv_std_logic_vector(21, 8),
9371 => conv_std_logic_vector(21, 8),
9372 => conv_std_logic_vector(21, 8),
9373 => conv_std_logic_vector(22, 8),
9374 => conv_std_logic_vector(22, 8),
9375 => conv_std_logic_vector(22, 8),
9376 => conv_std_logic_vector(22, 8),
9377 => conv_std_logic_vector(22, 8),
9378 => conv_std_logic_vector(22, 8),
9379 => conv_std_logic_vector(22, 8),
9380 => conv_std_logic_vector(23, 8),
9381 => conv_std_logic_vector(23, 8),
9382 => conv_std_logic_vector(23, 8),
9383 => conv_std_logic_vector(23, 8),
9384 => conv_std_logic_vector(23, 8),
9385 => conv_std_logic_vector(23, 8),
9386 => conv_std_logic_vector(23, 8),
9387 => conv_std_logic_vector(24, 8),
9388 => conv_std_logic_vector(24, 8),
9389 => conv_std_logic_vector(24, 8),
9390 => conv_std_logic_vector(24, 8),
9391 => conv_std_logic_vector(24, 8),
9392 => conv_std_logic_vector(24, 8),
9393 => conv_std_logic_vector(24, 8),
9394 => conv_std_logic_vector(25, 8),
9395 => conv_std_logic_vector(25, 8),
9396 => conv_std_logic_vector(25, 8),
9397 => conv_std_logic_vector(25, 8),
9398 => conv_std_logic_vector(25, 8),
9399 => conv_std_logic_vector(25, 8),
9400 => conv_std_logic_vector(25, 8),
9401 => conv_std_logic_vector(26, 8),
9402 => conv_std_logic_vector(26, 8),
9403 => conv_std_logic_vector(26, 8),
9404 => conv_std_logic_vector(26, 8),
9405 => conv_std_logic_vector(26, 8),
9406 => conv_std_logic_vector(26, 8),
9407 => conv_std_logic_vector(26, 8),
9408 => conv_std_logic_vector(27, 8),
9409 => conv_std_logic_vector(27, 8),
9410 => conv_std_logic_vector(27, 8),
9411 => conv_std_logic_vector(27, 8),
9412 => conv_std_logic_vector(27, 8),
9413 => conv_std_logic_vector(27, 8),
9414 => conv_std_logic_vector(27, 8),
9415 => conv_std_logic_vector(27, 8),
9416 => conv_std_logic_vector(28, 8),
9417 => conv_std_logic_vector(28, 8),
9418 => conv_std_logic_vector(28, 8),
9419 => conv_std_logic_vector(28, 8),
9420 => conv_std_logic_vector(28, 8),
9421 => conv_std_logic_vector(28, 8),
9422 => conv_std_logic_vector(28, 8),
9423 => conv_std_logic_vector(29, 8),
9424 => conv_std_logic_vector(29, 8),
9425 => conv_std_logic_vector(29, 8),
9426 => conv_std_logic_vector(29, 8),
9427 => conv_std_logic_vector(29, 8),
9428 => conv_std_logic_vector(29, 8),
9429 => conv_std_logic_vector(29, 8),
9430 => conv_std_logic_vector(30, 8),
9431 => conv_std_logic_vector(30, 8),
9432 => conv_std_logic_vector(30, 8),
9433 => conv_std_logic_vector(30, 8),
9434 => conv_std_logic_vector(30, 8),
9435 => conv_std_logic_vector(30, 8),
9436 => conv_std_logic_vector(30, 8),
9437 => conv_std_logic_vector(31, 8),
9438 => conv_std_logic_vector(31, 8),
9439 => conv_std_logic_vector(31, 8),
9440 => conv_std_logic_vector(31, 8),
9441 => conv_std_logic_vector(31, 8),
9442 => conv_std_logic_vector(31, 8),
9443 => conv_std_logic_vector(31, 8),
9444 => conv_std_logic_vector(32, 8),
9445 => conv_std_logic_vector(32, 8),
9446 => conv_std_logic_vector(32, 8),
9447 => conv_std_logic_vector(32, 8),
9448 => conv_std_logic_vector(32, 8),
9449 => conv_std_logic_vector(32, 8),
9450 => conv_std_logic_vector(32, 8),
9451 => conv_std_logic_vector(33, 8),
9452 => conv_std_logic_vector(33, 8),
9453 => conv_std_logic_vector(33, 8),
9454 => conv_std_logic_vector(33, 8),
9455 => conv_std_logic_vector(33, 8),
9456 => conv_std_logic_vector(33, 8),
9457 => conv_std_logic_vector(33, 8),
9458 => conv_std_logic_vector(34, 8),
9459 => conv_std_logic_vector(34, 8),
9460 => conv_std_logic_vector(34, 8),
9461 => conv_std_logic_vector(34, 8),
9462 => conv_std_logic_vector(34, 8),
9463 => conv_std_logic_vector(34, 8),
9464 => conv_std_logic_vector(34, 8),
9465 => conv_std_logic_vector(35, 8),
9466 => conv_std_logic_vector(35, 8),
9467 => conv_std_logic_vector(35, 8),
9468 => conv_std_logic_vector(35, 8),
9469 => conv_std_logic_vector(35, 8),
9470 => conv_std_logic_vector(35, 8),
9471 => conv_std_logic_vector(35, 8),
9472 => conv_std_logic_vector(0, 8),
9473 => conv_std_logic_vector(0, 8),
9474 => conv_std_logic_vector(0, 8),
9475 => conv_std_logic_vector(0, 8),
9476 => conv_std_logic_vector(0, 8),
9477 => conv_std_logic_vector(0, 8),
9478 => conv_std_logic_vector(0, 8),
9479 => conv_std_logic_vector(1, 8),
9480 => conv_std_logic_vector(1, 8),
9481 => conv_std_logic_vector(1, 8),
9482 => conv_std_logic_vector(1, 8),
9483 => conv_std_logic_vector(1, 8),
9484 => conv_std_logic_vector(1, 8),
9485 => conv_std_logic_vector(1, 8),
9486 => conv_std_logic_vector(2, 8),
9487 => conv_std_logic_vector(2, 8),
9488 => conv_std_logic_vector(2, 8),
9489 => conv_std_logic_vector(2, 8),
9490 => conv_std_logic_vector(2, 8),
9491 => conv_std_logic_vector(2, 8),
9492 => conv_std_logic_vector(2, 8),
9493 => conv_std_logic_vector(3, 8),
9494 => conv_std_logic_vector(3, 8),
9495 => conv_std_logic_vector(3, 8),
9496 => conv_std_logic_vector(3, 8),
9497 => conv_std_logic_vector(3, 8),
9498 => conv_std_logic_vector(3, 8),
9499 => conv_std_logic_vector(3, 8),
9500 => conv_std_logic_vector(4, 8),
9501 => conv_std_logic_vector(4, 8),
9502 => conv_std_logic_vector(4, 8),
9503 => conv_std_logic_vector(4, 8),
9504 => conv_std_logic_vector(4, 8),
9505 => conv_std_logic_vector(4, 8),
9506 => conv_std_logic_vector(4, 8),
9507 => conv_std_logic_vector(5, 8),
9508 => conv_std_logic_vector(5, 8),
9509 => conv_std_logic_vector(5, 8),
9510 => conv_std_logic_vector(5, 8),
9511 => conv_std_logic_vector(5, 8),
9512 => conv_std_logic_vector(5, 8),
9513 => conv_std_logic_vector(5, 8),
9514 => conv_std_logic_vector(6, 8),
9515 => conv_std_logic_vector(6, 8),
9516 => conv_std_logic_vector(6, 8),
9517 => conv_std_logic_vector(6, 8),
9518 => conv_std_logic_vector(6, 8),
9519 => conv_std_logic_vector(6, 8),
9520 => conv_std_logic_vector(6, 8),
9521 => conv_std_logic_vector(7, 8),
9522 => conv_std_logic_vector(7, 8),
9523 => conv_std_logic_vector(7, 8),
9524 => conv_std_logic_vector(7, 8),
9525 => conv_std_logic_vector(7, 8),
9526 => conv_std_logic_vector(7, 8),
9527 => conv_std_logic_vector(7, 8),
9528 => conv_std_logic_vector(8, 8),
9529 => conv_std_logic_vector(8, 8),
9530 => conv_std_logic_vector(8, 8),
9531 => conv_std_logic_vector(8, 8),
9532 => conv_std_logic_vector(8, 8),
9533 => conv_std_logic_vector(8, 8),
9534 => conv_std_logic_vector(8, 8),
9535 => conv_std_logic_vector(9, 8),
9536 => conv_std_logic_vector(9, 8),
9537 => conv_std_logic_vector(9, 8),
9538 => conv_std_logic_vector(9, 8),
9539 => conv_std_logic_vector(9, 8),
9540 => conv_std_logic_vector(9, 8),
9541 => conv_std_logic_vector(9, 8),
9542 => conv_std_logic_vector(10, 8),
9543 => conv_std_logic_vector(10, 8),
9544 => conv_std_logic_vector(10, 8),
9545 => conv_std_logic_vector(10, 8),
9546 => conv_std_logic_vector(10, 8),
9547 => conv_std_logic_vector(10, 8),
9548 => conv_std_logic_vector(10, 8),
9549 => conv_std_logic_vector(11, 8),
9550 => conv_std_logic_vector(11, 8),
9551 => conv_std_logic_vector(11, 8),
9552 => conv_std_logic_vector(11, 8),
9553 => conv_std_logic_vector(11, 8),
9554 => conv_std_logic_vector(11, 8),
9555 => conv_std_logic_vector(11, 8),
9556 => conv_std_logic_vector(12, 8),
9557 => conv_std_logic_vector(12, 8),
9558 => conv_std_logic_vector(12, 8),
9559 => conv_std_logic_vector(12, 8),
9560 => conv_std_logic_vector(12, 8),
9561 => conv_std_logic_vector(12, 8),
9562 => conv_std_logic_vector(13, 8),
9563 => conv_std_logic_vector(13, 8),
9564 => conv_std_logic_vector(13, 8),
9565 => conv_std_logic_vector(13, 8),
9566 => conv_std_logic_vector(13, 8),
9567 => conv_std_logic_vector(13, 8),
9568 => conv_std_logic_vector(13, 8),
9569 => conv_std_logic_vector(14, 8),
9570 => conv_std_logic_vector(14, 8),
9571 => conv_std_logic_vector(14, 8),
9572 => conv_std_logic_vector(14, 8),
9573 => conv_std_logic_vector(14, 8),
9574 => conv_std_logic_vector(14, 8),
9575 => conv_std_logic_vector(14, 8),
9576 => conv_std_logic_vector(15, 8),
9577 => conv_std_logic_vector(15, 8),
9578 => conv_std_logic_vector(15, 8),
9579 => conv_std_logic_vector(15, 8),
9580 => conv_std_logic_vector(15, 8),
9581 => conv_std_logic_vector(15, 8),
9582 => conv_std_logic_vector(15, 8),
9583 => conv_std_logic_vector(16, 8),
9584 => conv_std_logic_vector(16, 8),
9585 => conv_std_logic_vector(16, 8),
9586 => conv_std_logic_vector(16, 8),
9587 => conv_std_logic_vector(16, 8),
9588 => conv_std_logic_vector(16, 8),
9589 => conv_std_logic_vector(16, 8),
9590 => conv_std_logic_vector(17, 8),
9591 => conv_std_logic_vector(17, 8),
9592 => conv_std_logic_vector(17, 8),
9593 => conv_std_logic_vector(17, 8),
9594 => conv_std_logic_vector(17, 8),
9595 => conv_std_logic_vector(17, 8),
9596 => conv_std_logic_vector(17, 8),
9597 => conv_std_logic_vector(18, 8),
9598 => conv_std_logic_vector(18, 8),
9599 => conv_std_logic_vector(18, 8),
9600 => conv_std_logic_vector(18, 8),
9601 => conv_std_logic_vector(18, 8),
9602 => conv_std_logic_vector(18, 8),
9603 => conv_std_logic_vector(18, 8),
9604 => conv_std_logic_vector(19, 8),
9605 => conv_std_logic_vector(19, 8),
9606 => conv_std_logic_vector(19, 8),
9607 => conv_std_logic_vector(19, 8),
9608 => conv_std_logic_vector(19, 8),
9609 => conv_std_logic_vector(19, 8),
9610 => conv_std_logic_vector(19, 8),
9611 => conv_std_logic_vector(20, 8),
9612 => conv_std_logic_vector(20, 8),
9613 => conv_std_logic_vector(20, 8),
9614 => conv_std_logic_vector(20, 8),
9615 => conv_std_logic_vector(20, 8),
9616 => conv_std_logic_vector(20, 8),
9617 => conv_std_logic_vector(20, 8),
9618 => conv_std_logic_vector(21, 8),
9619 => conv_std_logic_vector(21, 8),
9620 => conv_std_logic_vector(21, 8),
9621 => conv_std_logic_vector(21, 8),
9622 => conv_std_logic_vector(21, 8),
9623 => conv_std_logic_vector(21, 8),
9624 => conv_std_logic_vector(21, 8),
9625 => conv_std_logic_vector(22, 8),
9626 => conv_std_logic_vector(22, 8),
9627 => conv_std_logic_vector(22, 8),
9628 => conv_std_logic_vector(22, 8),
9629 => conv_std_logic_vector(22, 8),
9630 => conv_std_logic_vector(22, 8),
9631 => conv_std_logic_vector(22, 8),
9632 => conv_std_logic_vector(23, 8),
9633 => conv_std_logic_vector(23, 8),
9634 => conv_std_logic_vector(23, 8),
9635 => conv_std_logic_vector(23, 8),
9636 => conv_std_logic_vector(23, 8),
9637 => conv_std_logic_vector(23, 8),
9638 => conv_std_logic_vector(23, 8),
9639 => conv_std_logic_vector(24, 8),
9640 => conv_std_logic_vector(24, 8),
9641 => conv_std_logic_vector(24, 8),
9642 => conv_std_logic_vector(24, 8),
9643 => conv_std_logic_vector(24, 8),
9644 => conv_std_logic_vector(24, 8),
9645 => conv_std_logic_vector(25, 8),
9646 => conv_std_logic_vector(25, 8),
9647 => conv_std_logic_vector(25, 8),
9648 => conv_std_logic_vector(25, 8),
9649 => conv_std_logic_vector(25, 8),
9650 => conv_std_logic_vector(25, 8),
9651 => conv_std_logic_vector(25, 8),
9652 => conv_std_logic_vector(26, 8),
9653 => conv_std_logic_vector(26, 8),
9654 => conv_std_logic_vector(26, 8),
9655 => conv_std_logic_vector(26, 8),
9656 => conv_std_logic_vector(26, 8),
9657 => conv_std_logic_vector(26, 8),
9658 => conv_std_logic_vector(26, 8),
9659 => conv_std_logic_vector(27, 8),
9660 => conv_std_logic_vector(27, 8),
9661 => conv_std_logic_vector(27, 8),
9662 => conv_std_logic_vector(27, 8),
9663 => conv_std_logic_vector(27, 8),
9664 => conv_std_logic_vector(27, 8),
9665 => conv_std_logic_vector(27, 8),
9666 => conv_std_logic_vector(28, 8),
9667 => conv_std_logic_vector(28, 8),
9668 => conv_std_logic_vector(28, 8),
9669 => conv_std_logic_vector(28, 8),
9670 => conv_std_logic_vector(28, 8),
9671 => conv_std_logic_vector(28, 8),
9672 => conv_std_logic_vector(28, 8),
9673 => conv_std_logic_vector(29, 8),
9674 => conv_std_logic_vector(29, 8),
9675 => conv_std_logic_vector(29, 8),
9676 => conv_std_logic_vector(29, 8),
9677 => conv_std_logic_vector(29, 8),
9678 => conv_std_logic_vector(29, 8),
9679 => conv_std_logic_vector(29, 8),
9680 => conv_std_logic_vector(30, 8),
9681 => conv_std_logic_vector(30, 8),
9682 => conv_std_logic_vector(30, 8),
9683 => conv_std_logic_vector(30, 8),
9684 => conv_std_logic_vector(30, 8),
9685 => conv_std_logic_vector(30, 8),
9686 => conv_std_logic_vector(30, 8),
9687 => conv_std_logic_vector(31, 8),
9688 => conv_std_logic_vector(31, 8),
9689 => conv_std_logic_vector(31, 8),
9690 => conv_std_logic_vector(31, 8),
9691 => conv_std_logic_vector(31, 8),
9692 => conv_std_logic_vector(31, 8),
9693 => conv_std_logic_vector(31, 8),
9694 => conv_std_logic_vector(32, 8),
9695 => conv_std_logic_vector(32, 8),
9696 => conv_std_logic_vector(32, 8),
9697 => conv_std_logic_vector(32, 8),
9698 => conv_std_logic_vector(32, 8),
9699 => conv_std_logic_vector(32, 8),
9700 => conv_std_logic_vector(32, 8),
9701 => conv_std_logic_vector(33, 8),
9702 => conv_std_logic_vector(33, 8),
9703 => conv_std_logic_vector(33, 8),
9704 => conv_std_logic_vector(33, 8),
9705 => conv_std_logic_vector(33, 8),
9706 => conv_std_logic_vector(33, 8),
9707 => conv_std_logic_vector(33, 8),
9708 => conv_std_logic_vector(34, 8),
9709 => conv_std_logic_vector(34, 8),
9710 => conv_std_logic_vector(34, 8),
9711 => conv_std_logic_vector(34, 8),
9712 => conv_std_logic_vector(34, 8),
9713 => conv_std_logic_vector(34, 8),
9714 => conv_std_logic_vector(34, 8),
9715 => conv_std_logic_vector(35, 8),
9716 => conv_std_logic_vector(35, 8),
9717 => conv_std_logic_vector(35, 8),
9718 => conv_std_logic_vector(35, 8),
9719 => conv_std_logic_vector(35, 8),
9720 => conv_std_logic_vector(35, 8),
9721 => conv_std_logic_vector(35, 8),
9722 => conv_std_logic_vector(36, 8),
9723 => conv_std_logic_vector(36, 8),
9724 => conv_std_logic_vector(36, 8),
9725 => conv_std_logic_vector(36, 8),
9726 => conv_std_logic_vector(36, 8),
9727 => conv_std_logic_vector(36, 8),
9728 => conv_std_logic_vector(0, 8),
9729 => conv_std_logic_vector(0, 8),
9730 => conv_std_logic_vector(0, 8),
9731 => conv_std_logic_vector(0, 8),
9732 => conv_std_logic_vector(0, 8),
9733 => conv_std_logic_vector(0, 8),
9734 => conv_std_logic_vector(0, 8),
9735 => conv_std_logic_vector(1, 8),
9736 => conv_std_logic_vector(1, 8),
9737 => conv_std_logic_vector(1, 8),
9738 => conv_std_logic_vector(1, 8),
9739 => conv_std_logic_vector(1, 8),
9740 => conv_std_logic_vector(1, 8),
9741 => conv_std_logic_vector(1, 8),
9742 => conv_std_logic_vector(2, 8),
9743 => conv_std_logic_vector(2, 8),
9744 => conv_std_logic_vector(2, 8),
9745 => conv_std_logic_vector(2, 8),
9746 => conv_std_logic_vector(2, 8),
9747 => conv_std_logic_vector(2, 8),
9748 => conv_std_logic_vector(2, 8),
9749 => conv_std_logic_vector(3, 8),
9750 => conv_std_logic_vector(3, 8),
9751 => conv_std_logic_vector(3, 8),
9752 => conv_std_logic_vector(3, 8),
9753 => conv_std_logic_vector(3, 8),
9754 => conv_std_logic_vector(3, 8),
9755 => conv_std_logic_vector(4, 8),
9756 => conv_std_logic_vector(4, 8),
9757 => conv_std_logic_vector(4, 8),
9758 => conv_std_logic_vector(4, 8),
9759 => conv_std_logic_vector(4, 8),
9760 => conv_std_logic_vector(4, 8),
9761 => conv_std_logic_vector(4, 8),
9762 => conv_std_logic_vector(5, 8),
9763 => conv_std_logic_vector(5, 8),
9764 => conv_std_logic_vector(5, 8),
9765 => conv_std_logic_vector(5, 8),
9766 => conv_std_logic_vector(5, 8),
9767 => conv_std_logic_vector(5, 8),
9768 => conv_std_logic_vector(5, 8),
9769 => conv_std_logic_vector(6, 8),
9770 => conv_std_logic_vector(6, 8),
9771 => conv_std_logic_vector(6, 8),
9772 => conv_std_logic_vector(6, 8),
9773 => conv_std_logic_vector(6, 8),
9774 => conv_std_logic_vector(6, 8),
9775 => conv_std_logic_vector(6, 8),
9776 => conv_std_logic_vector(7, 8),
9777 => conv_std_logic_vector(7, 8),
9778 => conv_std_logic_vector(7, 8),
9779 => conv_std_logic_vector(7, 8),
9780 => conv_std_logic_vector(7, 8),
9781 => conv_std_logic_vector(7, 8),
9782 => conv_std_logic_vector(8, 8),
9783 => conv_std_logic_vector(8, 8),
9784 => conv_std_logic_vector(8, 8),
9785 => conv_std_logic_vector(8, 8),
9786 => conv_std_logic_vector(8, 8),
9787 => conv_std_logic_vector(8, 8),
9788 => conv_std_logic_vector(8, 8),
9789 => conv_std_logic_vector(9, 8),
9790 => conv_std_logic_vector(9, 8),
9791 => conv_std_logic_vector(9, 8),
9792 => conv_std_logic_vector(9, 8),
9793 => conv_std_logic_vector(9, 8),
9794 => conv_std_logic_vector(9, 8),
9795 => conv_std_logic_vector(9, 8),
9796 => conv_std_logic_vector(10, 8),
9797 => conv_std_logic_vector(10, 8),
9798 => conv_std_logic_vector(10, 8),
9799 => conv_std_logic_vector(10, 8),
9800 => conv_std_logic_vector(10, 8),
9801 => conv_std_logic_vector(10, 8),
9802 => conv_std_logic_vector(10, 8),
9803 => conv_std_logic_vector(11, 8),
9804 => conv_std_logic_vector(11, 8),
9805 => conv_std_logic_vector(11, 8),
9806 => conv_std_logic_vector(11, 8),
9807 => conv_std_logic_vector(11, 8),
9808 => conv_std_logic_vector(11, 8),
9809 => conv_std_logic_vector(12, 8),
9810 => conv_std_logic_vector(12, 8),
9811 => conv_std_logic_vector(12, 8),
9812 => conv_std_logic_vector(12, 8),
9813 => conv_std_logic_vector(12, 8),
9814 => conv_std_logic_vector(12, 8),
9815 => conv_std_logic_vector(12, 8),
9816 => conv_std_logic_vector(13, 8),
9817 => conv_std_logic_vector(13, 8),
9818 => conv_std_logic_vector(13, 8),
9819 => conv_std_logic_vector(13, 8),
9820 => conv_std_logic_vector(13, 8),
9821 => conv_std_logic_vector(13, 8),
9822 => conv_std_logic_vector(13, 8),
9823 => conv_std_logic_vector(14, 8),
9824 => conv_std_logic_vector(14, 8),
9825 => conv_std_logic_vector(14, 8),
9826 => conv_std_logic_vector(14, 8),
9827 => conv_std_logic_vector(14, 8),
9828 => conv_std_logic_vector(14, 8),
9829 => conv_std_logic_vector(14, 8),
9830 => conv_std_logic_vector(15, 8),
9831 => conv_std_logic_vector(15, 8),
9832 => conv_std_logic_vector(15, 8),
9833 => conv_std_logic_vector(15, 8),
9834 => conv_std_logic_vector(15, 8),
9835 => conv_std_logic_vector(15, 8),
9836 => conv_std_logic_vector(16, 8),
9837 => conv_std_logic_vector(16, 8),
9838 => conv_std_logic_vector(16, 8),
9839 => conv_std_logic_vector(16, 8),
9840 => conv_std_logic_vector(16, 8),
9841 => conv_std_logic_vector(16, 8),
9842 => conv_std_logic_vector(16, 8),
9843 => conv_std_logic_vector(17, 8),
9844 => conv_std_logic_vector(17, 8),
9845 => conv_std_logic_vector(17, 8),
9846 => conv_std_logic_vector(17, 8),
9847 => conv_std_logic_vector(17, 8),
9848 => conv_std_logic_vector(17, 8),
9849 => conv_std_logic_vector(17, 8),
9850 => conv_std_logic_vector(18, 8),
9851 => conv_std_logic_vector(18, 8),
9852 => conv_std_logic_vector(18, 8),
9853 => conv_std_logic_vector(18, 8),
9854 => conv_std_logic_vector(18, 8),
9855 => conv_std_logic_vector(18, 8),
9856 => conv_std_logic_vector(19, 8),
9857 => conv_std_logic_vector(19, 8),
9858 => conv_std_logic_vector(19, 8),
9859 => conv_std_logic_vector(19, 8),
9860 => conv_std_logic_vector(19, 8),
9861 => conv_std_logic_vector(19, 8),
9862 => conv_std_logic_vector(19, 8),
9863 => conv_std_logic_vector(20, 8),
9864 => conv_std_logic_vector(20, 8),
9865 => conv_std_logic_vector(20, 8),
9866 => conv_std_logic_vector(20, 8),
9867 => conv_std_logic_vector(20, 8),
9868 => conv_std_logic_vector(20, 8),
9869 => conv_std_logic_vector(20, 8),
9870 => conv_std_logic_vector(21, 8),
9871 => conv_std_logic_vector(21, 8),
9872 => conv_std_logic_vector(21, 8),
9873 => conv_std_logic_vector(21, 8),
9874 => conv_std_logic_vector(21, 8),
9875 => conv_std_logic_vector(21, 8),
9876 => conv_std_logic_vector(21, 8),
9877 => conv_std_logic_vector(22, 8),
9878 => conv_std_logic_vector(22, 8),
9879 => conv_std_logic_vector(22, 8),
9880 => conv_std_logic_vector(22, 8),
9881 => conv_std_logic_vector(22, 8),
9882 => conv_std_logic_vector(22, 8),
9883 => conv_std_logic_vector(23, 8),
9884 => conv_std_logic_vector(23, 8),
9885 => conv_std_logic_vector(23, 8),
9886 => conv_std_logic_vector(23, 8),
9887 => conv_std_logic_vector(23, 8),
9888 => conv_std_logic_vector(23, 8),
9889 => conv_std_logic_vector(23, 8),
9890 => conv_std_logic_vector(24, 8),
9891 => conv_std_logic_vector(24, 8),
9892 => conv_std_logic_vector(24, 8),
9893 => conv_std_logic_vector(24, 8),
9894 => conv_std_logic_vector(24, 8),
9895 => conv_std_logic_vector(24, 8),
9896 => conv_std_logic_vector(24, 8),
9897 => conv_std_logic_vector(25, 8),
9898 => conv_std_logic_vector(25, 8),
9899 => conv_std_logic_vector(25, 8),
9900 => conv_std_logic_vector(25, 8),
9901 => conv_std_logic_vector(25, 8),
9902 => conv_std_logic_vector(25, 8),
9903 => conv_std_logic_vector(25, 8),
9904 => conv_std_logic_vector(26, 8),
9905 => conv_std_logic_vector(26, 8),
9906 => conv_std_logic_vector(26, 8),
9907 => conv_std_logic_vector(26, 8),
9908 => conv_std_logic_vector(26, 8),
9909 => conv_std_logic_vector(26, 8),
9910 => conv_std_logic_vector(27, 8),
9911 => conv_std_logic_vector(27, 8),
9912 => conv_std_logic_vector(27, 8),
9913 => conv_std_logic_vector(27, 8),
9914 => conv_std_logic_vector(27, 8),
9915 => conv_std_logic_vector(27, 8),
9916 => conv_std_logic_vector(27, 8),
9917 => conv_std_logic_vector(28, 8),
9918 => conv_std_logic_vector(28, 8),
9919 => conv_std_logic_vector(28, 8),
9920 => conv_std_logic_vector(28, 8),
9921 => conv_std_logic_vector(28, 8),
9922 => conv_std_logic_vector(28, 8),
9923 => conv_std_logic_vector(28, 8),
9924 => conv_std_logic_vector(29, 8),
9925 => conv_std_logic_vector(29, 8),
9926 => conv_std_logic_vector(29, 8),
9927 => conv_std_logic_vector(29, 8),
9928 => conv_std_logic_vector(29, 8),
9929 => conv_std_logic_vector(29, 8),
9930 => conv_std_logic_vector(29, 8),
9931 => conv_std_logic_vector(30, 8),
9932 => conv_std_logic_vector(30, 8),
9933 => conv_std_logic_vector(30, 8),
9934 => conv_std_logic_vector(30, 8),
9935 => conv_std_logic_vector(30, 8),
9936 => conv_std_logic_vector(30, 8),
9937 => conv_std_logic_vector(31, 8),
9938 => conv_std_logic_vector(31, 8),
9939 => conv_std_logic_vector(31, 8),
9940 => conv_std_logic_vector(31, 8),
9941 => conv_std_logic_vector(31, 8),
9942 => conv_std_logic_vector(31, 8),
9943 => conv_std_logic_vector(31, 8),
9944 => conv_std_logic_vector(32, 8),
9945 => conv_std_logic_vector(32, 8),
9946 => conv_std_logic_vector(32, 8),
9947 => conv_std_logic_vector(32, 8),
9948 => conv_std_logic_vector(32, 8),
9949 => conv_std_logic_vector(32, 8),
9950 => conv_std_logic_vector(32, 8),
9951 => conv_std_logic_vector(33, 8),
9952 => conv_std_logic_vector(33, 8),
9953 => conv_std_logic_vector(33, 8),
9954 => conv_std_logic_vector(33, 8),
9955 => conv_std_logic_vector(33, 8),
9956 => conv_std_logic_vector(33, 8),
9957 => conv_std_logic_vector(33, 8),
9958 => conv_std_logic_vector(34, 8),
9959 => conv_std_logic_vector(34, 8),
9960 => conv_std_logic_vector(34, 8),
9961 => conv_std_logic_vector(34, 8),
9962 => conv_std_logic_vector(34, 8),
9963 => conv_std_logic_vector(34, 8),
9964 => conv_std_logic_vector(35, 8),
9965 => conv_std_logic_vector(35, 8),
9966 => conv_std_logic_vector(35, 8),
9967 => conv_std_logic_vector(35, 8),
9968 => conv_std_logic_vector(35, 8),
9969 => conv_std_logic_vector(35, 8),
9970 => conv_std_logic_vector(35, 8),
9971 => conv_std_logic_vector(36, 8),
9972 => conv_std_logic_vector(36, 8),
9973 => conv_std_logic_vector(36, 8),
9974 => conv_std_logic_vector(36, 8),
9975 => conv_std_logic_vector(36, 8),
9976 => conv_std_logic_vector(36, 8),
9977 => conv_std_logic_vector(36, 8),
9978 => conv_std_logic_vector(37, 8),
9979 => conv_std_logic_vector(37, 8),
9980 => conv_std_logic_vector(37, 8),
9981 => conv_std_logic_vector(37, 8),
9982 => conv_std_logic_vector(37, 8),
9983 => conv_std_logic_vector(37, 8),
9984 => conv_std_logic_vector(0, 8),
9985 => conv_std_logic_vector(0, 8),
9986 => conv_std_logic_vector(0, 8),
9987 => conv_std_logic_vector(0, 8),
9988 => conv_std_logic_vector(0, 8),
9989 => conv_std_logic_vector(0, 8),
9990 => conv_std_logic_vector(0, 8),
9991 => conv_std_logic_vector(1, 8),
9992 => conv_std_logic_vector(1, 8),
9993 => conv_std_logic_vector(1, 8),
9994 => conv_std_logic_vector(1, 8),
9995 => conv_std_logic_vector(1, 8),
9996 => conv_std_logic_vector(1, 8),
9997 => conv_std_logic_vector(1, 8),
9998 => conv_std_logic_vector(2, 8),
9999 => conv_std_logic_vector(2, 8),
10000 => conv_std_logic_vector(2, 8),
10001 => conv_std_logic_vector(2, 8),
10002 => conv_std_logic_vector(2, 8),
10003 => conv_std_logic_vector(2, 8),
10004 => conv_std_logic_vector(3, 8),
10005 => conv_std_logic_vector(3, 8),
10006 => conv_std_logic_vector(3, 8),
10007 => conv_std_logic_vector(3, 8),
10008 => conv_std_logic_vector(3, 8),
10009 => conv_std_logic_vector(3, 8),
10010 => conv_std_logic_vector(3, 8),
10011 => conv_std_logic_vector(4, 8),
10012 => conv_std_logic_vector(4, 8),
10013 => conv_std_logic_vector(4, 8),
10014 => conv_std_logic_vector(4, 8),
10015 => conv_std_logic_vector(4, 8),
10016 => conv_std_logic_vector(4, 8),
10017 => conv_std_logic_vector(5, 8),
10018 => conv_std_logic_vector(5, 8),
10019 => conv_std_logic_vector(5, 8),
10020 => conv_std_logic_vector(5, 8),
10021 => conv_std_logic_vector(5, 8),
10022 => conv_std_logic_vector(5, 8),
10023 => conv_std_logic_vector(5, 8),
10024 => conv_std_logic_vector(6, 8),
10025 => conv_std_logic_vector(6, 8),
10026 => conv_std_logic_vector(6, 8),
10027 => conv_std_logic_vector(6, 8),
10028 => conv_std_logic_vector(6, 8),
10029 => conv_std_logic_vector(6, 8),
10030 => conv_std_logic_vector(7, 8),
10031 => conv_std_logic_vector(7, 8),
10032 => conv_std_logic_vector(7, 8),
10033 => conv_std_logic_vector(7, 8),
10034 => conv_std_logic_vector(7, 8),
10035 => conv_std_logic_vector(7, 8),
10036 => conv_std_logic_vector(7, 8),
10037 => conv_std_logic_vector(8, 8),
10038 => conv_std_logic_vector(8, 8),
10039 => conv_std_logic_vector(8, 8),
10040 => conv_std_logic_vector(8, 8),
10041 => conv_std_logic_vector(8, 8),
10042 => conv_std_logic_vector(8, 8),
10043 => conv_std_logic_vector(8, 8),
10044 => conv_std_logic_vector(9, 8),
10045 => conv_std_logic_vector(9, 8),
10046 => conv_std_logic_vector(9, 8),
10047 => conv_std_logic_vector(9, 8),
10048 => conv_std_logic_vector(9, 8),
10049 => conv_std_logic_vector(9, 8),
10050 => conv_std_logic_vector(10, 8),
10051 => conv_std_logic_vector(10, 8),
10052 => conv_std_logic_vector(10, 8),
10053 => conv_std_logic_vector(10, 8),
10054 => conv_std_logic_vector(10, 8),
10055 => conv_std_logic_vector(10, 8),
10056 => conv_std_logic_vector(10, 8),
10057 => conv_std_logic_vector(11, 8),
10058 => conv_std_logic_vector(11, 8),
10059 => conv_std_logic_vector(11, 8),
10060 => conv_std_logic_vector(11, 8),
10061 => conv_std_logic_vector(11, 8),
10062 => conv_std_logic_vector(11, 8),
10063 => conv_std_logic_vector(12, 8),
10064 => conv_std_logic_vector(12, 8),
10065 => conv_std_logic_vector(12, 8),
10066 => conv_std_logic_vector(12, 8),
10067 => conv_std_logic_vector(12, 8),
10068 => conv_std_logic_vector(12, 8),
10069 => conv_std_logic_vector(12, 8),
10070 => conv_std_logic_vector(13, 8),
10071 => conv_std_logic_vector(13, 8),
10072 => conv_std_logic_vector(13, 8),
10073 => conv_std_logic_vector(13, 8),
10074 => conv_std_logic_vector(13, 8),
10075 => conv_std_logic_vector(13, 8),
10076 => conv_std_logic_vector(14, 8),
10077 => conv_std_logic_vector(14, 8),
10078 => conv_std_logic_vector(14, 8),
10079 => conv_std_logic_vector(14, 8),
10080 => conv_std_logic_vector(14, 8),
10081 => conv_std_logic_vector(14, 8),
10082 => conv_std_logic_vector(14, 8),
10083 => conv_std_logic_vector(15, 8),
10084 => conv_std_logic_vector(15, 8),
10085 => conv_std_logic_vector(15, 8),
10086 => conv_std_logic_vector(15, 8),
10087 => conv_std_logic_vector(15, 8),
10088 => conv_std_logic_vector(15, 8),
10089 => conv_std_logic_vector(15, 8),
10090 => conv_std_logic_vector(16, 8),
10091 => conv_std_logic_vector(16, 8),
10092 => conv_std_logic_vector(16, 8),
10093 => conv_std_logic_vector(16, 8),
10094 => conv_std_logic_vector(16, 8),
10095 => conv_std_logic_vector(16, 8),
10096 => conv_std_logic_vector(17, 8),
10097 => conv_std_logic_vector(17, 8),
10098 => conv_std_logic_vector(17, 8),
10099 => conv_std_logic_vector(17, 8),
10100 => conv_std_logic_vector(17, 8),
10101 => conv_std_logic_vector(17, 8),
10102 => conv_std_logic_vector(17, 8),
10103 => conv_std_logic_vector(18, 8),
10104 => conv_std_logic_vector(18, 8),
10105 => conv_std_logic_vector(18, 8),
10106 => conv_std_logic_vector(18, 8),
10107 => conv_std_logic_vector(18, 8),
10108 => conv_std_logic_vector(18, 8),
10109 => conv_std_logic_vector(19, 8),
10110 => conv_std_logic_vector(19, 8),
10111 => conv_std_logic_vector(19, 8),
10112 => conv_std_logic_vector(19, 8),
10113 => conv_std_logic_vector(19, 8),
10114 => conv_std_logic_vector(19, 8),
10115 => conv_std_logic_vector(19, 8),
10116 => conv_std_logic_vector(20, 8),
10117 => conv_std_logic_vector(20, 8),
10118 => conv_std_logic_vector(20, 8),
10119 => conv_std_logic_vector(20, 8),
10120 => conv_std_logic_vector(20, 8),
10121 => conv_std_logic_vector(20, 8),
10122 => conv_std_logic_vector(21, 8),
10123 => conv_std_logic_vector(21, 8),
10124 => conv_std_logic_vector(21, 8),
10125 => conv_std_logic_vector(21, 8),
10126 => conv_std_logic_vector(21, 8),
10127 => conv_std_logic_vector(21, 8),
10128 => conv_std_logic_vector(21, 8),
10129 => conv_std_logic_vector(22, 8),
10130 => conv_std_logic_vector(22, 8),
10131 => conv_std_logic_vector(22, 8),
10132 => conv_std_logic_vector(22, 8),
10133 => conv_std_logic_vector(22, 8),
10134 => conv_std_logic_vector(22, 8),
10135 => conv_std_logic_vector(23, 8),
10136 => conv_std_logic_vector(23, 8),
10137 => conv_std_logic_vector(23, 8),
10138 => conv_std_logic_vector(23, 8),
10139 => conv_std_logic_vector(23, 8),
10140 => conv_std_logic_vector(23, 8),
10141 => conv_std_logic_vector(23, 8),
10142 => conv_std_logic_vector(24, 8),
10143 => conv_std_logic_vector(24, 8),
10144 => conv_std_logic_vector(24, 8),
10145 => conv_std_logic_vector(24, 8),
10146 => conv_std_logic_vector(24, 8),
10147 => conv_std_logic_vector(24, 8),
10148 => conv_std_logic_vector(24, 8),
10149 => conv_std_logic_vector(25, 8),
10150 => conv_std_logic_vector(25, 8),
10151 => conv_std_logic_vector(25, 8),
10152 => conv_std_logic_vector(25, 8),
10153 => conv_std_logic_vector(25, 8),
10154 => conv_std_logic_vector(25, 8),
10155 => conv_std_logic_vector(26, 8),
10156 => conv_std_logic_vector(26, 8),
10157 => conv_std_logic_vector(26, 8),
10158 => conv_std_logic_vector(26, 8),
10159 => conv_std_logic_vector(26, 8),
10160 => conv_std_logic_vector(26, 8),
10161 => conv_std_logic_vector(26, 8),
10162 => conv_std_logic_vector(27, 8),
10163 => conv_std_logic_vector(27, 8),
10164 => conv_std_logic_vector(27, 8),
10165 => conv_std_logic_vector(27, 8),
10166 => conv_std_logic_vector(27, 8),
10167 => conv_std_logic_vector(27, 8),
10168 => conv_std_logic_vector(28, 8),
10169 => conv_std_logic_vector(28, 8),
10170 => conv_std_logic_vector(28, 8),
10171 => conv_std_logic_vector(28, 8),
10172 => conv_std_logic_vector(28, 8),
10173 => conv_std_logic_vector(28, 8),
10174 => conv_std_logic_vector(28, 8),
10175 => conv_std_logic_vector(29, 8),
10176 => conv_std_logic_vector(29, 8),
10177 => conv_std_logic_vector(29, 8),
10178 => conv_std_logic_vector(29, 8),
10179 => conv_std_logic_vector(29, 8),
10180 => conv_std_logic_vector(29, 8),
10181 => conv_std_logic_vector(30, 8),
10182 => conv_std_logic_vector(30, 8),
10183 => conv_std_logic_vector(30, 8),
10184 => conv_std_logic_vector(30, 8),
10185 => conv_std_logic_vector(30, 8),
10186 => conv_std_logic_vector(30, 8),
10187 => conv_std_logic_vector(30, 8),
10188 => conv_std_logic_vector(31, 8),
10189 => conv_std_logic_vector(31, 8),
10190 => conv_std_logic_vector(31, 8),
10191 => conv_std_logic_vector(31, 8),
10192 => conv_std_logic_vector(31, 8),
10193 => conv_std_logic_vector(31, 8),
10194 => conv_std_logic_vector(31, 8),
10195 => conv_std_logic_vector(32, 8),
10196 => conv_std_logic_vector(32, 8),
10197 => conv_std_logic_vector(32, 8),
10198 => conv_std_logic_vector(32, 8),
10199 => conv_std_logic_vector(32, 8),
10200 => conv_std_logic_vector(32, 8),
10201 => conv_std_logic_vector(33, 8),
10202 => conv_std_logic_vector(33, 8),
10203 => conv_std_logic_vector(33, 8),
10204 => conv_std_logic_vector(33, 8),
10205 => conv_std_logic_vector(33, 8),
10206 => conv_std_logic_vector(33, 8),
10207 => conv_std_logic_vector(33, 8),
10208 => conv_std_logic_vector(34, 8),
10209 => conv_std_logic_vector(34, 8),
10210 => conv_std_logic_vector(34, 8),
10211 => conv_std_logic_vector(34, 8),
10212 => conv_std_logic_vector(34, 8),
10213 => conv_std_logic_vector(34, 8),
10214 => conv_std_logic_vector(35, 8),
10215 => conv_std_logic_vector(35, 8),
10216 => conv_std_logic_vector(35, 8),
10217 => conv_std_logic_vector(35, 8),
10218 => conv_std_logic_vector(35, 8),
10219 => conv_std_logic_vector(35, 8),
10220 => conv_std_logic_vector(35, 8),
10221 => conv_std_logic_vector(36, 8),
10222 => conv_std_logic_vector(36, 8),
10223 => conv_std_logic_vector(36, 8),
10224 => conv_std_logic_vector(36, 8),
10225 => conv_std_logic_vector(36, 8),
10226 => conv_std_logic_vector(36, 8),
10227 => conv_std_logic_vector(37, 8),
10228 => conv_std_logic_vector(37, 8),
10229 => conv_std_logic_vector(37, 8),
10230 => conv_std_logic_vector(37, 8),
10231 => conv_std_logic_vector(37, 8),
10232 => conv_std_logic_vector(37, 8),
10233 => conv_std_logic_vector(37, 8),
10234 => conv_std_logic_vector(38, 8),
10235 => conv_std_logic_vector(38, 8),
10236 => conv_std_logic_vector(38, 8),
10237 => conv_std_logic_vector(38, 8),
10238 => conv_std_logic_vector(38, 8),
10239 => conv_std_logic_vector(38, 8),
10240 => conv_std_logic_vector(0, 8),
10241 => conv_std_logic_vector(0, 8),
10242 => conv_std_logic_vector(0, 8),
10243 => conv_std_logic_vector(0, 8),
10244 => conv_std_logic_vector(0, 8),
10245 => conv_std_logic_vector(0, 8),
10246 => conv_std_logic_vector(0, 8),
10247 => conv_std_logic_vector(1, 8),
10248 => conv_std_logic_vector(1, 8),
10249 => conv_std_logic_vector(1, 8),
10250 => conv_std_logic_vector(1, 8),
10251 => conv_std_logic_vector(1, 8),
10252 => conv_std_logic_vector(1, 8),
10253 => conv_std_logic_vector(2, 8),
10254 => conv_std_logic_vector(2, 8),
10255 => conv_std_logic_vector(2, 8),
10256 => conv_std_logic_vector(2, 8),
10257 => conv_std_logic_vector(2, 8),
10258 => conv_std_logic_vector(2, 8),
10259 => conv_std_logic_vector(2, 8),
10260 => conv_std_logic_vector(3, 8),
10261 => conv_std_logic_vector(3, 8),
10262 => conv_std_logic_vector(3, 8),
10263 => conv_std_logic_vector(3, 8),
10264 => conv_std_logic_vector(3, 8),
10265 => conv_std_logic_vector(3, 8),
10266 => conv_std_logic_vector(4, 8),
10267 => conv_std_logic_vector(4, 8),
10268 => conv_std_logic_vector(4, 8),
10269 => conv_std_logic_vector(4, 8),
10270 => conv_std_logic_vector(4, 8),
10271 => conv_std_logic_vector(4, 8),
10272 => conv_std_logic_vector(5, 8),
10273 => conv_std_logic_vector(5, 8),
10274 => conv_std_logic_vector(5, 8),
10275 => conv_std_logic_vector(5, 8),
10276 => conv_std_logic_vector(5, 8),
10277 => conv_std_logic_vector(5, 8),
10278 => conv_std_logic_vector(5, 8),
10279 => conv_std_logic_vector(6, 8),
10280 => conv_std_logic_vector(6, 8),
10281 => conv_std_logic_vector(6, 8),
10282 => conv_std_logic_vector(6, 8),
10283 => conv_std_logic_vector(6, 8),
10284 => conv_std_logic_vector(6, 8),
10285 => conv_std_logic_vector(7, 8),
10286 => conv_std_logic_vector(7, 8),
10287 => conv_std_logic_vector(7, 8),
10288 => conv_std_logic_vector(7, 8),
10289 => conv_std_logic_vector(7, 8),
10290 => conv_std_logic_vector(7, 8),
10291 => conv_std_logic_vector(7, 8),
10292 => conv_std_logic_vector(8, 8),
10293 => conv_std_logic_vector(8, 8),
10294 => conv_std_logic_vector(8, 8),
10295 => conv_std_logic_vector(8, 8),
10296 => conv_std_logic_vector(8, 8),
10297 => conv_std_logic_vector(8, 8),
10298 => conv_std_logic_vector(9, 8),
10299 => conv_std_logic_vector(9, 8),
10300 => conv_std_logic_vector(9, 8),
10301 => conv_std_logic_vector(9, 8),
10302 => conv_std_logic_vector(9, 8),
10303 => conv_std_logic_vector(9, 8),
10304 => conv_std_logic_vector(10, 8),
10305 => conv_std_logic_vector(10, 8),
10306 => conv_std_logic_vector(10, 8),
10307 => conv_std_logic_vector(10, 8),
10308 => conv_std_logic_vector(10, 8),
10309 => conv_std_logic_vector(10, 8),
10310 => conv_std_logic_vector(10, 8),
10311 => conv_std_logic_vector(11, 8),
10312 => conv_std_logic_vector(11, 8),
10313 => conv_std_logic_vector(11, 8),
10314 => conv_std_logic_vector(11, 8),
10315 => conv_std_logic_vector(11, 8),
10316 => conv_std_logic_vector(11, 8),
10317 => conv_std_logic_vector(12, 8),
10318 => conv_std_logic_vector(12, 8),
10319 => conv_std_logic_vector(12, 8),
10320 => conv_std_logic_vector(12, 8),
10321 => conv_std_logic_vector(12, 8),
10322 => conv_std_logic_vector(12, 8),
10323 => conv_std_logic_vector(12, 8),
10324 => conv_std_logic_vector(13, 8),
10325 => conv_std_logic_vector(13, 8),
10326 => conv_std_logic_vector(13, 8),
10327 => conv_std_logic_vector(13, 8),
10328 => conv_std_logic_vector(13, 8),
10329 => conv_std_logic_vector(13, 8),
10330 => conv_std_logic_vector(14, 8),
10331 => conv_std_logic_vector(14, 8),
10332 => conv_std_logic_vector(14, 8),
10333 => conv_std_logic_vector(14, 8),
10334 => conv_std_logic_vector(14, 8),
10335 => conv_std_logic_vector(14, 8),
10336 => conv_std_logic_vector(15, 8),
10337 => conv_std_logic_vector(15, 8),
10338 => conv_std_logic_vector(15, 8),
10339 => conv_std_logic_vector(15, 8),
10340 => conv_std_logic_vector(15, 8),
10341 => conv_std_logic_vector(15, 8),
10342 => conv_std_logic_vector(15, 8),
10343 => conv_std_logic_vector(16, 8),
10344 => conv_std_logic_vector(16, 8),
10345 => conv_std_logic_vector(16, 8),
10346 => conv_std_logic_vector(16, 8),
10347 => conv_std_logic_vector(16, 8),
10348 => conv_std_logic_vector(16, 8),
10349 => conv_std_logic_vector(17, 8),
10350 => conv_std_logic_vector(17, 8),
10351 => conv_std_logic_vector(17, 8),
10352 => conv_std_logic_vector(17, 8),
10353 => conv_std_logic_vector(17, 8),
10354 => conv_std_logic_vector(17, 8),
10355 => conv_std_logic_vector(17, 8),
10356 => conv_std_logic_vector(18, 8),
10357 => conv_std_logic_vector(18, 8),
10358 => conv_std_logic_vector(18, 8),
10359 => conv_std_logic_vector(18, 8),
10360 => conv_std_logic_vector(18, 8),
10361 => conv_std_logic_vector(18, 8),
10362 => conv_std_logic_vector(19, 8),
10363 => conv_std_logic_vector(19, 8),
10364 => conv_std_logic_vector(19, 8),
10365 => conv_std_logic_vector(19, 8),
10366 => conv_std_logic_vector(19, 8),
10367 => conv_std_logic_vector(19, 8),
10368 => conv_std_logic_vector(20, 8),
10369 => conv_std_logic_vector(20, 8),
10370 => conv_std_logic_vector(20, 8),
10371 => conv_std_logic_vector(20, 8),
10372 => conv_std_logic_vector(20, 8),
10373 => conv_std_logic_vector(20, 8),
10374 => conv_std_logic_vector(20, 8),
10375 => conv_std_logic_vector(21, 8),
10376 => conv_std_logic_vector(21, 8),
10377 => conv_std_logic_vector(21, 8),
10378 => conv_std_logic_vector(21, 8),
10379 => conv_std_logic_vector(21, 8),
10380 => conv_std_logic_vector(21, 8),
10381 => conv_std_logic_vector(22, 8),
10382 => conv_std_logic_vector(22, 8),
10383 => conv_std_logic_vector(22, 8),
10384 => conv_std_logic_vector(22, 8),
10385 => conv_std_logic_vector(22, 8),
10386 => conv_std_logic_vector(22, 8),
10387 => conv_std_logic_vector(22, 8),
10388 => conv_std_logic_vector(23, 8),
10389 => conv_std_logic_vector(23, 8),
10390 => conv_std_logic_vector(23, 8),
10391 => conv_std_logic_vector(23, 8),
10392 => conv_std_logic_vector(23, 8),
10393 => conv_std_logic_vector(23, 8),
10394 => conv_std_logic_vector(24, 8),
10395 => conv_std_logic_vector(24, 8),
10396 => conv_std_logic_vector(24, 8),
10397 => conv_std_logic_vector(24, 8),
10398 => conv_std_logic_vector(24, 8),
10399 => conv_std_logic_vector(24, 8),
10400 => conv_std_logic_vector(25, 8),
10401 => conv_std_logic_vector(25, 8),
10402 => conv_std_logic_vector(25, 8),
10403 => conv_std_logic_vector(25, 8),
10404 => conv_std_logic_vector(25, 8),
10405 => conv_std_logic_vector(25, 8),
10406 => conv_std_logic_vector(25, 8),
10407 => conv_std_logic_vector(26, 8),
10408 => conv_std_logic_vector(26, 8),
10409 => conv_std_logic_vector(26, 8),
10410 => conv_std_logic_vector(26, 8),
10411 => conv_std_logic_vector(26, 8),
10412 => conv_std_logic_vector(26, 8),
10413 => conv_std_logic_vector(27, 8),
10414 => conv_std_logic_vector(27, 8),
10415 => conv_std_logic_vector(27, 8),
10416 => conv_std_logic_vector(27, 8),
10417 => conv_std_logic_vector(27, 8),
10418 => conv_std_logic_vector(27, 8),
10419 => conv_std_logic_vector(27, 8),
10420 => conv_std_logic_vector(28, 8),
10421 => conv_std_logic_vector(28, 8),
10422 => conv_std_logic_vector(28, 8),
10423 => conv_std_logic_vector(28, 8),
10424 => conv_std_logic_vector(28, 8),
10425 => conv_std_logic_vector(28, 8),
10426 => conv_std_logic_vector(29, 8),
10427 => conv_std_logic_vector(29, 8),
10428 => conv_std_logic_vector(29, 8),
10429 => conv_std_logic_vector(29, 8),
10430 => conv_std_logic_vector(29, 8),
10431 => conv_std_logic_vector(29, 8),
10432 => conv_std_logic_vector(30, 8),
10433 => conv_std_logic_vector(30, 8),
10434 => conv_std_logic_vector(30, 8),
10435 => conv_std_logic_vector(30, 8),
10436 => conv_std_logic_vector(30, 8),
10437 => conv_std_logic_vector(30, 8),
10438 => conv_std_logic_vector(30, 8),
10439 => conv_std_logic_vector(31, 8),
10440 => conv_std_logic_vector(31, 8),
10441 => conv_std_logic_vector(31, 8),
10442 => conv_std_logic_vector(31, 8),
10443 => conv_std_logic_vector(31, 8),
10444 => conv_std_logic_vector(31, 8),
10445 => conv_std_logic_vector(32, 8),
10446 => conv_std_logic_vector(32, 8),
10447 => conv_std_logic_vector(32, 8),
10448 => conv_std_logic_vector(32, 8),
10449 => conv_std_logic_vector(32, 8),
10450 => conv_std_logic_vector(32, 8),
10451 => conv_std_logic_vector(32, 8),
10452 => conv_std_logic_vector(33, 8),
10453 => conv_std_logic_vector(33, 8),
10454 => conv_std_logic_vector(33, 8),
10455 => conv_std_logic_vector(33, 8),
10456 => conv_std_logic_vector(33, 8),
10457 => conv_std_logic_vector(33, 8),
10458 => conv_std_logic_vector(34, 8),
10459 => conv_std_logic_vector(34, 8),
10460 => conv_std_logic_vector(34, 8),
10461 => conv_std_logic_vector(34, 8),
10462 => conv_std_logic_vector(34, 8),
10463 => conv_std_logic_vector(34, 8),
10464 => conv_std_logic_vector(35, 8),
10465 => conv_std_logic_vector(35, 8),
10466 => conv_std_logic_vector(35, 8),
10467 => conv_std_logic_vector(35, 8),
10468 => conv_std_logic_vector(35, 8),
10469 => conv_std_logic_vector(35, 8),
10470 => conv_std_logic_vector(35, 8),
10471 => conv_std_logic_vector(36, 8),
10472 => conv_std_logic_vector(36, 8),
10473 => conv_std_logic_vector(36, 8),
10474 => conv_std_logic_vector(36, 8),
10475 => conv_std_logic_vector(36, 8),
10476 => conv_std_logic_vector(36, 8),
10477 => conv_std_logic_vector(37, 8),
10478 => conv_std_logic_vector(37, 8),
10479 => conv_std_logic_vector(37, 8),
10480 => conv_std_logic_vector(37, 8),
10481 => conv_std_logic_vector(37, 8),
10482 => conv_std_logic_vector(37, 8),
10483 => conv_std_logic_vector(37, 8),
10484 => conv_std_logic_vector(38, 8),
10485 => conv_std_logic_vector(38, 8),
10486 => conv_std_logic_vector(38, 8),
10487 => conv_std_logic_vector(38, 8),
10488 => conv_std_logic_vector(38, 8),
10489 => conv_std_logic_vector(38, 8),
10490 => conv_std_logic_vector(39, 8),
10491 => conv_std_logic_vector(39, 8),
10492 => conv_std_logic_vector(39, 8),
10493 => conv_std_logic_vector(39, 8),
10494 => conv_std_logic_vector(39, 8),
10495 => conv_std_logic_vector(39, 8),
10496 => conv_std_logic_vector(0, 8),
10497 => conv_std_logic_vector(0, 8),
10498 => conv_std_logic_vector(0, 8),
10499 => conv_std_logic_vector(0, 8),
10500 => conv_std_logic_vector(0, 8),
10501 => conv_std_logic_vector(0, 8),
10502 => conv_std_logic_vector(0, 8),
10503 => conv_std_logic_vector(1, 8),
10504 => conv_std_logic_vector(1, 8),
10505 => conv_std_logic_vector(1, 8),
10506 => conv_std_logic_vector(1, 8),
10507 => conv_std_logic_vector(1, 8),
10508 => conv_std_logic_vector(1, 8),
10509 => conv_std_logic_vector(2, 8),
10510 => conv_std_logic_vector(2, 8),
10511 => conv_std_logic_vector(2, 8),
10512 => conv_std_logic_vector(2, 8),
10513 => conv_std_logic_vector(2, 8),
10514 => conv_std_logic_vector(2, 8),
10515 => conv_std_logic_vector(3, 8),
10516 => conv_std_logic_vector(3, 8),
10517 => conv_std_logic_vector(3, 8),
10518 => conv_std_logic_vector(3, 8),
10519 => conv_std_logic_vector(3, 8),
10520 => conv_std_logic_vector(3, 8),
10521 => conv_std_logic_vector(4, 8),
10522 => conv_std_logic_vector(4, 8),
10523 => conv_std_logic_vector(4, 8),
10524 => conv_std_logic_vector(4, 8),
10525 => conv_std_logic_vector(4, 8),
10526 => conv_std_logic_vector(4, 8),
10527 => conv_std_logic_vector(4, 8),
10528 => conv_std_logic_vector(5, 8),
10529 => conv_std_logic_vector(5, 8),
10530 => conv_std_logic_vector(5, 8),
10531 => conv_std_logic_vector(5, 8),
10532 => conv_std_logic_vector(5, 8),
10533 => conv_std_logic_vector(5, 8),
10534 => conv_std_logic_vector(6, 8),
10535 => conv_std_logic_vector(6, 8),
10536 => conv_std_logic_vector(6, 8),
10537 => conv_std_logic_vector(6, 8),
10538 => conv_std_logic_vector(6, 8),
10539 => conv_std_logic_vector(6, 8),
10540 => conv_std_logic_vector(7, 8),
10541 => conv_std_logic_vector(7, 8),
10542 => conv_std_logic_vector(7, 8),
10543 => conv_std_logic_vector(7, 8),
10544 => conv_std_logic_vector(7, 8),
10545 => conv_std_logic_vector(7, 8),
10546 => conv_std_logic_vector(8, 8),
10547 => conv_std_logic_vector(8, 8),
10548 => conv_std_logic_vector(8, 8),
10549 => conv_std_logic_vector(8, 8),
10550 => conv_std_logic_vector(8, 8),
10551 => conv_std_logic_vector(8, 8),
10552 => conv_std_logic_vector(8, 8),
10553 => conv_std_logic_vector(9, 8),
10554 => conv_std_logic_vector(9, 8),
10555 => conv_std_logic_vector(9, 8),
10556 => conv_std_logic_vector(9, 8),
10557 => conv_std_logic_vector(9, 8),
10558 => conv_std_logic_vector(9, 8),
10559 => conv_std_logic_vector(10, 8),
10560 => conv_std_logic_vector(10, 8),
10561 => conv_std_logic_vector(10, 8),
10562 => conv_std_logic_vector(10, 8),
10563 => conv_std_logic_vector(10, 8),
10564 => conv_std_logic_vector(10, 8),
10565 => conv_std_logic_vector(11, 8),
10566 => conv_std_logic_vector(11, 8),
10567 => conv_std_logic_vector(11, 8),
10568 => conv_std_logic_vector(11, 8),
10569 => conv_std_logic_vector(11, 8),
10570 => conv_std_logic_vector(11, 8),
10571 => conv_std_logic_vector(12, 8),
10572 => conv_std_logic_vector(12, 8),
10573 => conv_std_logic_vector(12, 8),
10574 => conv_std_logic_vector(12, 8),
10575 => conv_std_logic_vector(12, 8),
10576 => conv_std_logic_vector(12, 8),
10577 => conv_std_logic_vector(12, 8),
10578 => conv_std_logic_vector(13, 8),
10579 => conv_std_logic_vector(13, 8),
10580 => conv_std_logic_vector(13, 8),
10581 => conv_std_logic_vector(13, 8),
10582 => conv_std_logic_vector(13, 8),
10583 => conv_std_logic_vector(13, 8),
10584 => conv_std_logic_vector(14, 8),
10585 => conv_std_logic_vector(14, 8),
10586 => conv_std_logic_vector(14, 8),
10587 => conv_std_logic_vector(14, 8),
10588 => conv_std_logic_vector(14, 8),
10589 => conv_std_logic_vector(14, 8),
10590 => conv_std_logic_vector(15, 8),
10591 => conv_std_logic_vector(15, 8),
10592 => conv_std_logic_vector(15, 8),
10593 => conv_std_logic_vector(15, 8),
10594 => conv_std_logic_vector(15, 8),
10595 => conv_std_logic_vector(15, 8),
10596 => conv_std_logic_vector(16, 8),
10597 => conv_std_logic_vector(16, 8),
10598 => conv_std_logic_vector(16, 8),
10599 => conv_std_logic_vector(16, 8),
10600 => conv_std_logic_vector(16, 8),
10601 => conv_std_logic_vector(16, 8),
10602 => conv_std_logic_vector(16, 8),
10603 => conv_std_logic_vector(17, 8),
10604 => conv_std_logic_vector(17, 8),
10605 => conv_std_logic_vector(17, 8),
10606 => conv_std_logic_vector(17, 8),
10607 => conv_std_logic_vector(17, 8),
10608 => conv_std_logic_vector(17, 8),
10609 => conv_std_logic_vector(18, 8),
10610 => conv_std_logic_vector(18, 8),
10611 => conv_std_logic_vector(18, 8),
10612 => conv_std_logic_vector(18, 8),
10613 => conv_std_logic_vector(18, 8),
10614 => conv_std_logic_vector(18, 8),
10615 => conv_std_logic_vector(19, 8),
10616 => conv_std_logic_vector(19, 8),
10617 => conv_std_logic_vector(19, 8),
10618 => conv_std_logic_vector(19, 8),
10619 => conv_std_logic_vector(19, 8),
10620 => conv_std_logic_vector(19, 8),
10621 => conv_std_logic_vector(20, 8),
10622 => conv_std_logic_vector(20, 8),
10623 => conv_std_logic_vector(20, 8),
10624 => conv_std_logic_vector(20, 8),
10625 => conv_std_logic_vector(20, 8),
10626 => conv_std_logic_vector(20, 8),
10627 => conv_std_logic_vector(20, 8),
10628 => conv_std_logic_vector(21, 8),
10629 => conv_std_logic_vector(21, 8),
10630 => conv_std_logic_vector(21, 8),
10631 => conv_std_logic_vector(21, 8),
10632 => conv_std_logic_vector(21, 8),
10633 => conv_std_logic_vector(21, 8),
10634 => conv_std_logic_vector(22, 8),
10635 => conv_std_logic_vector(22, 8),
10636 => conv_std_logic_vector(22, 8),
10637 => conv_std_logic_vector(22, 8),
10638 => conv_std_logic_vector(22, 8),
10639 => conv_std_logic_vector(22, 8),
10640 => conv_std_logic_vector(23, 8),
10641 => conv_std_logic_vector(23, 8),
10642 => conv_std_logic_vector(23, 8),
10643 => conv_std_logic_vector(23, 8),
10644 => conv_std_logic_vector(23, 8),
10645 => conv_std_logic_vector(23, 8),
10646 => conv_std_logic_vector(24, 8),
10647 => conv_std_logic_vector(24, 8),
10648 => conv_std_logic_vector(24, 8),
10649 => conv_std_logic_vector(24, 8),
10650 => conv_std_logic_vector(24, 8),
10651 => conv_std_logic_vector(24, 8),
10652 => conv_std_logic_vector(24, 8),
10653 => conv_std_logic_vector(25, 8),
10654 => conv_std_logic_vector(25, 8),
10655 => conv_std_logic_vector(25, 8),
10656 => conv_std_logic_vector(25, 8),
10657 => conv_std_logic_vector(25, 8),
10658 => conv_std_logic_vector(25, 8),
10659 => conv_std_logic_vector(26, 8),
10660 => conv_std_logic_vector(26, 8),
10661 => conv_std_logic_vector(26, 8),
10662 => conv_std_logic_vector(26, 8),
10663 => conv_std_logic_vector(26, 8),
10664 => conv_std_logic_vector(26, 8),
10665 => conv_std_logic_vector(27, 8),
10666 => conv_std_logic_vector(27, 8),
10667 => conv_std_logic_vector(27, 8),
10668 => conv_std_logic_vector(27, 8),
10669 => conv_std_logic_vector(27, 8),
10670 => conv_std_logic_vector(27, 8),
10671 => conv_std_logic_vector(28, 8),
10672 => conv_std_logic_vector(28, 8),
10673 => conv_std_logic_vector(28, 8),
10674 => conv_std_logic_vector(28, 8),
10675 => conv_std_logic_vector(28, 8),
10676 => conv_std_logic_vector(28, 8),
10677 => conv_std_logic_vector(28, 8),
10678 => conv_std_logic_vector(29, 8),
10679 => conv_std_logic_vector(29, 8),
10680 => conv_std_logic_vector(29, 8),
10681 => conv_std_logic_vector(29, 8),
10682 => conv_std_logic_vector(29, 8),
10683 => conv_std_logic_vector(29, 8),
10684 => conv_std_logic_vector(30, 8),
10685 => conv_std_logic_vector(30, 8),
10686 => conv_std_logic_vector(30, 8),
10687 => conv_std_logic_vector(30, 8),
10688 => conv_std_logic_vector(30, 8),
10689 => conv_std_logic_vector(30, 8),
10690 => conv_std_logic_vector(31, 8),
10691 => conv_std_logic_vector(31, 8),
10692 => conv_std_logic_vector(31, 8),
10693 => conv_std_logic_vector(31, 8),
10694 => conv_std_logic_vector(31, 8),
10695 => conv_std_logic_vector(31, 8),
10696 => conv_std_logic_vector(32, 8),
10697 => conv_std_logic_vector(32, 8),
10698 => conv_std_logic_vector(32, 8),
10699 => conv_std_logic_vector(32, 8),
10700 => conv_std_logic_vector(32, 8),
10701 => conv_std_logic_vector(32, 8),
10702 => conv_std_logic_vector(32, 8),
10703 => conv_std_logic_vector(33, 8),
10704 => conv_std_logic_vector(33, 8),
10705 => conv_std_logic_vector(33, 8),
10706 => conv_std_logic_vector(33, 8),
10707 => conv_std_logic_vector(33, 8),
10708 => conv_std_logic_vector(33, 8),
10709 => conv_std_logic_vector(34, 8),
10710 => conv_std_logic_vector(34, 8),
10711 => conv_std_logic_vector(34, 8),
10712 => conv_std_logic_vector(34, 8),
10713 => conv_std_logic_vector(34, 8),
10714 => conv_std_logic_vector(34, 8),
10715 => conv_std_logic_vector(35, 8),
10716 => conv_std_logic_vector(35, 8),
10717 => conv_std_logic_vector(35, 8),
10718 => conv_std_logic_vector(35, 8),
10719 => conv_std_logic_vector(35, 8),
10720 => conv_std_logic_vector(35, 8),
10721 => conv_std_logic_vector(36, 8),
10722 => conv_std_logic_vector(36, 8),
10723 => conv_std_logic_vector(36, 8),
10724 => conv_std_logic_vector(36, 8),
10725 => conv_std_logic_vector(36, 8),
10726 => conv_std_logic_vector(36, 8),
10727 => conv_std_logic_vector(36, 8),
10728 => conv_std_logic_vector(37, 8),
10729 => conv_std_logic_vector(37, 8),
10730 => conv_std_logic_vector(37, 8),
10731 => conv_std_logic_vector(37, 8),
10732 => conv_std_logic_vector(37, 8),
10733 => conv_std_logic_vector(37, 8),
10734 => conv_std_logic_vector(38, 8),
10735 => conv_std_logic_vector(38, 8),
10736 => conv_std_logic_vector(38, 8),
10737 => conv_std_logic_vector(38, 8),
10738 => conv_std_logic_vector(38, 8),
10739 => conv_std_logic_vector(38, 8),
10740 => conv_std_logic_vector(39, 8),
10741 => conv_std_logic_vector(39, 8),
10742 => conv_std_logic_vector(39, 8),
10743 => conv_std_logic_vector(39, 8),
10744 => conv_std_logic_vector(39, 8),
10745 => conv_std_logic_vector(39, 8),
10746 => conv_std_logic_vector(40, 8),
10747 => conv_std_logic_vector(40, 8),
10748 => conv_std_logic_vector(40, 8),
10749 => conv_std_logic_vector(40, 8),
10750 => conv_std_logic_vector(40, 8),
10751 => conv_std_logic_vector(40, 8),
10752 => conv_std_logic_vector(0, 8),
10753 => conv_std_logic_vector(0, 8),
10754 => conv_std_logic_vector(0, 8),
10755 => conv_std_logic_vector(0, 8),
10756 => conv_std_logic_vector(0, 8),
10757 => conv_std_logic_vector(0, 8),
10758 => conv_std_logic_vector(0, 8),
10759 => conv_std_logic_vector(1, 8),
10760 => conv_std_logic_vector(1, 8),
10761 => conv_std_logic_vector(1, 8),
10762 => conv_std_logic_vector(1, 8),
10763 => conv_std_logic_vector(1, 8),
10764 => conv_std_logic_vector(1, 8),
10765 => conv_std_logic_vector(2, 8),
10766 => conv_std_logic_vector(2, 8),
10767 => conv_std_logic_vector(2, 8),
10768 => conv_std_logic_vector(2, 8),
10769 => conv_std_logic_vector(2, 8),
10770 => conv_std_logic_vector(2, 8),
10771 => conv_std_logic_vector(3, 8),
10772 => conv_std_logic_vector(3, 8),
10773 => conv_std_logic_vector(3, 8),
10774 => conv_std_logic_vector(3, 8),
10775 => conv_std_logic_vector(3, 8),
10776 => conv_std_logic_vector(3, 8),
10777 => conv_std_logic_vector(4, 8),
10778 => conv_std_logic_vector(4, 8),
10779 => conv_std_logic_vector(4, 8),
10780 => conv_std_logic_vector(4, 8),
10781 => conv_std_logic_vector(4, 8),
10782 => conv_std_logic_vector(4, 8),
10783 => conv_std_logic_vector(5, 8),
10784 => conv_std_logic_vector(5, 8),
10785 => conv_std_logic_vector(5, 8),
10786 => conv_std_logic_vector(5, 8),
10787 => conv_std_logic_vector(5, 8),
10788 => conv_std_logic_vector(5, 8),
10789 => conv_std_logic_vector(6, 8),
10790 => conv_std_logic_vector(6, 8),
10791 => conv_std_logic_vector(6, 8),
10792 => conv_std_logic_vector(6, 8),
10793 => conv_std_logic_vector(6, 8),
10794 => conv_std_logic_vector(6, 8),
10795 => conv_std_logic_vector(7, 8),
10796 => conv_std_logic_vector(7, 8),
10797 => conv_std_logic_vector(7, 8),
10798 => conv_std_logic_vector(7, 8),
10799 => conv_std_logic_vector(7, 8),
10800 => conv_std_logic_vector(7, 8),
10801 => conv_std_logic_vector(8, 8),
10802 => conv_std_logic_vector(8, 8),
10803 => conv_std_logic_vector(8, 8),
10804 => conv_std_logic_vector(8, 8),
10805 => conv_std_logic_vector(8, 8),
10806 => conv_std_logic_vector(8, 8),
10807 => conv_std_logic_vector(9, 8),
10808 => conv_std_logic_vector(9, 8),
10809 => conv_std_logic_vector(9, 8),
10810 => conv_std_logic_vector(9, 8),
10811 => conv_std_logic_vector(9, 8),
10812 => conv_std_logic_vector(9, 8),
10813 => conv_std_logic_vector(10, 8),
10814 => conv_std_logic_vector(10, 8),
10815 => conv_std_logic_vector(10, 8),
10816 => conv_std_logic_vector(10, 8),
10817 => conv_std_logic_vector(10, 8),
10818 => conv_std_logic_vector(10, 8),
10819 => conv_std_logic_vector(10, 8),
10820 => conv_std_logic_vector(11, 8),
10821 => conv_std_logic_vector(11, 8),
10822 => conv_std_logic_vector(11, 8),
10823 => conv_std_logic_vector(11, 8),
10824 => conv_std_logic_vector(11, 8),
10825 => conv_std_logic_vector(11, 8),
10826 => conv_std_logic_vector(12, 8),
10827 => conv_std_logic_vector(12, 8),
10828 => conv_std_logic_vector(12, 8),
10829 => conv_std_logic_vector(12, 8),
10830 => conv_std_logic_vector(12, 8),
10831 => conv_std_logic_vector(12, 8),
10832 => conv_std_logic_vector(13, 8),
10833 => conv_std_logic_vector(13, 8),
10834 => conv_std_logic_vector(13, 8),
10835 => conv_std_logic_vector(13, 8),
10836 => conv_std_logic_vector(13, 8),
10837 => conv_std_logic_vector(13, 8),
10838 => conv_std_logic_vector(14, 8),
10839 => conv_std_logic_vector(14, 8),
10840 => conv_std_logic_vector(14, 8),
10841 => conv_std_logic_vector(14, 8),
10842 => conv_std_logic_vector(14, 8),
10843 => conv_std_logic_vector(14, 8),
10844 => conv_std_logic_vector(15, 8),
10845 => conv_std_logic_vector(15, 8),
10846 => conv_std_logic_vector(15, 8),
10847 => conv_std_logic_vector(15, 8),
10848 => conv_std_logic_vector(15, 8),
10849 => conv_std_logic_vector(15, 8),
10850 => conv_std_logic_vector(16, 8),
10851 => conv_std_logic_vector(16, 8),
10852 => conv_std_logic_vector(16, 8),
10853 => conv_std_logic_vector(16, 8),
10854 => conv_std_logic_vector(16, 8),
10855 => conv_std_logic_vector(16, 8),
10856 => conv_std_logic_vector(17, 8),
10857 => conv_std_logic_vector(17, 8),
10858 => conv_std_logic_vector(17, 8),
10859 => conv_std_logic_vector(17, 8),
10860 => conv_std_logic_vector(17, 8),
10861 => conv_std_logic_vector(17, 8),
10862 => conv_std_logic_vector(18, 8),
10863 => conv_std_logic_vector(18, 8),
10864 => conv_std_logic_vector(18, 8),
10865 => conv_std_logic_vector(18, 8),
10866 => conv_std_logic_vector(18, 8),
10867 => conv_std_logic_vector(18, 8),
10868 => conv_std_logic_vector(19, 8),
10869 => conv_std_logic_vector(19, 8),
10870 => conv_std_logic_vector(19, 8),
10871 => conv_std_logic_vector(19, 8),
10872 => conv_std_logic_vector(19, 8),
10873 => conv_std_logic_vector(19, 8),
10874 => conv_std_logic_vector(20, 8),
10875 => conv_std_logic_vector(20, 8),
10876 => conv_std_logic_vector(20, 8),
10877 => conv_std_logic_vector(20, 8),
10878 => conv_std_logic_vector(20, 8),
10879 => conv_std_logic_vector(20, 8),
10880 => conv_std_logic_vector(21, 8),
10881 => conv_std_logic_vector(21, 8),
10882 => conv_std_logic_vector(21, 8),
10883 => conv_std_logic_vector(21, 8),
10884 => conv_std_logic_vector(21, 8),
10885 => conv_std_logic_vector(21, 8),
10886 => conv_std_logic_vector(21, 8),
10887 => conv_std_logic_vector(22, 8),
10888 => conv_std_logic_vector(22, 8),
10889 => conv_std_logic_vector(22, 8),
10890 => conv_std_logic_vector(22, 8),
10891 => conv_std_logic_vector(22, 8),
10892 => conv_std_logic_vector(22, 8),
10893 => conv_std_logic_vector(23, 8),
10894 => conv_std_logic_vector(23, 8),
10895 => conv_std_logic_vector(23, 8),
10896 => conv_std_logic_vector(23, 8),
10897 => conv_std_logic_vector(23, 8),
10898 => conv_std_logic_vector(23, 8),
10899 => conv_std_logic_vector(24, 8),
10900 => conv_std_logic_vector(24, 8),
10901 => conv_std_logic_vector(24, 8),
10902 => conv_std_logic_vector(24, 8),
10903 => conv_std_logic_vector(24, 8),
10904 => conv_std_logic_vector(24, 8),
10905 => conv_std_logic_vector(25, 8),
10906 => conv_std_logic_vector(25, 8),
10907 => conv_std_logic_vector(25, 8),
10908 => conv_std_logic_vector(25, 8),
10909 => conv_std_logic_vector(25, 8),
10910 => conv_std_logic_vector(25, 8),
10911 => conv_std_logic_vector(26, 8),
10912 => conv_std_logic_vector(26, 8),
10913 => conv_std_logic_vector(26, 8),
10914 => conv_std_logic_vector(26, 8),
10915 => conv_std_logic_vector(26, 8),
10916 => conv_std_logic_vector(26, 8),
10917 => conv_std_logic_vector(27, 8),
10918 => conv_std_logic_vector(27, 8),
10919 => conv_std_logic_vector(27, 8),
10920 => conv_std_logic_vector(27, 8),
10921 => conv_std_logic_vector(27, 8),
10922 => conv_std_logic_vector(27, 8),
10923 => conv_std_logic_vector(28, 8),
10924 => conv_std_logic_vector(28, 8),
10925 => conv_std_logic_vector(28, 8),
10926 => conv_std_logic_vector(28, 8),
10927 => conv_std_logic_vector(28, 8),
10928 => conv_std_logic_vector(28, 8),
10929 => conv_std_logic_vector(29, 8),
10930 => conv_std_logic_vector(29, 8),
10931 => conv_std_logic_vector(29, 8),
10932 => conv_std_logic_vector(29, 8),
10933 => conv_std_logic_vector(29, 8),
10934 => conv_std_logic_vector(29, 8),
10935 => conv_std_logic_vector(30, 8),
10936 => conv_std_logic_vector(30, 8),
10937 => conv_std_logic_vector(30, 8),
10938 => conv_std_logic_vector(30, 8),
10939 => conv_std_logic_vector(30, 8),
10940 => conv_std_logic_vector(30, 8),
10941 => conv_std_logic_vector(31, 8),
10942 => conv_std_logic_vector(31, 8),
10943 => conv_std_logic_vector(31, 8),
10944 => conv_std_logic_vector(31, 8),
10945 => conv_std_logic_vector(31, 8),
10946 => conv_std_logic_vector(31, 8),
10947 => conv_std_logic_vector(31, 8),
10948 => conv_std_logic_vector(32, 8),
10949 => conv_std_logic_vector(32, 8),
10950 => conv_std_logic_vector(32, 8),
10951 => conv_std_logic_vector(32, 8),
10952 => conv_std_logic_vector(32, 8),
10953 => conv_std_logic_vector(32, 8),
10954 => conv_std_logic_vector(33, 8),
10955 => conv_std_logic_vector(33, 8),
10956 => conv_std_logic_vector(33, 8),
10957 => conv_std_logic_vector(33, 8),
10958 => conv_std_logic_vector(33, 8),
10959 => conv_std_logic_vector(33, 8),
10960 => conv_std_logic_vector(34, 8),
10961 => conv_std_logic_vector(34, 8),
10962 => conv_std_logic_vector(34, 8),
10963 => conv_std_logic_vector(34, 8),
10964 => conv_std_logic_vector(34, 8),
10965 => conv_std_logic_vector(34, 8),
10966 => conv_std_logic_vector(35, 8),
10967 => conv_std_logic_vector(35, 8),
10968 => conv_std_logic_vector(35, 8),
10969 => conv_std_logic_vector(35, 8),
10970 => conv_std_logic_vector(35, 8),
10971 => conv_std_logic_vector(35, 8),
10972 => conv_std_logic_vector(36, 8),
10973 => conv_std_logic_vector(36, 8),
10974 => conv_std_logic_vector(36, 8),
10975 => conv_std_logic_vector(36, 8),
10976 => conv_std_logic_vector(36, 8),
10977 => conv_std_logic_vector(36, 8),
10978 => conv_std_logic_vector(37, 8),
10979 => conv_std_logic_vector(37, 8),
10980 => conv_std_logic_vector(37, 8),
10981 => conv_std_logic_vector(37, 8),
10982 => conv_std_logic_vector(37, 8),
10983 => conv_std_logic_vector(37, 8),
10984 => conv_std_logic_vector(38, 8),
10985 => conv_std_logic_vector(38, 8),
10986 => conv_std_logic_vector(38, 8),
10987 => conv_std_logic_vector(38, 8),
10988 => conv_std_logic_vector(38, 8),
10989 => conv_std_logic_vector(38, 8),
10990 => conv_std_logic_vector(39, 8),
10991 => conv_std_logic_vector(39, 8),
10992 => conv_std_logic_vector(39, 8),
10993 => conv_std_logic_vector(39, 8),
10994 => conv_std_logic_vector(39, 8),
10995 => conv_std_logic_vector(39, 8),
10996 => conv_std_logic_vector(40, 8),
10997 => conv_std_logic_vector(40, 8),
10998 => conv_std_logic_vector(40, 8),
10999 => conv_std_logic_vector(40, 8),
11000 => conv_std_logic_vector(40, 8),
11001 => conv_std_logic_vector(40, 8),
11002 => conv_std_logic_vector(41, 8),
11003 => conv_std_logic_vector(41, 8),
11004 => conv_std_logic_vector(41, 8),
11005 => conv_std_logic_vector(41, 8),
11006 => conv_std_logic_vector(41, 8),
11007 => conv_std_logic_vector(41, 8),
11008 => conv_std_logic_vector(0, 8),
11009 => conv_std_logic_vector(0, 8),
11010 => conv_std_logic_vector(0, 8),
11011 => conv_std_logic_vector(0, 8),
11012 => conv_std_logic_vector(0, 8),
11013 => conv_std_logic_vector(0, 8),
11014 => conv_std_logic_vector(1, 8),
11015 => conv_std_logic_vector(1, 8),
11016 => conv_std_logic_vector(1, 8),
11017 => conv_std_logic_vector(1, 8),
11018 => conv_std_logic_vector(1, 8),
11019 => conv_std_logic_vector(1, 8),
11020 => conv_std_logic_vector(2, 8),
11021 => conv_std_logic_vector(2, 8),
11022 => conv_std_logic_vector(2, 8),
11023 => conv_std_logic_vector(2, 8),
11024 => conv_std_logic_vector(2, 8),
11025 => conv_std_logic_vector(2, 8),
11026 => conv_std_logic_vector(3, 8),
11027 => conv_std_logic_vector(3, 8),
11028 => conv_std_logic_vector(3, 8),
11029 => conv_std_logic_vector(3, 8),
11030 => conv_std_logic_vector(3, 8),
11031 => conv_std_logic_vector(3, 8),
11032 => conv_std_logic_vector(4, 8),
11033 => conv_std_logic_vector(4, 8),
11034 => conv_std_logic_vector(4, 8),
11035 => conv_std_logic_vector(4, 8),
11036 => conv_std_logic_vector(4, 8),
11037 => conv_std_logic_vector(4, 8),
11038 => conv_std_logic_vector(5, 8),
11039 => conv_std_logic_vector(5, 8),
11040 => conv_std_logic_vector(5, 8),
11041 => conv_std_logic_vector(5, 8),
11042 => conv_std_logic_vector(5, 8),
11043 => conv_std_logic_vector(5, 8),
11044 => conv_std_logic_vector(6, 8),
11045 => conv_std_logic_vector(6, 8),
11046 => conv_std_logic_vector(6, 8),
11047 => conv_std_logic_vector(6, 8),
11048 => conv_std_logic_vector(6, 8),
11049 => conv_std_logic_vector(6, 8),
11050 => conv_std_logic_vector(7, 8),
11051 => conv_std_logic_vector(7, 8),
11052 => conv_std_logic_vector(7, 8),
11053 => conv_std_logic_vector(7, 8),
11054 => conv_std_logic_vector(7, 8),
11055 => conv_std_logic_vector(7, 8),
11056 => conv_std_logic_vector(8, 8),
11057 => conv_std_logic_vector(8, 8),
11058 => conv_std_logic_vector(8, 8),
11059 => conv_std_logic_vector(8, 8),
11060 => conv_std_logic_vector(8, 8),
11061 => conv_std_logic_vector(8, 8),
11062 => conv_std_logic_vector(9, 8),
11063 => conv_std_logic_vector(9, 8),
11064 => conv_std_logic_vector(9, 8),
11065 => conv_std_logic_vector(9, 8),
11066 => conv_std_logic_vector(9, 8),
11067 => conv_std_logic_vector(9, 8),
11068 => conv_std_logic_vector(10, 8),
11069 => conv_std_logic_vector(10, 8),
11070 => conv_std_logic_vector(10, 8),
11071 => conv_std_logic_vector(10, 8),
11072 => conv_std_logic_vector(10, 8),
11073 => conv_std_logic_vector(10, 8),
11074 => conv_std_logic_vector(11, 8),
11075 => conv_std_logic_vector(11, 8),
11076 => conv_std_logic_vector(11, 8),
11077 => conv_std_logic_vector(11, 8),
11078 => conv_std_logic_vector(11, 8),
11079 => conv_std_logic_vector(11, 8),
11080 => conv_std_logic_vector(12, 8),
11081 => conv_std_logic_vector(12, 8),
11082 => conv_std_logic_vector(12, 8),
11083 => conv_std_logic_vector(12, 8),
11084 => conv_std_logic_vector(12, 8),
11085 => conv_std_logic_vector(12, 8),
11086 => conv_std_logic_vector(13, 8),
11087 => conv_std_logic_vector(13, 8),
11088 => conv_std_logic_vector(13, 8),
11089 => conv_std_logic_vector(13, 8),
11090 => conv_std_logic_vector(13, 8),
11091 => conv_std_logic_vector(13, 8),
11092 => conv_std_logic_vector(14, 8),
11093 => conv_std_logic_vector(14, 8),
11094 => conv_std_logic_vector(14, 8),
11095 => conv_std_logic_vector(14, 8),
11096 => conv_std_logic_vector(14, 8),
11097 => conv_std_logic_vector(14, 8),
11098 => conv_std_logic_vector(15, 8),
11099 => conv_std_logic_vector(15, 8),
11100 => conv_std_logic_vector(15, 8),
11101 => conv_std_logic_vector(15, 8),
11102 => conv_std_logic_vector(15, 8),
11103 => conv_std_logic_vector(15, 8),
11104 => conv_std_logic_vector(16, 8),
11105 => conv_std_logic_vector(16, 8),
11106 => conv_std_logic_vector(16, 8),
11107 => conv_std_logic_vector(16, 8),
11108 => conv_std_logic_vector(16, 8),
11109 => conv_std_logic_vector(16, 8),
11110 => conv_std_logic_vector(17, 8),
11111 => conv_std_logic_vector(17, 8),
11112 => conv_std_logic_vector(17, 8),
11113 => conv_std_logic_vector(17, 8),
11114 => conv_std_logic_vector(17, 8),
11115 => conv_std_logic_vector(17, 8),
11116 => conv_std_logic_vector(18, 8),
11117 => conv_std_logic_vector(18, 8),
11118 => conv_std_logic_vector(18, 8),
11119 => conv_std_logic_vector(18, 8),
11120 => conv_std_logic_vector(18, 8),
11121 => conv_std_logic_vector(18, 8),
11122 => conv_std_logic_vector(19, 8),
11123 => conv_std_logic_vector(19, 8),
11124 => conv_std_logic_vector(19, 8),
11125 => conv_std_logic_vector(19, 8),
11126 => conv_std_logic_vector(19, 8),
11127 => conv_std_logic_vector(19, 8),
11128 => conv_std_logic_vector(20, 8),
11129 => conv_std_logic_vector(20, 8),
11130 => conv_std_logic_vector(20, 8),
11131 => conv_std_logic_vector(20, 8),
11132 => conv_std_logic_vector(20, 8),
11133 => conv_std_logic_vector(20, 8),
11134 => conv_std_logic_vector(21, 8),
11135 => conv_std_logic_vector(21, 8),
11136 => conv_std_logic_vector(21, 8),
11137 => conv_std_logic_vector(21, 8),
11138 => conv_std_logic_vector(21, 8),
11139 => conv_std_logic_vector(22, 8),
11140 => conv_std_logic_vector(22, 8),
11141 => conv_std_logic_vector(22, 8),
11142 => conv_std_logic_vector(22, 8),
11143 => conv_std_logic_vector(22, 8),
11144 => conv_std_logic_vector(22, 8),
11145 => conv_std_logic_vector(23, 8),
11146 => conv_std_logic_vector(23, 8),
11147 => conv_std_logic_vector(23, 8),
11148 => conv_std_logic_vector(23, 8),
11149 => conv_std_logic_vector(23, 8),
11150 => conv_std_logic_vector(23, 8),
11151 => conv_std_logic_vector(24, 8),
11152 => conv_std_logic_vector(24, 8),
11153 => conv_std_logic_vector(24, 8),
11154 => conv_std_logic_vector(24, 8),
11155 => conv_std_logic_vector(24, 8),
11156 => conv_std_logic_vector(24, 8),
11157 => conv_std_logic_vector(25, 8),
11158 => conv_std_logic_vector(25, 8),
11159 => conv_std_logic_vector(25, 8),
11160 => conv_std_logic_vector(25, 8),
11161 => conv_std_logic_vector(25, 8),
11162 => conv_std_logic_vector(25, 8),
11163 => conv_std_logic_vector(26, 8),
11164 => conv_std_logic_vector(26, 8),
11165 => conv_std_logic_vector(26, 8),
11166 => conv_std_logic_vector(26, 8),
11167 => conv_std_logic_vector(26, 8),
11168 => conv_std_logic_vector(26, 8),
11169 => conv_std_logic_vector(27, 8),
11170 => conv_std_logic_vector(27, 8),
11171 => conv_std_logic_vector(27, 8),
11172 => conv_std_logic_vector(27, 8),
11173 => conv_std_logic_vector(27, 8),
11174 => conv_std_logic_vector(27, 8),
11175 => conv_std_logic_vector(28, 8),
11176 => conv_std_logic_vector(28, 8),
11177 => conv_std_logic_vector(28, 8),
11178 => conv_std_logic_vector(28, 8),
11179 => conv_std_logic_vector(28, 8),
11180 => conv_std_logic_vector(28, 8),
11181 => conv_std_logic_vector(29, 8),
11182 => conv_std_logic_vector(29, 8),
11183 => conv_std_logic_vector(29, 8),
11184 => conv_std_logic_vector(29, 8),
11185 => conv_std_logic_vector(29, 8),
11186 => conv_std_logic_vector(29, 8),
11187 => conv_std_logic_vector(30, 8),
11188 => conv_std_logic_vector(30, 8),
11189 => conv_std_logic_vector(30, 8),
11190 => conv_std_logic_vector(30, 8),
11191 => conv_std_logic_vector(30, 8),
11192 => conv_std_logic_vector(30, 8),
11193 => conv_std_logic_vector(31, 8),
11194 => conv_std_logic_vector(31, 8),
11195 => conv_std_logic_vector(31, 8),
11196 => conv_std_logic_vector(31, 8),
11197 => conv_std_logic_vector(31, 8),
11198 => conv_std_logic_vector(31, 8),
11199 => conv_std_logic_vector(32, 8),
11200 => conv_std_logic_vector(32, 8),
11201 => conv_std_logic_vector(32, 8),
11202 => conv_std_logic_vector(32, 8),
11203 => conv_std_logic_vector(32, 8),
11204 => conv_std_logic_vector(32, 8),
11205 => conv_std_logic_vector(33, 8),
11206 => conv_std_logic_vector(33, 8),
11207 => conv_std_logic_vector(33, 8),
11208 => conv_std_logic_vector(33, 8),
11209 => conv_std_logic_vector(33, 8),
11210 => conv_std_logic_vector(33, 8),
11211 => conv_std_logic_vector(34, 8),
11212 => conv_std_logic_vector(34, 8),
11213 => conv_std_logic_vector(34, 8),
11214 => conv_std_logic_vector(34, 8),
11215 => conv_std_logic_vector(34, 8),
11216 => conv_std_logic_vector(34, 8),
11217 => conv_std_logic_vector(35, 8),
11218 => conv_std_logic_vector(35, 8),
11219 => conv_std_logic_vector(35, 8),
11220 => conv_std_logic_vector(35, 8),
11221 => conv_std_logic_vector(35, 8),
11222 => conv_std_logic_vector(35, 8),
11223 => conv_std_logic_vector(36, 8),
11224 => conv_std_logic_vector(36, 8),
11225 => conv_std_logic_vector(36, 8),
11226 => conv_std_logic_vector(36, 8),
11227 => conv_std_logic_vector(36, 8),
11228 => conv_std_logic_vector(36, 8),
11229 => conv_std_logic_vector(37, 8),
11230 => conv_std_logic_vector(37, 8),
11231 => conv_std_logic_vector(37, 8),
11232 => conv_std_logic_vector(37, 8),
11233 => conv_std_logic_vector(37, 8),
11234 => conv_std_logic_vector(37, 8),
11235 => conv_std_logic_vector(38, 8),
11236 => conv_std_logic_vector(38, 8),
11237 => conv_std_logic_vector(38, 8),
11238 => conv_std_logic_vector(38, 8),
11239 => conv_std_logic_vector(38, 8),
11240 => conv_std_logic_vector(38, 8),
11241 => conv_std_logic_vector(39, 8),
11242 => conv_std_logic_vector(39, 8),
11243 => conv_std_logic_vector(39, 8),
11244 => conv_std_logic_vector(39, 8),
11245 => conv_std_logic_vector(39, 8),
11246 => conv_std_logic_vector(39, 8),
11247 => conv_std_logic_vector(40, 8),
11248 => conv_std_logic_vector(40, 8),
11249 => conv_std_logic_vector(40, 8),
11250 => conv_std_logic_vector(40, 8),
11251 => conv_std_logic_vector(40, 8),
11252 => conv_std_logic_vector(40, 8),
11253 => conv_std_logic_vector(41, 8),
11254 => conv_std_logic_vector(41, 8),
11255 => conv_std_logic_vector(41, 8),
11256 => conv_std_logic_vector(41, 8),
11257 => conv_std_logic_vector(41, 8),
11258 => conv_std_logic_vector(41, 8),
11259 => conv_std_logic_vector(42, 8),
11260 => conv_std_logic_vector(42, 8),
11261 => conv_std_logic_vector(42, 8),
11262 => conv_std_logic_vector(42, 8),
11263 => conv_std_logic_vector(42, 8),
11264 => conv_std_logic_vector(0, 8),
11265 => conv_std_logic_vector(0, 8),
11266 => conv_std_logic_vector(0, 8),
11267 => conv_std_logic_vector(0, 8),
11268 => conv_std_logic_vector(0, 8),
11269 => conv_std_logic_vector(0, 8),
11270 => conv_std_logic_vector(1, 8),
11271 => conv_std_logic_vector(1, 8),
11272 => conv_std_logic_vector(1, 8),
11273 => conv_std_logic_vector(1, 8),
11274 => conv_std_logic_vector(1, 8),
11275 => conv_std_logic_vector(1, 8),
11276 => conv_std_logic_vector(2, 8),
11277 => conv_std_logic_vector(2, 8),
11278 => conv_std_logic_vector(2, 8),
11279 => conv_std_logic_vector(2, 8),
11280 => conv_std_logic_vector(2, 8),
11281 => conv_std_logic_vector(2, 8),
11282 => conv_std_logic_vector(3, 8),
11283 => conv_std_logic_vector(3, 8),
11284 => conv_std_logic_vector(3, 8),
11285 => conv_std_logic_vector(3, 8),
11286 => conv_std_logic_vector(3, 8),
11287 => conv_std_logic_vector(3, 8),
11288 => conv_std_logic_vector(4, 8),
11289 => conv_std_logic_vector(4, 8),
11290 => conv_std_logic_vector(4, 8),
11291 => conv_std_logic_vector(4, 8),
11292 => conv_std_logic_vector(4, 8),
11293 => conv_std_logic_vector(4, 8),
11294 => conv_std_logic_vector(5, 8),
11295 => conv_std_logic_vector(5, 8),
11296 => conv_std_logic_vector(5, 8),
11297 => conv_std_logic_vector(5, 8),
11298 => conv_std_logic_vector(5, 8),
11299 => conv_std_logic_vector(6, 8),
11300 => conv_std_logic_vector(6, 8),
11301 => conv_std_logic_vector(6, 8),
11302 => conv_std_logic_vector(6, 8),
11303 => conv_std_logic_vector(6, 8),
11304 => conv_std_logic_vector(6, 8),
11305 => conv_std_logic_vector(7, 8),
11306 => conv_std_logic_vector(7, 8),
11307 => conv_std_logic_vector(7, 8),
11308 => conv_std_logic_vector(7, 8),
11309 => conv_std_logic_vector(7, 8),
11310 => conv_std_logic_vector(7, 8),
11311 => conv_std_logic_vector(8, 8),
11312 => conv_std_logic_vector(8, 8),
11313 => conv_std_logic_vector(8, 8),
11314 => conv_std_logic_vector(8, 8),
11315 => conv_std_logic_vector(8, 8),
11316 => conv_std_logic_vector(8, 8),
11317 => conv_std_logic_vector(9, 8),
11318 => conv_std_logic_vector(9, 8),
11319 => conv_std_logic_vector(9, 8),
11320 => conv_std_logic_vector(9, 8),
11321 => conv_std_logic_vector(9, 8),
11322 => conv_std_logic_vector(9, 8),
11323 => conv_std_logic_vector(10, 8),
11324 => conv_std_logic_vector(10, 8),
11325 => conv_std_logic_vector(10, 8),
11326 => conv_std_logic_vector(10, 8),
11327 => conv_std_logic_vector(10, 8),
11328 => conv_std_logic_vector(11, 8),
11329 => conv_std_logic_vector(11, 8),
11330 => conv_std_logic_vector(11, 8),
11331 => conv_std_logic_vector(11, 8),
11332 => conv_std_logic_vector(11, 8),
11333 => conv_std_logic_vector(11, 8),
11334 => conv_std_logic_vector(12, 8),
11335 => conv_std_logic_vector(12, 8),
11336 => conv_std_logic_vector(12, 8),
11337 => conv_std_logic_vector(12, 8),
11338 => conv_std_logic_vector(12, 8),
11339 => conv_std_logic_vector(12, 8),
11340 => conv_std_logic_vector(13, 8),
11341 => conv_std_logic_vector(13, 8),
11342 => conv_std_logic_vector(13, 8),
11343 => conv_std_logic_vector(13, 8),
11344 => conv_std_logic_vector(13, 8),
11345 => conv_std_logic_vector(13, 8),
11346 => conv_std_logic_vector(14, 8),
11347 => conv_std_logic_vector(14, 8),
11348 => conv_std_logic_vector(14, 8),
11349 => conv_std_logic_vector(14, 8),
11350 => conv_std_logic_vector(14, 8),
11351 => conv_std_logic_vector(14, 8),
11352 => conv_std_logic_vector(15, 8),
11353 => conv_std_logic_vector(15, 8),
11354 => conv_std_logic_vector(15, 8),
11355 => conv_std_logic_vector(15, 8),
11356 => conv_std_logic_vector(15, 8),
11357 => conv_std_logic_vector(15, 8),
11358 => conv_std_logic_vector(16, 8),
11359 => conv_std_logic_vector(16, 8),
11360 => conv_std_logic_vector(16, 8),
11361 => conv_std_logic_vector(16, 8),
11362 => conv_std_logic_vector(16, 8),
11363 => conv_std_logic_vector(17, 8),
11364 => conv_std_logic_vector(17, 8),
11365 => conv_std_logic_vector(17, 8),
11366 => conv_std_logic_vector(17, 8),
11367 => conv_std_logic_vector(17, 8),
11368 => conv_std_logic_vector(17, 8),
11369 => conv_std_logic_vector(18, 8),
11370 => conv_std_logic_vector(18, 8),
11371 => conv_std_logic_vector(18, 8),
11372 => conv_std_logic_vector(18, 8),
11373 => conv_std_logic_vector(18, 8),
11374 => conv_std_logic_vector(18, 8),
11375 => conv_std_logic_vector(19, 8),
11376 => conv_std_logic_vector(19, 8),
11377 => conv_std_logic_vector(19, 8),
11378 => conv_std_logic_vector(19, 8),
11379 => conv_std_logic_vector(19, 8),
11380 => conv_std_logic_vector(19, 8),
11381 => conv_std_logic_vector(20, 8),
11382 => conv_std_logic_vector(20, 8),
11383 => conv_std_logic_vector(20, 8),
11384 => conv_std_logic_vector(20, 8),
11385 => conv_std_logic_vector(20, 8),
11386 => conv_std_logic_vector(20, 8),
11387 => conv_std_logic_vector(21, 8),
11388 => conv_std_logic_vector(21, 8),
11389 => conv_std_logic_vector(21, 8),
11390 => conv_std_logic_vector(21, 8),
11391 => conv_std_logic_vector(21, 8),
11392 => conv_std_logic_vector(22, 8),
11393 => conv_std_logic_vector(22, 8),
11394 => conv_std_logic_vector(22, 8),
11395 => conv_std_logic_vector(22, 8),
11396 => conv_std_logic_vector(22, 8),
11397 => conv_std_logic_vector(22, 8),
11398 => conv_std_logic_vector(23, 8),
11399 => conv_std_logic_vector(23, 8),
11400 => conv_std_logic_vector(23, 8),
11401 => conv_std_logic_vector(23, 8),
11402 => conv_std_logic_vector(23, 8),
11403 => conv_std_logic_vector(23, 8),
11404 => conv_std_logic_vector(24, 8),
11405 => conv_std_logic_vector(24, 8),
11406 => conv_std_logic_vector(24, 8),
11407 => conv_std_logic_vector(24, 8),
11408 => conv_std_logic_vector(24, 8),
11409 => conv_std_logic_vector(24, 8),
11410 => conv_std_logic_vector(25, 8),
11411 => conv_std_logic_vector(25, 8),
11412 => conv_std_logic_vector(25, 8),
11413 => conv_std_logic_vector(25, 8),
11414 => conv_std_logic_vector(25, 8),
11415 => conv_std_logic_vector(25, 8),
11416 => conv_std_logic_vector(26, 8),
11417 => conv_std_logic_vector(26, 8),
11418 => conv_std_logic_vector(26, 8),
11419 => conv_std_logic_vector(26, 8),
11420 => conv_std_logic_vector(26, 8),
11421 => conv_std_logic_vector(26, 8),
11422 => conv_std_logic_vector(27, 8),
11423 => conv_std_logic_vector(27, 8),
11424 => conv_std_logic_vector(27, 8),
11425 => conv_std_logic_vector(27, 8),
11426 => conv_std_logic_vector(27, 8),
11427 => conv_std_logic_vector(28, 8),
11428 => conv_std_logic_vector(28, 8),
11429 => conv_std_logic_vector(28, 8),
11430 => conv_std_logic_vector(28, 8),
11431 => conv_std_logic_vector(28, 8),
11432 => conv_std_logic_vector(28, 8),
11433 => conv_std_logic_vector(29, 8),
11434 => conv_std_logic_vector(29, 8),
11435 => conv_std_logic_vector(29, 8),
11436 => conv_std_logic_vector(29, 8),
11437 => conv_std_logic_vector(29, 8),
11438 => conv_std_logic_vector(29, 8),
11439 => conv_std_logic_vector(30, 8),
11440 => conv_std_logic_vector(30, 8),
11441 => conv_std_logic_vector(30, 8),
11442 => conv_std_logic_vector(30, 8),
11443 => conv_std_logic_vector(30, 8),
11444 => conv_std_logic_vector(30, 8),
11445 => conv_std_logic_vector(31, 8),
11446 => conv_std_logic_vector(31, 8),
11447 => conv_std_logic_vector(31, 8),
11448 => conv_std_logic_vector(31, 8),
11449 => conv_std_logic_vector(31, 8),
11450 => conv_std_logic_vector(31, 8),
11451 => conv_std_logic_vector(32, 8),
11452 => conv_std_logic_vector(32, 8),
11453 => conv_std_logic_vector(32, 8),
11454 => conv_std_logic_vector(32, 8),
11455 => conv_std_logic_vector(32, 8),
11456 => conv_std_logic_vector(33, 8),
11457 => conv_std_logic_vector(33, 8),
11458 => conv_std_logic_vector(33, 8),
11459 => conv_std_logic_vector(33, 8),
11460 => conv_std_logic_vector(33, 8),
11461 => conv_std_logic_vector(33, 8),
11462 => conv_std_logic_vector(34, 8),
11463 => conv_std_logic_vector(34, 8),
11464 => conv_std_logic_vector(34, 8),
11465 => conv_std_logic_vector(34, 8),
11466 => conv_std_logic_vector(34, 8),
11467 => conv_std_logic_vector(34, 8),
11468 => conv_std_logic_vector(35, 8),
11469 => conv_std_logic_vector(35, 8),
11470 => conv_std_logic_vector(35, 8),
11471 => conv_std_logic_vector(35, 8),
11472 => conv_std_logic_vector(35, 8),
11473 => conv_std_logic_vector(35, 8),
11474 => conv_std_logic_vector(36, 8),
11475 => conv_std_logic_vector(36, 8),
11476 => conv_std_logic_vector(36, 8),
11477 => conv_std_logic_vector(36, 8),
11478 => conv_std_logic_vector(36, 8),
11479 => conv_std_logic_vector(36, 8),
11480 => conv_std_logic_vector(37, 8),
11481 => conv_std_logic_vector(37, 8),
11482 => conv_std_logic_vector(37, 8),
11483 => conv_std_logic_vector(37, 8),
11484 => conv_std_logic_vector(37, 8),
11485 => conv_std_logic_vector(37, 8),
11486 => conv_std_logic_vector(38, 8),
11487 => conv_std_logic_vector(38, 8),
11488 => conv_std_logic_vector(38, 8),
11489 => conv_std_logic_vector(38, 8),
11490 => conv_std_logic_vector(38, 8),
11491 => conv_std_logic_vector(39, 8),
11492 => conv_std_logic_vector(39, 8),
11493 => conv_std_logic_vector(39, 8),
11494 => conv_std_logic_vector(39, 8),
11495 => conv_std_logic_vector(39, 8),
11496 => conv_std_logic_vector(39, 8),
11497 => conv_std_logic_vector(40, 8),
11498 => conv_std_logic_vector(40, 8),
11499 => conv_std_logic_vector(40, 8),
11500 => conv_std_logic_vector(40, 8),
11501 => conv_std_logic_vector(40, 8),
11502 => conv_std_logic_vector(40, 8),
11503 => conv_std_logic_vector(41, 8),
11504 => conv_std_logic_vector(41, 8),
11505 => conv_std_logic_vector(41, 8),
11506 => conv_std_logic_vector(41, 8),
11507 => conv_std_logic_vector(41, 8),
11508 => conv_std_logic_vector(41, 8),
11509 => conv_std_logic_vector(42, 8),
11510 => conv_std_logic_vector(42, 8),
11511 => conv_std_logic_vector(42, 8),
11512 => conv_std_logic_vector(42, 8),
11513 => conv_std_logic_vector(42, 8),
11514 => conv_std_logic_vector(42, 8),
11515 => conv_std_logic_vector(43, 8),
11516 => conv_std_logic_vector(43, 8),
11517 => conv_std_logic_vector(43, 8),
11518 => conv_std_logic_vector(43, 8),
11519 => conv_std_logic_vector(43, 8),
11520 => conv_std_logic_vector(0, 8),
11521 => conv_std_logic_vector(0, 8),
11522 => conv_std_logic_vector(0, 8),
11523 => conv_std_logic_vector(0, 8),
11524 => conv_std_logic_vector(0, 8),
11525 => conv_std_logic_vector(0, 8),
11526 => conv_std_logic_vector(1, 8),
11527 => conv_std_logic_vector(1, 8),
11528 => conv_std_logic_vector(1, 8),
11529 => conv_std_logic_vector(1, 8),
11530 => conv_std_logic_vector(1, 8),
11531 => conv_std_logic_vector(1, 8),
11532 => conv_std_logic_vector(2, 8),
11533 => conv_std_logic_vector(2, 8),
11534 => conv_std_logic_vector(2, 8),
11535 => conv_std_logic_vector(2, 8),
11536 => conv_std_logic_vector(2, 8),
11537 => conv_std_logic_vector(2, 8),
11538 => conv_std_logic_vector(3, 8),
11539 => conv_std_logic_vector(3, 8),
11540 => conv_std_logic_vector(3, 8),
11541 => conv_std_logic_vector(3, 8),
11542 => conv_std_logic_vector(3, 8),
11543 => conv_std_logic_vector(4, 8),
11544 => conv_std_logic_vector(4, 8),
11545 => conv_std_logic_vector(4, 8),
11546 => conv_std_logic_vector(4, 8),
11547 => conv_std_logic_vector(4, 8),
11548 => conv_std_logic_vector(4, 8),
11549 => conv_std_logic_vector(5, 8),
11550 => conv_std_logic_vector(5, 8),
11551 => conv_std_logic_vector(5, 8),
11552 => conv_std_logic_vector(5, 8),
11553 => conv_std_logic_vector(5, 8),
11554 => conv_std_logic_vector(5, 8),
11555 => conv_std_logic_vector(6, 8),
11556 => conv_std_logic_vector(6, 8),
11557 => conv_std_logic_vector(6, 8),
11558 => conv_std_logic_vector(6, 8),
11559 => conv_std_logic_vector(6, 8),
11560 => conv_std_logic_vector(7, 8),
11561 => conv_std_logic_vector(7, 8),
11562 => conv_std_logic_vector(7, 8),
11563 => conv_std_logic_vector(7, 8),
11564 => conv_std_logic_vector(7, 8),
11565 => conv_std_logic_vector(7, 8),
11566 => conv_std_logic_vector(8, 8),
11567 => conv_std_logic_vector(8, 8),
11568 => conv_std_logic_vector(8, 8),
11569 => conv_std_logic_vector(8, 8),
11570 => conv_std_logic_vector(8, 8),
11571 => conv_std_logic_vector(8, 8),
11572 => conv_std_logic_vector(9, 8),
11573 => conv_std_logic_vector(9, 8),
11574 => conv_std_logic_vector(9, 8),
11575 => conv_std_logic_vector(9, 8),
11576 => conv_std_logic_vector(9, 8),
11577 => conv_std_logic_vector(10, 8),
11578 => conv_std_logic_vector(10, 8),
11579 => conv_std_logic_vector(10, 8),
11580 => conv_std_logic_vector(10, 8),
11581 => conv_std_logic_vector(10, 8),
11582 => conv_std_logic_vector(10, 8),
11583 => conv_std_logic_vector(11, 8),
11584 => conv_std_logic_vector(11, 8),
11585 => conv_std_logic_vector(11, 8),
11586 => conv_std_logic_vector(11, 8),
11587 => conv_std_logic_vector(11, 8),
11588 => conv_std_logic_vector(11, 8),
11589 => conv_std_logic_vector(12, 8),
11590 => conv_std_logic_vector(12, 8),
11591 => conv_std_logic_vector(12, 8),
11592 => conv_std_logic_vector(12, 8),
11593 => conv_std_logic_vector(12, 8),
11594 => conv_std_logic_vector(13, 8),
11595 => conv_std_logic_vector(13, 8),
11596 => conv_std_logic_vector(13, 8),
11597 => conv_std_logic_vector(13, 8),
11598 => conv_std_logic_vector(13, 8),
11599 => conv_std_logic_vector(13, 8),
11600 => conv_std_logic_vector(14, 8),
11601 => conv_std_logic_vector(14, 8),
11602 => conv_std_logic_vector(14, 8),
11603 => conv_std_logic_vector(14, 8),
11604 => conv_std_logic_vector(14, 8),
11605 => conv_std_logic_vector(14, 8),
11606 => conv_std_logic_vector(15, 8),
11607 => conv_std_logic_vector(15, 8),
11608 => conv_std_logic_vector(15, 8),
11609 => conv_std_logic_vector(15, 8),
11610 => conv_std_logic_vector(15, 8),
11611 => conv_std_logic_vector(15, 8),
11612 => conv_std_logic_vector(16, 8),
11613 => conv_std_logic_vector(16, 8),
11614 => conv_std_logic_vector(16, 8),
11615 => conv_std_logic_vector(16, 8),
11616 => conv_std_logic_vector(16, 8),
11617 => conv_std_logic_vector(17, 8),
11618 => conv_std_logic_vector(17, 8),
11619 => conv_std_logic_vector(17, 8),
11620 => conv_std_logic_vector(17, 8),
11621 => conv_std_logic_vector(17, 8),
11622 => conv_std_logic_vector(17, 8),
11623 => conv_std_logic_vector(18, 8),
11624 => conv_std_logic_vector(18, 8),
11625 => conv_std_logic_vector(18, 8),
11626 => conv_std_logic_vector(18, 8),
11627 => conv_std_logic_vector(18, 8),
11628 => conv_std_logic_vector(18, 8),
11629 => conv_std_logic_vector(19, 8),
11630 => conv_std_logic_vector(19, 8),
11631 => conv_std_logic_vector(19, 8),
11632 => conv_std_logic_vector(19, 8),
11633 => conv_std_logic_vector(19, 8),
11634 => conv_std_logic_vector(20, 8),
11635 => conv_std_logic_vector(20, 8),
11636 => conv_std_logic_vector(20, 8),
11637 => conv_std_logic_vector(20, 8),
11638 => conv_std_logic_vector(20, 8),
11639 => conv_std_logic_vector(20, 8),
11640 => conv_std_logic_vector(21, 8),
11641 => conv_std_logic_vector(21, 8),
11642 => conv_std_logic_vector(21, 8),
11643 => conv_std_logic_vector(21, 8),
11644 => conv_std_logic_vector(21, 8),
11645 => conv_std_logic_vector(21, 8),
11646 => conv_std_logic_vector(22, 8),
11647 => conv_std_logic_vector(22, 8),
11648 => conv_std_logic_vector(22, 8),
11649 => conv_std_logic_vector(22, 8),
11650 => conv_std_logic_vector(22, 8),
11651 => conv_std_logic_vector(23, 8),
11652 => conv_std_logic_vector(23, 8),
11653 => conv_std_logic_vector(23, 8),
11654 => conv_std_logic_vector(23, 8),
11655 => conv_std_logic_vector(23, 8),
11656 => conv_std_logic_vector(23, 8),
11657 => conv_std_logic_vector(24, 8),
11658 => conv_std_logic_vector(24, 8),
11659 => conv_std_logic_vector(24, 8),
11660 => conv_std_logic_vector(24, 8),
11661 => conv_std_logic_vector(24, 8),
11662 => conv_std_logic_vector(24, 8),
11663 => conv_std_logic_vector(25, 8),
11664 => conv_std_logic_vector(25, 8),
11665 => conv_std_logic_vector(25, 8),
11666 => conv_std_logic_vector(25, 8),
11667 => conv_std_logic_vector(25, 8),
11668 => conv_std_logic_vector(26, 8),
11669 => conv_std_logic_vector(26, 8),
11670 => conv_std_logic_vector(26, 8),
11671 => conv_std_logic_vector(26, 8),
11672 => conv_std_logic_vector(26, 8),
11673 => conv_std_logic_vector(26, 8),
11674 => conv_std_logic_vector(27, 8),
11675 => conv_std_logic_vector(27, 8),
11676 => conv_std_logic_vector(27, 8),
11677 => conv_std_logic_vector(27, 8),
11678 => conv_std_logic_vector(27, 8),
11679 => conv_std_logic_vector(27, 8),
11680 => conv_std_logic_vector(28, 8),
11681 => conv_std_logic_vector(28, 8),
11682 => conv_std_logic_vector(28, 8),
11683 => conv_std_logic_vector(28, 8),
11684 => conv_std_logic_vector(28, 8),
11685 => conv_std_logic_vector(29, 8),
11686 => conv_std_logic_vector(29, 8),
11687 => conv_std_logic_vector(29, 8),
11688 => conv_std_logic_vector(29, 8),
11689 => conv_std_logic_vector(29, 8),
11690 => conv_std_logic_vector(29, 8),
11691 => conv_std_logic_vector(30, 8),
11692 => conv_std_logic_vector(30, 8),
11693 => conv_std_logic_vector(30, 8),
11694 => conv_std_logic_vector(30, 8),
11695 => conv_std_logic_vector(30, 8),
11696 => conv_std_logic_vector(30, 8),
11697 => conv_std_logic_vector(31, 8),
11698 => conv_std_logic_vector(31, 8),
11699 => conv_std_logic_vector(31, 8),
11700 => conv_std_logic_vector(31, 8),
11701 => conv_std_logic_vector(31, 8),
11702 => conv_std_logic_vector(31, 8),
11703 => conv_std_logic_vector(32, 8),
11704 => conv_std_logic_vector(32, 8),
11705 => conv_std_logic_vector(32, 8),
11706 => conv_std_logic_vector(32, 8),
11707 => conv_std_logic_vector(32, 8),
11708 => conv_std_logic_vector(33, 8),
11709 => conv_std_logic_vector(33, 8),
11710 => conv_std_logic_vector(33, 8),
11711 => conv_std_logic_vector(33, 8),
11712 => conv_std_logic_vector(33, 8),
11713 => conv_std_logic_vector(33, 8),
11714 => conv_std_logic_vector(34, 8),
11715 => conv_std_logic_vector(34, 8),
11716 => conv_std_logic_vector(34, 8),
11717 => conv_std_logic_vector(34, 8),
11718 => conv_std_logic_vector(34, 8),
11719 => conv_std_logic_vector(34, 8),
11720 => conv_std_logic_vector(35, 8),
11721 => conv_std_logic_vector(35, 8),
11722 => conv_std_logic_vector(35, 8),
11723 => conv_std_logic_vector(35, 8),
11724 => conv_std_logic_vector(35, 8),
11725 => conv_std_logic_vector(36, 8),
11726 => conv_std_logic_vector(36, 8),
11727 => conv_std_logic_vector(36, 8),
11728 => conv_std_logic_vector(36, 8),
11729 => conv_std_logic_vector(36, 8),
11730 => conv_std_logic_vector(36, 8),
11731 => conv_std_logic_vector(37, 8),
11732 => conv_std_logic_vector(37, 8),
11733 => conv_std_logic_vector(37, 8),
11734 => conv_std_logic_vector(37, 8),
11735 => conv_std_logic_vector(37, 8),
11736 => conv_std_logic_vector(37, 8),
11737 => conv_std_logic_vector(38, 8),
11738 => conv_std_logic_vector(38, 8),
11739 => conv_std_logic_vector(38, 8),
11740 => conv_std_logic_vector(38, 8),
11741 => conv_std_logic_vector(38, 8),
11742 => conv_std_logic_vector(39, 8),
11743 => conv_std_logic_vector(39, 8),
11744 => conv_std_logic_vector(39, 8),
11745 => conv_std_logic_vector(39, 8),
11746 => conv_std_logic_vector(39, 8),
11747 => conv_std_logic_vector(39, 8),
11748 => conv_std_logic_vector(40, 8),
11749 => conv_std_logic_vector(40, 8),
11750 => conv_std_logic_vector(40, 8),
11751 => conv_std_logic_vector(40, 8),
11752 => conv_std_logic_vector(40, 8),
11753 => conv_std_logic_vector(40, 8),
11754 => conv_std_logic_vector(41, 8),
11755 => conv_std_logic_vector(41, 8),
11756 => conv_std_logic_vector(41, 8),
11757 => conv_std_logic_vector(41, 8),
11758 => conv_std_logic_vector(41, 8),
11759 => conv_std_logic_vector(42, 8),
11760 => conv_std_logic_vector(42, 8),
11761 => conv_std_logic_vector(42, 8),
11762 => conv_std_logic_vector(42, 8),
11763 => conv_std_logic_vector(42, 8),
11764 => conv_std_logic_vector(42, 8),
11765 => conv_std_logic_vector(43, 8),
11766 => conv_std_logic_vector(43, 8),
11767 => conv_std_logic_vector(43, 8),
11768 => conv_std_logic_vector(43, 8),
11769 => conv_std_logic_vector(43, 8),
11770 => conv_std_logic_vector(43, 8),
11771 => conv_std_logic_vector(44, 8),
11772 => conv_std_logic_vector(44, 8),
11773 => conv_std_logic_vector(44, 8),
11774 => conv_std_logic_vector(44, 8),
11775 => conv_std_logic_vector(44, 8),
11776 => conv_std_logic_vector(0, 8),
11777 => conv_std_logic_vector(0, 8),
11778 => conv_std_logic_vector(0, 8),
11779 => conv_std_logic_vector(0, 8),
11780 => conv_std_logic_vector(0, 8),
11781 => conv_std_logic_vector(0, 8),
11782 => conv_std_logic_vector(1, 8),
11783 => conv_std_logic_vector(1, 8),
11784 => conv_std_logic_vector(1, 8),
11785 => conv_std_logic_vector(1, 8),
11786 => conv_std_logic_vector(1, 8),
11787 => conv_std_logic_vector(1, 8),
11788 => conv_std_logic_vector(2, 8),
11789 => conv_std_logic_vector(2, 8),
11790 => conv_std_logic_vector(2, 8),
11791 => conv_std_logic_vector(2, 8),
11792 => conv_std_logic_vector(2, 8),
11793 => conv_std_logic_vector(3, 8),
11794 => conv_std_logic_vector(3, 8),
11795 => conv_std_logic_vector(3, 8),
11796 => conv_std_logic_vector(3, 8),
11797 => conv_std_logic_vector(3, 8),
11798 => conv_std_logic_vector(3, 8),
11799 => conv_std_logic_vector(4, 8),
11800 => conv_std_logic_vector(4, 8),
11801 => conv_std_logic_vector(4, 8),
11802 => conv_std_logic_vector(4, 8),
11803 => conv_std_logic_vector(4, 8),
11804 => conv_std_logic_vector(5, 8),
11805 => conv_std_logic_vector(5, 8),
11806 => conv_std_logic_vector(5, 8),
11807 => conv_std_logic_vector(5, 8),
11808 => conv_std_logic_vector(5, 8),
11809 => conv_std_logic_vector(5, 8),
11810 => conv_std_logic_vector(6, 8),
11811 => conv_std_logic_vector(6, 8),
11812 => conv_std_logic_vector(6, 8),
11813 => conv_std_logic_vector(6, 8),
11814 => conv_std_logic_vector(6, 8),
11815 => conv_std_logic_vector(7, 8),
11816 => conv_std_logic_vector(7, 8),
11817 => conv_std_logic_vector(7, 8),
11818 => conv_std_logic_vector(7, 8),
11819 => conv_std_logic_vector(7, 8),
11820 => conv_std_logic_vector(7, 8),
11821 => conv_std_logic_vector(8, 8),
11822 => conv_std_logic_vector(8, 8),
11823 => conv_std_logic_vector(8, 8),
11824 => conv_std_logic_vector(8, 8),
11825 => conv_std_logic_vector(8, 8),
11826 => conv_std_logic_vector(8, 8),
11827 => conv_std_logic_vector(9, 8),
11828 => conv_std_logic_vector(9, 8),
11829 => conv_std_logic_vector(9, 8),
11830 => conv_std_logic_vector(9, 8),
11831 => conv_std_logic_vector(9, 8),
11832 => conv_std_logic_vector(10, 8),
11833 => conv_std_logic_vector(10, 8),
11834 => conv_std_logic_vector(10, 8),
11835 => conv_std_logic_vector(10, 8),
11836 => conv_std_logic_vector(10, 8),
11837 => conv_std_logic_vector(10, 8),
11838 => conv_std_logic_vector(11, 8),
11839 => conv_std_logic_vector(11, 8),
11840 => conv_std_logic_vector(11, 8),
11841 => conv_std_logic_vector(11, 8),
11842 => conv_std_logic_vector(11, 8),
11843 => conv_std_logic_vector(12, 8),
11844 => conv_std_logic_vector(12, 8),
11845 => conv_std_logic_vector(12, 8),
11846 => conv_std_logic_vector(12, 8),
11847 => conv_std_logic_vector(12, 8),
11848 => conv_std_logic_vector(12, 8),
11849 => conv_std_logic_vector(13, 8),
11850 => conv_std_logic_vector(13, 8),
11851 => conv_std_logic_vector(13, 8),
11852 => conv_std_logic_vector(13, 8),
11853 => conv_std_logic_vector(13, 8),
11854 => conv_std_logic_vector(14, 8),
11855 => conv_std_logic_vector(14, 8),
11856 => conv_std_logic_vector(14, 8),
11857 => conv_std_logic_vector(14, 8),
11858 => conv_std_logic_vector(14, 8),
11859 => conv_std_logic_vector(14, 8),
11860 => conv_std_logic_vector(15, 8),
11861 => conv_std_logic_vector(15, 8),
11862 => conv_std_logic_vector(15, 8),
11863 => conv_std_logic_vector(15, 8),
11864 => conv_std_logic_vector(15, 8),
11865 => conv_std_logic_vector(15, 8),
11866 => conv_std_logic_vector(16, 8),
11867 => conv_std_logic_vector(16, 8),
11868 => conv_std_logic_vector(16, 8),
11869 => conv_std_logic_vector(16, 8),
11870 => conv_std_logic_vector(16, 8),
11871 => conv_std_logic_vector(17, 8),
11872 => conv_std_logic_vector(17, 8),
11873 => conv_std_logic_vector(17, 8),
11874 => conv_std_logic_vector(17, 8),
11875 => conv_std_logic_vector(17, 8),
11876 => conv_std_logic_vector(17, 8),
11877 => conv_std_logic_vector(18, 8),
11878 => conv_std_logic_vector(18, 8),
11879 => conv_std_logic_vector(18, 8),
11880 => conv_std_logic_vector(18, 8),
11881 => conv_std_logic_vector(18, 8),
11882 => conv_std_logic_vector(19, 8),
11883 => conv_std_logic_vector(19, 8),
11884 => conv_std_logic_vector(19, 8),
11885 => conv_std_logic_vector(19, 8),
11886 => conv_std_logic_vector(19, 8),
11887 => conv_std_logic_vector(19, 8),
11888 => conv_std_logic_vector(20, 8),
11889 => conv_std_logic_vector(20, 8),
11890 => conv_std_logic_vector(20, 8),
11891 => conv_std_logic_vector(20, 8),
11892 => conv_std_logic_vector(20, 8),
11893 => conv_std_logic_vector(21, 8),
11894 => conv_std_logic_vector(21, 8),
11895 => conv_std_logic_vector(21, 8),
11896 => conv_std_logic_vector(21, 8),
11897 => conv_std_logic_vector(21, 8),
11898 => conv_std_logic_vector(21, 8),
11899 => conv_std_logic_vector(22, 8),
11900 => conv_std_logic_vector(22, 8),
11901 => conv_std_logic_vector(22, 8),
11902 => conv_std_logic_vector(22, 8),
11903 => conv_std_logic_vector(22, 8),
11904 => conv_std_logic_vector(23, 8),
11905 => conv_std_logic_vector(23, 8),
11906 => conv_std_logic_vector(23, 8),
11907 => conv_std_logic_vector(23, 8),
11908 => conv_std_logic_vector(23, 8),
11909 => conv_std_logic_vector(23, 8),
11910 => conv_std_logic_vector(24, 8),
11911 => conv_std_logic_vector(24, 8),
11912 => conv_std_logic_vector(24, 8),
11913 => conv_std_logic_vector(24, 8),
11914 => conv_std_logic_vector(24, 8),
11915 => conv_std_logic_vector(24, 8),
11916 => conv_std_logic_vector(25, 8),
11917 => conv_std_logic_vector(25, 8),
11918 => conv_std_logic_vector(25, 8),
11919 => conv_std_logic_vector(25, 8),
11920 => conv_std_logic_vector(25, 8),
11921 => conv_std_logic_vector(26, 8),
11922 => conv_std_logic_vector(26, 8),
11923 => conv_std_logic_vector(26, 8),
11924 => conv_std_logic_vector(26, 8),
11925 => conv_std_logic_vector(26, 8),
11926 => conv_std_logic_vector(26, 8),
11927 => conv_std_logic_vector(27, 8),
11928 => conv_std_logic_vector(27, 8),
11929 => conv_std_logic_vector(27, 8),
11930 => conv_std_logic_vector(27, 8),
11931 => conv_std_logic_vector(27, 8),
11932 => conv_std_logic_vector(28, 8),
11933 => conv_std_logic_vector(28, 8),
11934 => conv_std_logic_vector(28, 8),
11935 => conv_std_logic_vector(28, 8),
11936 => conv_std_logic_vector(28, 8),
11937 => conv_std_logic_vector(28, 8),
11938 => conv_std_logic_vector(29, 8),
11939 => conv_std_logic_vector(29, 8),
11940 => conv_std_logic_vector(29, 8),
11941 => conv_std_logic_vector(29, 8),
11942 => conv_std_logic_vector(29, 8),
11943 => conv_std_logic_vector(30, 8),
11944 => conv_std_logic_vector(30, 8),
11945 => conv_std_logic_vector(30, 8),
11946 => conv_std_logic_vector(30, 8),
11947 => conv_std_logic_vector(30, 8),
11948 => conv_std_logic_vector(30, 8),
11949 => conv_std_logic_vector(31, 8),
11950 => conv_std_logic_vector(31, 8),
11951 => conv_std_logic_vector(31, 8),
11952 => conv_std_logic_vector(31, 8),
11953 => conv_std_logic_vector(31, 8),
11954 => conv_std_logic_vector(31, 8),
11955 => conv_std_logic_vector(32, 8),
11956 => conv_std_logic_vector(32, 8),
11957 => conv_std_logic_vector(32, 8),
11958 => conv_std_logic_vector(32, 8),
11959 => conv_std_logic_vector(32, 8),
11960 => conv_std_logic_vector(33, 8),
11961 => conv_std_logic_vector(33, 8),
11962 => conv_std_logic_vector(33, 8),
11963 => conv_std_logic_vector(33, 8),
11964 => conv_std_logic_vector(33, 8),
11965 => conv_std_logic_vector(33, 8),
11966 => conv_std_logic_vector(34, 8),
11967 => conv_std_logic_vector(34, 8),
11968 => conv_std_logic_vector(34, 8),
11969 => conv_std_logic_vector(34, 8),
11970 => conv_std_logic_vector(34, 8),
11971 => conv_std_logic_vector(35, 8),
11972 => conv_std_logic_vector(35, 8),
11973 => conv_std_logic_vector(35, 8),
11974 => conv_std_logic_vector(35, 8),
11975 => conv_std_logic_vector(35, 8),
11976 => conv_std_logic_vector(35, 8),
11977 => conv_std_logic_vector(36, 8),
11978 => conv_std_logic_vector(36, 8),
11979 => conv_std_logic_vector(36, 8),
11980 => conv_std_logic_vector(36, 8),
11981 => conv_std_logic_vector(36, 8),
11982 => conv_std_logic_vector(37, 8),
11983 => conv_std_logic_vector(37, 8),
11984 => conv_std_logic_vector(37, 8),
11985 => conv_std_logic_vector(37, 8),
11986 => conv_std_logic_vector(37, 8),
11987 => conv_std_logic_vector(37, 8),
11988 => conv_std_logic_vector(38, 8),
11989 => conv_std_logic_vector(38, 8),
11990 => conv_std_logic_vector(38, 8),
11991 => conv_std_logic_vector(38, 8),
11992 => conv_std_logic_vector(38, 8),
11993 => conv_std_logic_vector(38, 8),
11994 => conv_std_logic_vector(39, 8),
11995 => conv_std_logic_vector(39, 8),
11996 => conv_std_logic_vector(39, 8),
11997 => conv_std_logic_vector(39, 8),
11998 => conv_std_logic_vector(39, 8),
11999 => conv_std_logic_vector(40, 8),
12000 => conv_std_logic_vector(40, 8),
12001 => conv_std_logic_vector(40, 8),
12002 => conv_std_logic_vector(40, 8),
12003 => conv_std_logic_vector(40, 8),
12004 => conv_std_logic_vector(40, 8),
12005 => conv_std_logic_vector(41, 8),
12006 => conv_std_logic_vector(41, 8),
12007 => conv_std_logic_vector(41, 8),
12008 => conv_std_logic_vector(41, 8),
12009 => conv_std_logic_vector(41, 8),
12010 => conv_std_logic_vector(42, 8),
12011 => conv_std_logic_vector(42, 8),
12012 => conv_std_logic_vector(42, 8),
12013 => conv_std_logic_vector(42, 8),
12014 => conv_std_logic_vector(42, 8),
12015 => conv_std_logic_vector(42, 8),
12016 => conv_std_logic_vector(43, 8),
12017 => conv_std_logic_vector(43, 8),
12018 => conv_std_logic_vector(43, 8),
12019 => conv_std_logic_vector(43, 8),
12020 => conv_std_logic_vector(43, 8),
12021 => conv_std_logic_vector(44, 8),
12022 => conv_std_logic_vector(44, 8),
12023 => conv_std_logic_vector(44, 8),
12024 => conv_std_logic_vector(44, 8),
12025 => conv_std_logic_vector(44, 8),
12026 => conv_std_logic_vector(44, 8),
12027 => conv_std_logic_vector(45, 8),
12028 => conv_std_logic_vector(45, 8),
12029 => conv_std_logic_vector(45, 8),
12030 => conv_std_logic_vector(45, 8),
12031 => conv_std_logic_vector(45, 8),
12032 => conv_std_logic_vector(0, 8),
12033 => conv_std_logic_vector(0, 8),
12034 => conv_std_logic_vector(0, 8),
12035 => conv_std_logic_vector(0, 8),
12036 => conv_std_logic_vector(0, 8),
12037 => conv_std_logic_vector(0, 8),
12038 => conv_std_logic_vector(1, 8),
12039 => conv_std_logic_vector(1, 8),
12040 => conv_std_logic_vector(1, 8),
12041 => conv_std_logic_vector(1, 8),
12042 => conv_std_logic_vector(1, 8),
12043 => conv_std_logic_vector(2, 8),
12044 => conv_std_logic_vector(2, 8),
12045 => conv_std_logic_vector(2, 8),
12046 => conv_std_logic_vector(2, 8),
12047 => conv_std_logic_vector(2, 8),
12048 => conv_std_logic_vector(2, 8),
12049 => conv_std_logic_vector(3, 8),
12050 => conv_std_logic_vector(3, 8),
12051 => conv_std_logic_vector(3, 8),
12052 => conv_std_logic_vector(3, 8),
12053 => conv_std_logic_vector(3, 8),
12054 => conv_std_logic_vector(4, 8),
12055 => conv_std_logic_vector(4, 8),
12056 => conv_std_logic_vector(4, 8),
12057 => conv_std_logic_vector(4, 8),
12058 => conv_std_logic_vector(4, 8),
12059 => conv_std_logic_vector(4, 8),
12060 => conv_std_logic_vector(5, 8),
12061 => conv_std_logic_vector(5, 8),
12062 => conv_std_logic_vector(5, 8),
12063 => conv_std_logic_vector(5, 8),
12064 => conv_std_logic_vector(5, 8),
12065 => conv_std_logic_vector(6, 8),
12066 => conv_std_logic_vector(6, 8),
12067 => conv_std_logic_vector(6, 8),
12068 => conv_std_logic_vector(6, 8),
12069 => conv_std_logic_vector(6, 8),
12070 => conv_std_logic_vector(6, 8),
12071 => conv_std_logic_vector(7, 8),
12072 => conv_std_logic_vector(7, 8),
12073 => conv_std_logic_vector(7, 8),
12074 => conv_std_logic_vector(7, 8),
12075 => conv_std_logic_vector(7, 8),
12076 => conv_std_logic_vector(8, 8),
12077 => conv_std_logic_vector(8, 8),
12078 => conv_std_logic_vector(8, 8),
12079 => conv_std_logic_vector(8, 8),
12080 => conv_std_logic_vector(8, 8),
12081 => conv_std_logic_vector(8, 8),
12082 => conv_std_logic_vector(9, 8),
12083 => conv_std_logic_vector(9, 8),
12084 => conv_std_logic_vector(9, 8),
12085 => conv_std_logic_vector(9, 8),
12086 => conv_std_logic_vector(9, 8),
12087 => conv_std_logic_vector(10, 8),
12088 => conv_std_logic_vector(10, 8),
12089 => conv_std_logic_vector(10, 8),
12090 => conv_std_logic_vector(10, 8),
12091 => conv_std_logic_vector(10, 8),
12092 => conv_std_logic_vector(11, 8),
12093 => conv_std_logic_vector(11, 8),
12094 => conv_std_logic_vector(11, 8),
12095 => conv_std_logic_vector(11, 8),
12096 => conv_std_logic_vector(11, 8),
12097 => conv_std_logic_vector(11, 8),
12098 => conv_std_logic_vector(12, 8),
12099 => conv_std_logic_vector(12, 8),
12100 => conv_std_logic_vector(12, 8),
12101 => conv_std_logic_vector(12, 8),
12102 => conv_std_logic_vector(12, 8),
12103 => conv_std_logic_vector(13, 8),
12104 => conv_std_logic_vector(13, 8),
12105 => conv_std_logic_vector(13, 8),
12106 => conv_std_logic_vector(13, 8),
12107 => conv_std_logic_vector(13, 8),
12108 => conv_std_logic_vector(13, 8),
12109 => conv_std_logic_vector(14, 8),
12110 => conv_std_logic_vector(14, 8),
12111 => conv_std_logic_vector(14, 8),
12112 => conv_std_logic_vector(14, 8),
12113 => conv_std_logic_vector(14, 8),
12114 => conv_std_logic_vector(15, 8),
12115 => conv_std_logic_vector(15, 8),
12116 => conv_std_logic_vector(15, 8),
12117 => conv_std_logic_vector(15, 8),
12118 => conv_std_logic_vector(15, 8),
12119 => conv_std_logic_vector(15, 8),
12120 => conv_std_logic_vector(16, 8),
12121 => conv_std_logic_vector(16, 8),
12122 => conv_std_logic_vector(16, 8),
12123 => conv_std_logic_vector(16, 8),
12124 => conv_std_logic_vector(16, 8),
12125 => conv_std_logic_vector(17, 8),
12126 => conv_std_logic_vector(17, 8),
12127 => conv_std_logic_vector(17, 8),
12128 => conv_std_logic_vector(17, 8),
12129 => conv_std_logic_vector(17, 8),
12130 => conv_std_logic_vector(17, 8),
12131 => conv_std_logic_vector(18, 8),
12132 => conv_std_logic_vector(18, 8),
12133 => conv_std_logic_vector(18, 8),
12134 => conv_std_logic_vector(18, 8),
12135 => conv_std_logic_vector(18, 8),
12136 => conv_std_logic_vector(19, 8),
12137 => conv_std_logic_vector(19, 8),
12138 => conv_std_logic_vector(19, 8),
12139 => conv_std_logic_vector(19, 8),
12140 => conv_std_logic_vector(19, 8),
12141 => conv_std_logic_vector(20, 8),
12142 => conv_std_logic_vector(20, 8),
12143 => conv_std_logic_vector(20, 8),
12144 => conv_std_logic_vector(20, 8),
12145 => conv_std_logic_vector(20, 8),
12146 => conv_std_logic_vector(20, 8),
12147 => conv_std_logic_vector(21, 8),
12148 => conv_std_logic_vector(21, 8),
12149 => conv_std_logic_vector(21, 8),
12150 => conv_std_logic_vector(21, 8),
12151 => conv_std_logic_vector(21, 8),
12152 => conv_std_logic_vector(22, 8),
12153 => conv_std_logic_vector(22, 8),
12154 => conv_std_logic_vector(22, 8),
12155 => conv_std_logic_vector(22, 8),
12156 => conv_std_logic_vector(22, 8),
12157 => conv_std_logic_vector(22, 8),
12158 => conv_std_logic_vector(23, 8),
12159 => conv_std_logic_vector(23, 8),
12160 => conv_std_logic_vector(23, 8),
12161 => conv_std_logic_vector(23, 8),
12162 => conv_std_logic_vector(23, 8),
12163 => conv_std_logic_vector(24, 8),
12164 => conv_std_logic_vector(24, 8),
12165 => conv_std_logic_vector(24, 8),
12166 => conv_std_logic_vector(24, 8),
12167 => conv_std_logic_vector(24, 8),
12168 => conv_std_logic_vector(24, 8),
12169 => conv_std_logic_vector(25, 8),
12170 => conv_std_logic_vector(25, 8),
12171 => conv_std_logic_vector(25, 8),
12172 => conv_std_logic_vector(25, 8),
12173 => conv_std_logic_vector(25, 8),
12174 => conv_std_logic_vector(26, 8),
12175 => conv_std_logic_vector(26, 8),
12176 => conv_std_logic_vector(26, 8),
12177 => conv_std_logic_vector(26, 8),
12178 => conv_std_logic_vector(26, 8),
12179 => conv_std_logic_vector(26, 8),
12180 => conv_std_logic_vector(27, 8),
12181 => conv_std_logic_vector(27, 8),
12182 => conv_std_logic_vector(27, 8),
12183 => conv_std_logic_vector(27, 8),
12184 => conv_std_logic_vector(27, 8),
12185 => conv_std_logic_vector(28, 8),
12186 => conv_std_logic_vector(28, 8),
12187 => conv_std_logic_vector(28, 8),
12188 => conv_std_logic_vector(28, 8),
12189 => conv_std_logic_vector(28, 8),
12190 => conv_std_logic_vector(29, 8),
12191 => conv_std_logic_vector(29, 8),
12192 => conv_std_logic_vector(29, 8),
12193 => conv_std_logic_vector(29, 8),
12194 => conv_std_logic_vector(29, 8),
12195 => conv_std_logic_vector(29, 8),
12196 => conv_std_logic_vector(30, 8),
12197 => conv_std_logic_vector(30, 8),
12198 => conv_std_logic_vector(30, 8),
12199 => conv_std_logic_vector(30, 8),
12200 => conv_std_logic_vector(30, 8),
12201 => conv_std_logic_vector(31, 8),
12202 => conv_std_logic_vector(31, 8),
12203 => conv_std_logic_vector(31, 8),
12204 => conv_std_logic_vector(31, 8),
12205 => conv_std_logic_vector(31, 8),
12206 => conv_std_logic_vector(31, 8),
12207 => conv_std_logic_vector(32, 8),
12208 => conv_std_logic_vector(32, 8),
12209 => conv_std_logic_vector(32, 8),
12210 => conv_std_logic_vector(32, 8),
12211 => conv_std_logic_vector(32, 8),
12212 => conv_std_logic_vector(33, 8),
12213 => conv_std_logic_vector(33, 8),
12214 => conv_std_logic_vector(33, 8),
12215 => conv_std_logic_vector(33, 8),
12216 => conv_std_logic_vector(33, 8),
12217 => conv_std_logic_vector(33, 8),
12218 => conv_std_logic_vector(34, 8),
12219 => conv_std_logic_vector(34, 8),
12220 => conv_std_logic_vector(34, 8),
12221 => conv_std_logic_vector(34, 8),
12222 => conv_std_logic_vector(34, 8),
12223 => conv_std_logic_vector(35, 8),
12224 => conv_std_logic_vector(35, 8),
12225 => conv_std_logic_vector(35, 8),
12226 => conv_std_logic_vector(35, 8),
12227 => conv_std_logic_vector(35, 8),
12228 => conv_std_logic_vector(35, 8),
12229 => conv_std_logic_vector(36, 8),
12230 => conv_std_logic_vector(36, 8),
12231 => conv_std_logic_vector(36, 8),
12232 => conv_std_logic_vector(36, 8),
12233 => conv_std_logic_vector(36, 8),
12234 => conv_std_logic_vector(37, 8),
12235 => conv_std_logic_vector(37, 8),
12236 => conv_std_logic_vector(37, 8),
12237 => conv_std_logic_vector(37, 8),
12238 => conv_std_logic_vector(37, 8),
12239 => conv_std_logic_vector(38, 8),
12240 => conv_std_logic_vector(38, 8),
12241 => conv_std_logic_vector(38, 8),
12242 => conv_std_logic_vector(38, 8),
12243 => conv_std_logic_vector(38, 8),
12244 => conv_std_logic_vector(38, 8),
12245 => conv_std_logic_vector(39, 8),
12246 => conv_std_logic_vector(39, 8),
12247 => conv_std_logic_vector(39, 8),
12248 => conv_std_logic_vector(39, 8),
12249 => conv_std_logic_vector(39, 8),
12250 => conv_std_logic_vector(40, 8),
12251 => conv_std_logic_vector(40, 8),
12252 => conv_std_logic_vector(40, 8),
12253 => conv_std_logic_vector(40, 8),
12254 => conv_std_logic_vector(40, 8),
12255 => conv_std_logic_vector(40, 8),
12256 => conv_std_logic_vector(41, 8),
12257 => conv_std_logic_vector(41, 8),
12258 => conv_std_logic_vector(41, 8),
12259 => conv_std_logic_vector(41, 8),
12260 => conv_std_logic_vector(41, 8),
12261 => conv_std_logic_vector(42, 8),
12262 => conv_std_logic_vector(42, 8),
12263 => conv_std_logic_vector(42, 8),
12264 => conv_std_logic_vector(42, 8),
12265 => conv_std_logic_vector(42, 8),
12266 => conv_std_logic_vector(42, 8),
12267 => conv_std_logic_vector(43, 8),
12268 => conv_std_logic_vector(43, 8),
12269 => conv_std_logic_vector(43, 8),
12270 => conv_std_logic_vector(43, 8),
12271 => conv_std_logic_vector(43, 8),
12272 => conv_std_logic_vector(44, 8),
12273 => conv_std_logic_vector(44, 8),
12274 => conv_std_logic_vector(44, 8),
12275 => conv_std_logic_vector(44, 8),
12276 => conv_std_logic_vector(44, 8),
12277 => conv_std_logic_vector(44, 8),
12278 => conv_std_logic_vector(45, 8),
12279 => conv_std_logic_vector(45, 8),
12280 => conv_std_logic_vector(45, 8),
12281 => conv_std_logic_vector(45, 8),
12282 => conv_std_logic_vector(45, 8),
12283 => conv_std_logic_vector(46, 8),
12284 => conv_std_logic_vector(46, 8),
12285 => conv_std_logic_vector(46, 8),
12286 => conv_std_logic_vector(46, 8),
12287 => conv_std_logic_vector(46, 8),
12288 => conv_std_logic_vector(0, 8),
12289 => conv_std_logic_vector(0, 8),
12290 => conv_std_logic_vector(0, 8),
12291 => conv_std_logic_vector(0, 8),
12292 => conv_std_logic_vector(0, 8),
12293 => conv_std_logic_vector(0, 8),
12294 => conv_std_logic_vector(1, 8),
12295 => conv_std_logic_vector(1, 8),
12296 => conv_std_logic_vector(1, 8),
12297 => conv_std_logic_vector(1, 8),
12298 => conv_std_logic_vector(1, 8),
12299 => conv_std_logic_vector(2, 8),
12300 => conv_std_logic_vector(2, 8),
12301 => conv_std_logic_vector(2, 8),
12302 => conv_std_logic_vector(2, 8),
12303 => conv_std_logic_vector(2, 8),
12304 => conv_std_logic_vector(3, 8),
12305 => conv_std_logic_vector(3, 8),
12306 => conv_std_logic_vector(3, 8),
12307 => conv_std_logic_vector(3, 8),
12308 => conv_std_logic_vector(3, 8),
12309 => conv_std_logic_vector(3, 8),
12310 => conv_std_logic_vector(4, 8),
12311 => conv_std_logic_vector(4, 8),
12312 => conv_std_logic_vector(4, 8),
12313 => conv_std_logic_vector(4, 8),
12314 => conv_std_logic_vector(4, 8),
12315 => conv_std_logic_vector(5, 8),
12316 => conv_std_logic_vector(5, 8),
12317 => conv_std_logic_vector(5, 8),
12318 => conv_std_logic_vector(5, 8),
12319 => conv_std_logic_vector(5, 8),
12320 => conv_std_logic_vector(6, 8),
12321 => conv_std_logic_vector(6, 8),
12322 => conv_std_logic_vector(6, 8),
12323 => conv_std_logic_vector(6, 8),
12324 => conv_std_logic_vector(6, 8),
12325 => conv_std_logic_vector(6, 8),
12326 => conv_std_logic_vector(7, 8),
12327 => conv_std_logic_vector(7, 8),
12328 => conv_std_logic_vector(7, 8),
12329 => conv_std_logic_vector(7, 8),
12330 => conv_std_logic_vector(7, 8),
12331 => conv_std_logic_vector(8, 8),
12332 => conv_std_logic_vector(8, 8),
12333 => conv_std_logic_vector(8, 8),
12334 => conv_std_logic_vector(8, 8),
12335 => conv_std_logic_vector(8, 8),
12336 => conv_std_logic_vector(9, 8),
12337 => conv_std_logic_vector(9, 8),
12338 => conv_std_logic_vector(9, 8),
12339 => conv_std_logic_vector(9, 8),
12340 => conv_std_logic_vector(9, 8),
12341 => conv_std_logic_vector(9, 8),
12342 => conv_std_logic_vector(10, 8),
12343 => conv_std_logic_vector(10, 8),
12344 => conv_std_logic_vector(10, 8),
12345 => conv_std_logic_vector(10, 8),
12346 => conv_std_logic_vector(10, 8),
12347 => conv_std_logic_vector(11, 8),
12348 => conv_std_logic_vector(11, 8),
12349 => conv_std_logic_vector(11, 8),
12350 => conv_std_logic_vector(11, 8),
12351 => conv_std_logic_vector(11, 8),
12352 => conv_std_logic_vector(12, 8),
12353 => conv_std_logic_vector(12, 8),
12354 => conv_std_logic_vector(12, 8),
12355 => conv_std_logic_vector(12, 8),
12356 => conv_std_logic_vector(12, 8),
12357 => conv_std_logic_vector(12, 8),
12358 => conv_std_logic_vector(13, 8),
12359 => conv_std_logic_vector(13, 8),
12360 => conv_std_logic_vector(13, 8),
12361 => conv_std_logic_vector(13, 8),
12362 => conv_std_logic_vector(13, 8),
12363 => conv_std_logic_vector(14, 8),
12364 => conv_std_logic_vector(14, 8),
12365 => conv_std_logic_vector(14, 8),
12366 => conv_std_logic_vector(14, 8),
12367 => conv_std_logic_vector(14, 8),
12368 => conv_std_logic_vector(15, 8),
12369 => conv_std_logic_vector(15, 8),
12370 => conv_std_logic_vector(15, 8),
12371 => conv_std_logic_vector(15, 8),
12372 => conv_std_logic_vector(15, 8),
12373 => conv_std_logic_vector(15, 8),
12374 => conv_std_logic_vector(16, 8),
12375 => conv_std_logic_vector(16, 8),
12376 => conv_std_logic_vector(16, 8),
12377 => conv_std_logic_vector(16, 8),
12378 => conv_std_logic_vector(16, 8),
12379 => conv_std_logic_vector(17, 8),
12380 => conv_std_logic_vector(17, 8),
12381 => conv_std_logic_vector(17, 8),
12382 => conv_std_logic_vector(17, 8),
12383 => conv_std_logic_vector(17, 8),
12384 => conv_std_logic_vector(18, 8),
12385 => conv_std_logic_vector(18, 8),
12386 => conv_std_logic_vector(18, 8),
12387 => conv_std_logic_vector(18, 8),
12388 => conv_std_logic_vector(18, 8),
12389 => conv_std_logic_vector(18, 8),
12390 => conv_std_logic_vector(19, 8),
12391 => conv_std_logic_vector(19, 8),
12392 => conv_std_logic_vector(19, 8),
12393 => conv_std_logic_vector(19, 8),
12394 => conv_std_logic_vector(19, 8),
12395 => conv_std_logic_vector(20, 8),
12396 => conv_std_logic_vector(20, 8),
12397 => conv_std_logic_vector(20, 8),
12398 => conv_std_logic_vector(20, 8),
12399 => conv_std_logic_vector(20, 8),
12400 => conv_std_logic_vector(21, 8),
12401 => conv_std_logic_vector(21, 8),
12402 => conv_std_logic_vector(21, 8),
12403 => conv_std_logic_vector(21, 8),
12404 => conv_std_logic_vector(21, 8),
12405 => conv_std_logic_vector(21, 8),
12406 => conv_std_logic_vector(22, 8),
12407 => conv_std_logic_vector(22, 8),
12408 => conv_std_logic_vector(22, 8),
12409 => conv_std_logic_vector(22, 8),
12410 => conv_std_logic_vector(22, 8),
12411 => conv_std_logic_vector(23, 8),
12412 => conv_std_logic_vector(23, 8),
12413 => conv_std_logic_vector(23, 8),
12414 => conv_std_logic_vector(23, 8),
12415 => conv_std_logic_vector(23, 8),
12416 => conv_std_logic_vector(24, 8),
12417 => conv_std_logic_vector(24, 8),
12418 => conv_std_logic_vector(24, 8),
12419 => conv_std_logic_vector(24, 8),
12420 => conv_std_logic_vector(24, 8),
12421 => conv_std_logic_vector(24, 8),
12422 => conv_std_logic_vector(25, 8),
12423 => conv_std_logic_vector(25, 8),
12424 => conv_std_logic_vector(25, 8),
12425 => conv_std_logic_vector(25, 8),
12426 => conv_std_logic_vector(25, 8),
12427 => conv_std_logic_vector(26, 8),
12428 => conv_std_logic_vector(26, 8),
12429 => conv_std_logic_vector(26, 8),
12430 => conv_std_logic_vector(26, 8),
12431 => conv_std_logic_vector(26, 8),
12432 => conv_std_logic_vector(27, 8),
12433 => conv_std_logic_vector(27, 8),
12434 => conv_std_logic_vector(27, 8),
12435 => conv_std_logic_vector(27, 8),
12436 => conv_std_logic_vector(27, 8),
12437 => conv_std_logic_vector(27, 8),
12438 => conv_std_logic_vector(28, 8),
12439 => conv_std_logic_vector(28, 8),
12440 => conv_std_logic_vector(28, 8),
12441 => conv_std_logic_vector(28, 8),
12442 => conv_std_logic_vector(28, 8),
12443 => conv_std_logic_vector(29, 8),
12444 => conv_std_logic_vector(29, 8),
12445 => conv_std_logic_vector(29, 8),
12446 => conv_std_logic_vector(29, 8),
12447 => conv_std_logic_vector(29, 8),
12448 => conv_std_logic_vector(30, 8),
12449 => conv_std_logic_vector(30, 8),
12450 => conv_std_logic_vector(30, 8),
12451 => conv_std_logic_vector(30, 8),
12452 => conv_std_logic_vector(30, 8),
12453 => conv_std_logic_vector(30, 8),
12454 => conv_std_logic_vector(31, 8),
12455 => conv_std_logic_vector(31, 8),
12456 => conv_std_logic_vector(31, 8),
12457 => conv_std_logic_vector(31, 8),
12458 => conv_std_logic_vector(31, 8),
12459 => conv_std_logic_vector(32, 8),
12460 => conv_std_logic_vector(32, 8),
12461 => conv_std_logic_vector(32, 8),
12462 => conv_std_logic_vector(32, 8),
12463 => conv_std_logic_vector(32, 8),
12464 => conv_std_logic_vector(33, 8),
12465 => conv_std_logic_vector(33, 8),
12466 => conv_std_logic_vector(33, 8),
12467 => conv_std_logic_vector(33, 8),
12468 => conv_std_logic_vector(33, 8),
12469 => conv_std_logic_vector(33, 8),
12470 => conv_std_logic_vector(34, 8),
12471 => conv_std_logic_vector(34, 8),
12472 => conv_std_logic_vector(34, 8),
12473 => conv_std_logic_vector(34, 8),
12474 => conv_std_logic_vector(34, 8),
12475 => conv_std_logic_vector(35, 8),
12476 => conv_std_logic_vector(35, 8),
12477 => conv_std_logic_vector(35, 8),
12478 => conv_std_logic_vector(35, 8),
12479 => conv_std_logic_vector(35, 8),
12480 => conv_std_logic_vector(36, 8),
12481 => conv_std_logic_vector(36, 8),
12482 => conv_std_logic_vector(36, 8),
12483 => conv_std_logic_vector(36, 8),
12484 => conv_std_logic_vector(36, 8),
12485 => conv_std_logic_vector(36, 8),
12486 => conv_std_logic_vector(37, 8),
12487 => conv_std_logic_vector(37, 8),
12488 => conv_std_logic_vector(37, 8),
12489 => conv_std_logic_vector(37, 8),
12490 => conv_std_logic_vector(37, 8),
12491 => conv_std_logic_vector(38, 8),
12492 => conv_std_logic_vector(38, 8),
12493 => conv_std_logic_vector(38, 8),
12494 => conv_std_logic_vector(38, 8),
12495 => conv_std_logic_vector(38, 8),
12496 => conv_std_logic_vector(39, 8),
12497 => conv_std_logic_vector(39, 8),
12498 => conv_std_logic_vector(39, 8),
12499 => conv_std_logic_vector(39, 8),
12500 => conv_std_logic_vector(39, 8),
12501 => conv_std_logic_vector(39, 8),
12502 => conv_std_logic_vector(40, 8),
12503 => conv_std_logic_vector(40, 8),
12504 => conv_std_logic_vector(40, 8),
12505 => conv_std_logic_vector(40, 8),
12506 => conv_std_logic_vector(40, 8),
12507 => conv_std_logic_vector(41, 8),
12508 => conv_std_logic_vector(41, 8),
12509 => conv_std_logic_vector(41, 8),
12510 => conv_std_logic_vector(41, 8),
12511 => conv_std_logic_vector(41, 8),
12512 => conv_std_logic_vector(42, 8),
12513 => conv_std_logic_vector(42, 8),
12514 => conv_std_logic_vector(42, 8),
12515 => conv_std_logic_vector(42, 8),
12516 => conv_std_logic_vector(42, 8),
12517 => conv_std_logic_vector(42, 8),
12518 => conv_std_logic_vector(43, 8),
12519 => conv_std_logic_vector(43, 8),
12520 => conv_std_logic_vector(43, 8),
12521 => conv_std_logic_vector(43, 8),
12522 => conv_std_logic_vector(43, 8),
12523 => conv_std_logic_vector(44, 8),
12524 => conv_std_logic_vector(44, 8),
12525 => conv_std_logic_vector(44, 8),
12526 => conv_std_logic_vector(44, 8),
12527 => conv_std_logic_vector(44, 8),
12528 => conv_std_logic_vector(45, 8),
12529 => conv_std_logic_vector(45, 8),
12530 => conv_std_logic_vector(45, 8),
12531 => conv_std_logic_vector(45, 8),
12532 => conv_std_logic_vector(45, 8),
12533 => conv_std_logic_vector(45, 8),
12534 => conv_std_logic_vector(46, 8),
12535 => conv_std_logic_vector(46, 8),
12536 => conv_std_logic_vector(46, 8),
12537 => conv_std_logic_vector(46, 8),
12538 => conv_std_logic_vector(46, 8),
12539 => conv_std_logic_vector(47, 8),
12540 => conv_std_logic_vector(47, 8),
12541 => conv_std_logic_vector(47, 8),
12542 => conv_std_logic_vector(47, 8),
12543 => conv_std_logic_vector(47, 8),
12544 => conv_std_logic_vector(0, 8),
12545 => conv_std_logic_vector(0, 8),
12546 => conv_std_logic_vector(0, 8),
12547 => conv_std_logic_vector(0, 8),
12548 => conv_std_logic_vector(0, 8),
12549 => conv_std_logic_vector(0, 8),
12550 => conv_std_logic_vector(1, 8),
12551 => conv_std_logic_vector(1, 8),
12552 => conv_std_logic_vector(1, 8),
12553 => conv_std_logic_vector(1, 8),
12554 => conv_std_logic_vector(1, 8),
12555 => conv_std_logic_vector(2, 8),
12556 => conv_std_logic_vector(2, 8),
12557 => conv_std_logic_vector(2, 8),
12558 => conv_std_logic_vector(2, 8),
12559 => conv_std_logic_vector(2, 8),
12560 => conv_std_logic_vector(3, 8),
12561 => conv_std_logic_vector(3, 8),
12562 => conv_std_logic_vector(3, 8),
12563 => conv_std_logic_vector(3, 8),
12564 => conv_std_logic_vector(3, 8),
12565 => conv_std_logic_vector(4, 8),
12566 => conv_std_logic_vector(4, 8),
12567 => conv_std_logic_vector(4, 8),
12568 => conv_std_logic_vector(4, 8),
12569 => conv_std_logic_vector(4, 8),
12570 => conv_std_logic_vector(4, 8),
12571 => conv_std_logic_vector(5, 8),
12572 => conv_std_logic_vector(5, 8),
12573 => conv_std_logic_vector(5, 8),
12574 => conv_std_logic_vector(5, 8),
12575 => conv_std_logic_vector(5, 8),
12576 => conv_std_logic_vector(6, 8),
12577 => conv_std_logic_vector(6, 8),
12578 => conv_std_logic_vector(6, 8),
12579 => conv_std_logic_vector(6, 8),
12580 => conv_std_logic_vector(6, 8),
12581 => conv_std_logic_vector(7, 8),
12582 => conv_std_logic_vector(7, 8),
12583 => conv_std_logic_vector(7, 8),
12584 => conv_std_logic_vector(7, 8),
12585 => conv_std_logic_vector(7, 8),
12586 => conv_std_logic_vector(8, 8),
12587 => conv_std_logic_vector(8, 8),
12588 => conv_std_logic_vector(8, 8),
12589 => conv_std_logic_vector(8, 8),
12590 => conv_std_logic_vector(8, 8),
12591 => conv_std_logic_vector(8, 8),
12592 => conv_std_logic_vector(9, 8),
12593 => conv_std_logic_vector(9, 8),
12594 => conv_std_logic_vector(9, 8),
12595 => conv_std_logic_vector(9, 8),
12596 => conv_std_logic_vector(9, 8),
12597 => conv_std_logic_vector(10, 8),
12598 => conv_std_logic_vector(10, 8),
12599 => conv_std_logic_vector(10, 8),
12600 => conv_std_logic_vector(10, 8),
12601 => conv_std_logic_vector(10, 8),
12602 => conv_std_logic_vector(11, 8),
12603 => conv_std_logic_vector(11, 8),
12604 => conv_std_logic_vector(11, 8),
12605 => conv_std_logic_vector(11, 8),
12606 => conv_std_logic_vector(11, 8),
12607 => conv_std_logic_vector(12, 8),
12608 => conv_std_logic_vector(12, 8),
12609 => conv_std_logic_vector(12, 8),
12610 => conv_std_logic_vector(12, 8),
12611 => conv_std_logic_vector(12, 8),
12612 => conv_std_logic_vector(13, 8),
12613 => conv_std_logic_vector(13, 8),
12614 => conv_std_logic_vector(13, 8),
12615 => conv_std_logic_vector(13, 8),
12616 => conv_std_logic_vector(13, 8),
12617 => conv_std_logic_vector(13, 8),
12618 => conv_std_logic_vector(14, 8),
12619 => conv_std_logic_vector(14, 8),
12620 => conv_std_logic_vector(14, 8),
12621 => conv_std_logic_vector(14, 8),
12622 => conv_std_logic_vector(14, 8),
12623 => conv_std_logic_vector(15, 8),
12624 => conv_std_logic_vector(15, 8),
12625 => conv_std_logic_vector(15, 8),
12626 => conv_std_logic_vector(15, 8),
12627 => conv_std_logic_vector(15, 8),
12628 => conv_std_logic_vector(16, 8),
12629 => conv_std_logic_vector(16, 8),
12630 => conv_std_logic_vector(16, 8),
12631 => conv_std_logic_vector(16, 8),
12632 => conv_std_logic_vector(16, 8),
12633 => conv_std_logic_vector(17, 8),
12634 => conv_std_logic_vector(17, 8),
12635 => conv_std_logic_vector(17, 8),
12636 => conv_std_logic_vector(17, 8),
12637 => conv_std_logic_vector(17, 8),
12638 => conv_std_logic_vector(17, 8),
12639 => conv_std_logic_vector(18, 8),
12640 => conv_std_logic_vector(18, 8),
12641 => conv_std_logic_vector(18, 8),
12642 => conv_std_logic_vector(18, 8),
12643 => conv_std_logic_vector(18, 8),
12644 => conv_std_logic_vector(19, 8),
12645 => conv_std_logic_vector(19, 8),
12646 => conv_std_logic_vector(19, 8),
12647 => conv_std_logic_vector(19, 8),
12648 => conv_std_logic_vector(19, 8),
12649 => conv_std_logic_vector(20, 8),
12650 => conv_std_logic_vector(20, 8),
12651 => conv_std_logic_vector(20, 8),
12652 => conv_std_logic_vector(20, 8),
12653 => conv_std_logic_vector(20, 8),
12654 => conv_std_logic_vector(21, 8),
12655 => conv_std_logic_vector(21, 8),
12656 => conv_std_logic_vector(21, 8),
12657 => conv_std_logic_vector(21, 8),
12658 => conv_std_logic_vector(21, 8),
12659 => conv_std_logic_vector(22, 8),
12660 => conv_std_logic_vector(22, 8),
12661 => conv_std_logic_vector(22, 8),
12662 => conv_std_logic_vector(22, 8),
12663 => conv_std_logic_vector(22, 8),
12664 => conv_std_logic_vector(22, 8),
12665 => conv_std_logic_vector(23, 8),
12666 => conv_std_logic_vector(23, 8),
12667 => conv_std_logic_vector(23, 8),
12668 => conv_std_logic_vector(23, 8),
12669 => conv_std_logic_vector(23, 8),
12670 => conv_std_logic_vector(24, 8),
12671 => conv_std_logic_vector(24, 8),
12672 => conv_std_logic_vector(24, 8),
12673 => conv_std_logic_vector(24, 8),
12674 => conv_std_logic_vector(24, 8),
12675 => conv_std_logic_vector(25, 8),
12676 => conv_std_logic_vector(25, 8),
12677 => conv_std_logic_vector(25, 8),
12678 => conv_std_logic_vector(25, 8),
12679 => conv_std_logic_vector(25, 8),
12680 => conv_std_logic_vector(26, 8),
12681 => conv_std_logic_vector(26, 8),
12682 => conv_std_logic_vector(26, 8),
12683 => conv_std_logic_vector(26, 8),
12684 => conv_std_logic_vector(26, 8),
12685 => conv_std_logic_vector(26, 8),
12686 => conv_std_logic_vector(27, 8),
12687 => conv_std_logic_vector(27, 8),
12688 => conv_std_logic_vector(27, 8),
12689 => conv_std_logic_vector(27, 8),
12690 => conv_std_logic_vector(27, 8),
12691 => conv_std_logic_vector(28, 8),
12692 => conv_std_logic_vector(28, 8),
12693 => conv_std_logic_vector(28, 8),
12694 => conv_std_logic_vector(28, 8),
12695 => conv_std_logic_vector(28, 8),
12696 => conv_std_logic_vector(29, 8),
12697 => conv_std_logic_vector(29, 8),
12698 => conv_std_logic_vector(29, 8),
12699 => conv_std_logic_vector(29, 8),
12700 => conv_std_logic_vector(29, 8),
12701 => conv_std_logic_vector(30, 8),
12702 => conv_std_logic_vector(30, 8),
12703 => conv_std_logic_vector(30, 8),
12704 => conv_std_logic_vector(30, 8),
12705 => conv_std_logic_vector(30, 8),
12706 => conv_std_logic_vector(31, 8),
12707 => conv_std_logic_vector(31, 8),
12708 => conv_std_logic_vector(31, 8),
12709 => conv_std_logic_vector(31, 8),
12710 => conv_std_logic_vector(31, 8),
12711 => conv_std_logic_vector(31, 8),
12712 => conv_std_logic_vector(32, 8),
12713 => conv_std_logic_vector(32, 8),
12714 => conv_std_logic_vector(32, 8),
12715 => conv_std_logic_vector(32, 8),
12716 => conv_std_logic_vector(32, 8),
12717 => conv_std_logic_vector(33, 8),
12718 => conv_std_logic_vector(33, 8),
12719 => conv_std_logic_vector(33, 8),
12720 => conv_std_logic_vector(33, 8),
12721 => conv_std_logic_vector(33, 8),
12722 => conv_std_logic_vector(34, 8),
12723 => conv_std_logic_vector(34, 8),
12724 => conv_std_logic_vector(34, 8),
12725 => conv_std_logic_vector(34, 8),
12726 => conv_std_logic_vector(34, 8),
12727 => conv_std_logic_vector(35, 8),
12728 => conv_std_logic_vector(35, 8),
12729 => conv_std_logic_vector(35, 8),
12730 => conv_std_logic_vector(35, 8),
12731 => conv_std_logic_vector(35, 8),
12732 => conv_std_logic_vector(35, 8),
12733 => conv_std_logic_vector(36, 8),
12734 => conv_std_logic_vector(36, 8),
12735 => conv_std_logic_vector(36, 8),
12736 => conv_std_logic_vector(36, 8),
12737 => conv_std_logic_vector(36, 8),
12738 => conv_std_logic_vector(37, 8),
12739 => conv_std_logic_vector(37, 8),
12740 => conv_std_logic_vector(37, 8),
12741 => conv_std_logic_vector(37, 8),
12742 => conv_std_logic_vector(37, 8),
12743 => conv_std_logic_vector(38, 8),
12744 => conv_std_logic_vector(38, 8),
12745 => conv_std_logic_vector(38, 8),
12746 => conv_std_logic_vector(38, 8),
12747 => conv_std_logic_vector(38, 8),
12748 => conv_std_logic_vector(39, 8),
12749 => conv_std_logic_vector(39, 8),
12750 => conv_std_logic_vector(39, 8),
12751 => conv_std_logic_vector(39, 8),
12752 => conv_std_logic_vector(39, 8),
12753 => conv_std_logic_vector(40, 8),
12754 => conv_std_logic_vector(40, 8),
12755 => conv_std_logic_vector(40, 8),
12756 => conv_std_logic_vector(40, 8),
12757 => conv_std_logic_vector(40, 8),
12758 => conv_std_logic_vector(40, 8),
12759 => conv_std_logic_vector(41, 8),
12760 => conv_std_logic_vector(41, 8),
12761 => conv_std_logic_vector(41, 8),
12762 => conv_std_logic_vector(41, 8),
12763 => conv_std_logic_vector(41, 8),
12764 => conv_std_logic_vector(42, 8),
12765 => conv_std_logic_vector(42, 8),
12766 => conv_std_logic_vector(42, 8),
12767 => conv_std_logic_vector(42, 8),
12768 => conv_std_logic_vector(42, 8),
12769 => conv_std_logic_vector(43, 8),
12770 => conv_std_logic_vector(43, 8),
12771 => conv_std_logic_vector(43, 8),
12772 => conv_std_logic_vector(43, 8),
12773 => conv_std_logic_vector(43, 8),
12774 => conv_std_logic_vector(44, 8),
12775 => conv_std_logic_vector(44, 8),
12776 => conv_std_logic_vector(44, 8),
12777 => conv_std_logic_vector(44, 8),
12778 => conv_std_logic_vector(44, 8),
12779 => conv_std_logic_vector(44, 8),
12780 => conv_std_logic_vector(45, 8),
12781 => conv_std_logic_vector(45, 8),
12782 => conv_std_logic_vector(45, 8),
12783 => conv_std_logic_vector(45, 8),
12784 => conv_std_logic_vector(45, 8),
12785 => conv_std_logic_vector(46, 8),
12786 => conv_std_logic_vector(46, 8),
12787 => conv_std_logic_vector(46, 8),
12788 => conv_std_logic_vector(46, 8),
12789 => conv_std_logic_vector(46, 8),
12790 => conv_std_logic_vector(47, 8),
12791 => conv_std_logic_vector(47, 8),
12792 => conv_std_logic_vector(47, 8),
12793 => conv_std_logic_vector(47, 8),
12794 => conv_std_logic_vector(47, 8),
12795 => conv_std_logic_vector(48, 8),
12796 => conv_std_logic_vector(48, 8),
12797 => conv_std_logic_vector(48, 8),
12798 => conv_std_logic_vector(48, 8),
12799 => conv_std_logic_vector(48, 8),
12800 => conv_std_logic_vector(0, 8),
12801 => conv_std_logic_vector(0, 8),
12802 => conv_std_logic_vector(0, 8),
12803 => conv_std_logic_vector(0, 8),
12804 => conv_std_logic_vector(0, 8),
12805 => conv_std_logic_vector(0, 8),
12806 => conv_std_logic_vector(1, 8),
12807 => conv_std_logic_vector(1, 8),
12808 => conv_std_logic_vector(1, 8),
12809 => conv_std_logic_vector(1, 8),
12810 => conv_std_logic_vector(1, 8),
12811 => conv_std_logic_vector(2, 8),
12812 => conv_std_logic_vector(2, 8),
12813 => conv_std_logic_vector(2, 8),
12814 => conv_std_logic_vector(2, 8),
12815 => conv_std_logic_vector(2, 8),
12816 => conv_std_logic_vector(3, 8),
12817 => conv_std_logic_vector(3, 8),
12818 => conv_std_logic_vector(3, 8),
12819 => conv_std_logic_vector(3, 8),
12820 => conv_std_logic_vector(3, 8),
12821 => conv_std_logic_vector(4, 8),
12822 => conv_std_logic_vector(4, 8),
12823 => conv_std_logic_vector(4, 8),
12824 => conv_std_logic_vector(4, 8),
12825 => conv_std_logic_vector(4, 8),
12826 => conv_std_logic_vector(5, 8),
12827 => conv_std_logic_vector(5, 8),
12828 => conv_std_logic_vector(5, 8),
12829 => conv_std_logic_vector(5, 8),
12830 => conv_std_logic_vector(5, 8),
12831 => conv_std_logic_vector(6, 8),
12832 => conv_std_logic_vector(6, 8),
12833 => conv_std_logic_vector(6, 8),
12834 => conv_std_logic_vector(6, 8),
12835 => conv_std_logic_vector(6, 8),
12836 => conv_std_logic_vector(7, 8),
12837 => conv_std_logic_vector(7, 8),
12838 => conv_std_logic_vector(7, 8),
12839 => conv_std_logic_vector(7, 8),
12840 => conv_std_logic_vector(7, 8),
12841 => conv_std_logic_vector(8, 8),
12842 => conv_std_logic_vector(8, 8),
12843 => conv_std_logic_vector(8, 8),
12844 => conv_std_logic_vector(8, 8),
12845 => conv_std_logic_vector(8, 8),
12846 => conv_std_logic_vector(8, 8),
12847 => conv_std_logic_vector(9, 8),
12848 => conv_std_logic_vector(9, 8),
12849 => conv_std_logic_vector(9, 8),
12850 => conv_std_logic_vector(9, 8),
12851 => conv_std_logic_vector(9, 8),
12852 => conv_std_logic_vector(10, 8),
12853 => conv_std_logic_vector(10, 8),
12854 => conv_std_logic_vector(10, 8),
12855 => conv_std_logic_vector(10, 8),
12856 => conv_std_logic_vector(10, 8),
12857 => conv_std_logic_vector(11, 8),
12858 => conv_std_logic_vector(11, 8),
12859 => conv_std_logic_vector(11, 8),
12860 => conv_std_logic_vector(11, 8),
12861 => conv_std_logic_vector(11, 8),
12862 => conv_std_logic_vector(12, 8),
12863 => conv_std_logic_vector(12, 8),
12864 => conv_std_logic_vector(12, 8),
12865 => conv_std_logic_vector(12, 8),
12866 => conv_std_logic_vector(12, 8),
12867 => conv_std_logic_vector(13, 8),
12868 => conv_std_logic_vector(13, 8),
12869 => conv_std_logic_vector(13, 8),
12870 => conv_std_logic_vector(13, 8),
12871 => conv_std_logic_vector(13, 8),
12872 => conv_std_logic_vector(14, 8),
12873 => conv_std_logic_vector(14, 8),
12874 => conv_std_logic_vector(14, 8),
12875 => conv_std_logic_vector(14, 8),
12876 => conv_std_logic_vector(14, 8),
12877 => conv_std_logic_vector(15, 8),
12878 => conv_std_logic_vector(15, 8),
12879 => conv_std_logic_vector(15, 8),
12880 => conv_std_logic_vector(15, 8),
12881 => conv_std_logic_vector(15, 8),
12882 => conv_std_logic_vector(16, 8),
12883 => conv_std_logic_vector(16, 8),
12884 => conv_std_logic_vector(16, 8),
12885 => conv_std_logic_vector(16, 8),
12886 => conv_std_logic_vector(16, 8),
12887 => conv_std_logic_vector(16, 8),
12888 => conv_std_logic_vector(17, 8),
12889 => conv_std_logic_vector(17, 8),
12890 => conv_std_logic_vector(17, 8),
12891 => conv_std_logic_vector(17, 8),
12892 => conv_std_logic_vector(17, 8),
12893 => conv_std_logic_vector(18, 8),
12894 => conv_std_logic_vector(18, 8),
12895 => conv_std_logic_vector(18, 8),
12896 => conv_std_logic_vector(18, 8),
12897 => conv_std_logic_vector(18, 8),
12898 => conv_std_logic_vector(19, 8),
12899 => conv_std_logic_vector(19, 8),
12900 => conv_std_logic_vector(19, 8),
12901 => conv_std_logic_vector(19, 8),
12902 => conv_std_logic_vector(19, 8),
12903 => conv_std_logic_vector(20, 8),
12904 => conv_std_logic_vector(20, 8),
12905 => conv_std_logic_vector(20, 8),
12906 => conv_std_logic_vector(20, 8),
12907 => conv_std_logic_vector(20, 8),
12908 => conv_std_logic_vector(21, 8),
12909 => conv_std_logic_vector(21, 8),
12910 => conv_std_logic_vector(21, 8),
12911 => conv_std_logic_vector(21, 8),
12912 => conv_std_logic_vector(21, 8),
12913 => conv_std_logic_vector(22, 8),
12914 => conv_std_logic_vector(22, 8),
12915 => conv_std_logic_vector(22, 8),
12916 => conv_std_logic_vector(22, 8),
12917 => conv_std_logic_vector(22, 8),
12918 => conv_std_logic_vector(23, 8),
12919 => conv_std_logic_vector(23, 8),
12920 => conv_std_logic_vector(23, 8),
12921 => conv_std_logic_vector(23, 8),
12922 => conv_std_logic_vector(23, 8),
12923 => conv_std_logic_vector(24, 8),
12924 => conv_std_logic_vector(24, 8),
12925 => conv_std_logic_vector(24, 8),
12926 => conv_std_logic_vector(24, 8),
12927 => conv_std_logic_vector(24, 8),
12928 => conv_std_logic_vector(25, 8),
12929 => conv_std_logic_vector(25, 8),
12930 => conv_std_logic_vector(25, 8),
12931 => conv_std_logic_vector(25, 8),
12932 => conv_std_logic_vector(25, 8),
12933 => conv_std_logic_vector(25, 8),
12934 => conv_std_logic_vector(26, 8),
12935 => conv_std_logic_vector(26, 8),
12936 => conv_std_logic_vector(26, 8),
12937 => conv_std_logic_vector(26, 8),
12938 => conv_std_logic_vector(26, 8),
12939 => conv_std_logic_vector(27, 8),
12940 => conv_std_logic_vector(27, 8),
12941 => conv_std_logic_vector(27, 8),
12942 => conv_std_logic_vector(27, 8),
12943 => conv_std_logic_vector(27, 8),
12944 => conv_std_logic_vector(28, 8),
12945 => conv_std_logic_vector(28, 8),
12946 => conv_std_logic_vector(28, 8),
12947 => conv_std_logic_vector(28, 8),
12948 => conv_std_logic_vector(28, 8),
12949 => conv_std_logic_vector(29, 8),
12950 => conv_std_logic_vector(29, 8),
12951 => conv_std_logic_vector(29, 8),
12952 => conv_std_logic_vector(29, 8),
12953 => conv_std_logic_vector(29, 8),
12954 => conv_std_logic_vector(30, 8),
12955 => conv_std_logic_vector(30, 8),
12956 => conv_std_logic_vector(30, 8),
12957 => conv_std_logic_vector(30, 8),
12958 => conv_std_logic_vector(30, 8),
12959 => conv_std_logic_vector(31, 8),
12960 => conv_std_logic_vector(31, 8),
12961 => conv_std_logic_vector(31, 8),
12962 => conv_std_logic_vector(31, 8),
12963 => conv_std_logic_vector(31, 8),
12964 => conv_std_logic_vector(32, 8),
12965 => conv_std_logic_vector(32, 8),
12966 => conv_std_logic_vector(32, 8),
12967 => conv_std_logic_vector(32, 8),
12968 => conv_std_logic_vector(32, 8),
12969 => conv_std_logic_vector(33, 8),
12970 => conv_std_logic_vector(33, 8),
12971 => conv_std_logic_vector(33, 8),
12972 => conv_std_logic_vector(33, 8),
12973 => conv_std_logic_vector(33, 8),
12974 => conv_std_logic_vector(33, 8),
12975 => conv_std_logic_vector(34, 8),
12976 => conv_std_logic_vector(34, 8),
12977 => conv_std_logic_vector(34, 8),
12978 => conv_std_logic_vector(34, 8),
12979 => conv_std_logic_vector(34, 8),
12980 => conv_std_logic_vector(35, 8),
12981 => conv_std_logic_vector(35, 8),
12982 => conv_std_logic_vector(35, 8),
12983 => conv_std_logic_vector(35, 8),
12984 => conv_std_logic_vector(35, 8),
12985 => conv_std_logic_vector(36, 8),
12986 => conv_std_logic_vector(36, 8),
12987 => conv_std_logic_vector(36, 8),
12988 => conv_std_logic_vector(36, 8),
12989 => conv_std_logic_vector(36, 8),
12990 => conv_std_logic_vector(37, 8),
12991 => conv_std_logic_vector(37, 8),
12992 => conv_std_logic_vector(37, 8),
12993 => conv_std_logic_vector(37, 8),
12994 => conv_std_logic_vector(37, 8),
12995 => conv_std_logic_vector(38, 8),
12996 => conv_std_logic_vector(38, 8),
12997 => conv_std_logic_vector(38, 8),
12998 => conv_std_logic_vector(38, 8),
12999 => conv_std_logic_vector(38, 8),
13000 => conv_std_logic_vector(39, 8),
13001 => conv_std_logic_vector(39, 8),
13002 => conv_std_logic_vector(39, 8),
13003 => conv_std_logic_vector(39, 8),
13004 => conv_std_logic_vector(39, 8),
13005 => conv_std_logic_vector(40, 8),
13006 => conv_std_logic_vector(40, 8),
13007 => conv_std_logic_vector(40, 8),
13008 => conv_std_logic_vector(40, 8),
13009 => conv_std_logic_vector(40, 8),
13010 => conv_std_logic_vector(41, 8),
13011 => conv_std_logic_vector(41, 8),
13012 => conv_std_logic_vector(41, 8),
13013 => conv_std_logic_vector(41, 8),
13014 => conv_std_logic_vector(41, 8),
13015 => conv_std_logic_vector(41, 8),
13016 => conv_std_logic_vector(42, 8),
13017 => conv_std_logic_vector(42, 8),
13018 => conv_std_logic_vector(42, 8),
13019 => conv_std_logic_vector(42, 8),
13020 => conv_std_logic_vector(42, 8),
13021 => conv_std_logic_vector(43, 8),
13022 => conv_std_logic_vector(43, 8),
13023 => conv_std_logic_vector(43, 8),
13024 => conv_std_logic_vector(43, 8),
13025 => conv_std_logic_vector(43, 8),
13026 => conv_std_logic_vector(44, 8),
13027 => conv_std_logic_vector(44, 8),
13028 => conv_std_logic_vector(44, 8),
13029 => conv_std_logic_vector(44, 8),
13030 => conv_std_logic_vector(44, 8),
13031 => conv_std_logic_vector(45, 8),
13032 => conv_std_logic_vector(45, 8),
13033 => conv_std_logic_vector(45, 8),
13034 => conv_std_logic_vector(45, 8),
13035 => conv_std_logic_vector(45, 8),
13036 => conv_std_logic_vector(46, 8),
13037 => conv_std_logic_vector(46, 8),
13038 => conv_std_logic_vector(46, 8),
13039 => conv_std_logic_vector(46, 8),
13040 => conv_std_logic_vector(46, 8),
13041 => conv_std_logic_vector(47, 8),
13042 => conv_std_logic_vector(47, 8),
13043 => conv_std_logic_vector(47, 8),
13044 => conv_std_logic_vector(47, 8),
13045 => conv_std_logic_vector(47, 8),
13046 => conv_std_logic_vector(48, 8),
13047 => conv_std_logic_vector(48, 8),
13048 => conv_std_logic_vector(48, 8),
13049 => conv_std_logic_vector(48, 8),
13050 => conv_std_logic_vector(48, 8),
13051 => conv_std_logic_vector(49, 8),
13052 => conv_std_logic_vector(49, 8),
13053 => conv_std_logic_vector(49, 8),
13054 => conv_std_logic_vector(49, 8),
13055 => conv_std_logic_vector(49, 8),
13056 => conv_std_logic_vector(0, 8),
13057 => conv_std_logic_vector(0, 8),
13058 => conv_std_logic_vector(0, 8),
13059 => conv_std_logic_vector(0, 8),
13060 => conv_std_logic_vector(0, 8),
13061 => conv_std_logic_vector(0, 8),
13062 => conv_std_logic_vector(1, 8),
13063 => conv_std_logic_vector(1, 8),
13064 => conv_std_logic_vector(1, 8),
13065 => conv_std_logic_vector(1, 8),
13066 => conv_std_logic_vector(1, 8),
13067 => conv_std_logic_vector(2, 8),
13068 => conv_std_logic_vector(2, 8),
13069 => conv_std_logic_vector(2, 8),
13070 => conv_std_logic_vector(2, 8),
13071 => conv_std_logic_vector(2, 8),
13072 => conv_std_logic_vector(3, 8),
13073 => conv_std_logic_vector(3, 8),
13074 => conv_std_logic_vector(3, 8),
13075 => conv_std_logic_vector(3, 8),
13076 => conv_std_logic_vector(3, 8),
13077 => conv_std_logic_vector(4, 8),
13078 => conv_std_logic_vector(4, 8),
13079 => conv_std_logic_vector(4, 8),
13080 => conv_std_logic_vector(4, 8),
13081 => conv_std_logic_vector(4, 8),
13082 => conv_std_logic_vector(5, 8),
13083 => conv_std_logic_vector(5, 8),
13084 => conv_std_logic_vector(5, 8),
13085 => conv_std_logic_vector(5, 8),
13086 => conv_std_logic_vector(5, 8),
13087 => conv_std_logic_vector(6, 8),
13088 => conv_std_logic_vector(6, 8),
13089 => conv_std_logic_vector(6, 8),
13090 => conv_std_logic_vector(6, 8),
13091 => conv_std_logic_vector(6, 8),
13092 => conv_std_logic_vector(7, 8),
13093 => conv_std_logic_vector(7, 8),
13094 => conv_std_logic_vector(7, 8),
13095 => conv_std_logic_vector(7, 8),
13096 => conv_std_logic_vector(7, 8),
13097 => conv_std_logic_vector(8, 8),
13098 => conv_std_logic_vector(8, 8),
13099 => conv_std_logic_vector(8, 8),
13100 => conv_std_logic_vector(8, 8),
13101 => conv_std_logic_vector(8, 8),
13102 => conv_std_logic_vector(9, 8),
13103 => conv_std_logic_vector(9, 8),
13104 => conv_std_logic_vector(9, 8),
13105 => conv_std_logic_vector(9, 8),
13106 => conv_std_logic_vector(9, 8),
13107 => conv_std_logic_vector(10, 8),
13108 => conv_std_logic_vector(10, 8),
13109 => conv_std_logic_vector(10, 8),
13110 => conv_std_logic_vector(10, 8),
13111 => conv_std_logic_vector(10, 8),
13112 => conv_std_logic_vector(11, 8),
13113 => conv_std_logic_vector(11, 8),
13114 => conv_std_logic_vector(11, 8),
13115 => conv_std_logic_vector(11, 8),
13116 => conv_std_logic_vector(11, 8),
13117 => conv_std_logic_vector(12, 8),
13118 => conv_std_logic_vector(12, 8),
13119 => conv_std_logic_vector(12, 8),
13120 => conv_std_logic_vector(12, 8),
13121 => conv_std_logic_vector(12, 8),
13122 => conv_std_logic_vector(13, 8),
13123 => conv_std_logic_vector(13, 8),
13124 => conv_std_logic_vector(13, 8),
13125 => conv_std_logic_vector(13, 8),
13126 => conv_std_logic_vector(13, 8),
13127 => conv_std_logic_vector(14, 8),
13128 => conv_std_logic_vector(14, 8),
13129 => conv_std_logic_vector(14, 8),
13130 => conv_std_logic_vector(14, 8),
13131 => conv_std_logic_vector(14, 8),
13132 => conv_std_logic_vector(15, 8),
13133 => conv_std_logic_vector(15, 8),
13134 => conv_std_logic_vector(15, 8),
13135 => conv_std_logic_vector(15, 8),
13136 => conv_std_logic_vector(15, 8),
13137 => conv_std_logic_vector(16, 8),
13138 => conv_std_logic_vector(16, 8),
13139 => conv_std_logic_vector(16, 8),
13140 => conv_std_logic_vector(16, 8),
13141 => conv_std_logic_vector(16, 8),
13142 => conv_std_logic_vector(17, 8),
13143 => conv_std_logic_vector(17, 8),
13144 => conv_std_logic_vector(17, 8),
13145 => conv_std_logic_vector(17, 8),
13146 => conv_std_logic_vector(17, 8),
13147 => conv_std_logic_vector(18, 8),
13148 => conv_std_logic_vector(18, 8),
13149 => conv_std_logic_vector(18, 8),
13150 => conv_std_logic_vector(18, 8),
13151 => conv_std_logic_vector(18, 8),
13152 => conv_std_logic_vector(19, 8),
13153 => conv_std_logic_vector(19, 8),
13154 => conv_std_logic_vector(19, 8),
13155 => conv_std_logic_vector(19, 8),
13156 => conv_std_logic_vector(19, 8),
13157 => conv_std_logic_vector(20, 8),
13158 => conv_std_logic_vector(20, 8),
13159 => conv_std_logic_vector(20, 8),
13160 => conv_std_logic_vector(20, 8),
13161 => conv_std_logic_vector(20, 8),
13162 => conv_std_logic_vector(21, 8),
13163 => conv_std_logic_vector(21, 8),
13164 => conv_std_logic_vector(21, 8),
13165 => conv_std_logic_vector(21, 8),
13166 => conv_std_logic_vector(21, 8),
13167 => conv_std_logic_vector(22, 8),
13168 => conv_std_logic_vector(22, 8),
13169 => conv_std_logic_vector(22, 8),
13170 => conv_std_logic_vector(22, 8),
13171 => conv_std_logic_vector(22, 8),
13172 => conv_std_logic_vector(23, 8),
13173 => conv_std_logic_vector(23, 8),
13174 => conv_std_logic_vector(23, 8),
13175 => conv_std_logic_vector(23, 8),
13176 => conv_std_logic_vector(23, 8),
13177 => conv_std_logic_vector(24, 8),
13178 => conv_std_logic_vector(24, 8),
13179 => conv_std_logic_vector(24, 8),
13180 => conv_std_logic_vector(24, 8),
13181 => conv_std_logic_vector(24, 8),
13182 => conv_std_logic_vector(25, 8),
13183 => conv_std_logic_vector(25, 8),
13184 => conv_std_logic_vector(25, 8),
13185 => conv_std_logic_vector(25, 8),
13186 => conv_std_logic_vector(25, 8),
13187 => conv_std_logic_vector(26, 8),
13188 => conv_std_logic_vector(26, 8),
13189 => conv_std_logic_vector(26, 8),
13190 => conv_std_logic_vector(26, 8),
13191 => conv_std_logic_vector(26, 8),
13192 => conv_std_logic_vector(27, 8),
13193 => conv_std_logic_vector(27, 8),
13194 => conv_std_logic_vector(27, 8),
13195 => conv_std_logic_vector(27, 8),
13196 => conv_std_logic_vector(27, 8),
13197 => conv_std_logic_vector(28, 8),
13198 => conv_std_logic_vector(28, 8),
13199 => conv_std_logic_vector(28, 8),
13200 => conv_std_logic_vector(28, 8),
13201 => conv_std_logic_vector(28, 8),
13202 => conv_std_logic_vector(29, 8),
13203 => conv_std_logic_vector(29, 8),
13204 => conv_std_logic_vector(29, 8),
13205 => conv_std_logic_vector(29, 8),
13206 => conv_std_logic_vector(29, 8),
13207 => conv_std_logic_vector(30, 8),
13208 => conv_std_logic_vector(30, 8),
13209 => conv_std_logic_vector(30, 8),
13210 => conv_std_logic_vector(30, 8),
13211 => conv_std_logic_vector(30, 8),
13212 => conv_std_logic_vector(31, 8),
13213 => conv_std_logic_vector(31, 8),
13214 => conv_std_logic_vector(31, 8),
13215 => conv_std_logic_vector(31, 8),
13216 => conv_std_logic_vector(31, 8),
13217 => conv_std_logic_vector(32, 8),
13218 => conv_std_logic_vector(32, 8),
13219 => conv_std_logic_vector(32, 8),
13220 => conv_std_logic_vector(32, 8),
13221 => conv_std_logic_vector(32, 8),
13222 => conv_std_logic_vector(33, 8),
13223 => conv_std_logic_vector(33, 8),
13224 => conv_std_logic_vector(33, 8),
13225 => conv_std_logic_vector(33, 8),
13226 => conv_std_logic_vector(33, 8),
13227 => conv_std_logic_vector(34, 8),
13228 => conv_std_logic_vector(34, 8),
13229 => conv_std_logic_vector(34, 8),
13230 => conv_std_logic_vector(34, 8),
13231 => conv_std_logic_vector(34, 8),
13232 => conv_std_logic_vector(35, 8),
13233 => conv_std_logic_vector(35, 8),
13234 => conv_std_logic_vector(35, 8),
13235 => conv_std_logic_vector(35, 8),
13236 => conv_std_logic_vector(35, 8),
13237 => conv_std_logic_vector(36, 8),
13238 => conv_std_logic_vector(36, 8),
13239 => conv_std_logic_vector(36, 8),
13240 => conv_std_logic_vector(36, 8),
13241 => conv_std_logic_vector(36, 8),
13242 => conv_std_logic_vector(37, 8),
13243 => conv_std_logic_vector(37, 8),
13244 => conv_std_logic_vector(37, 8),
13245 => conv_std_logic_vector(37, 8),
13246 => conv_std_logic_vector(37, 8),
13247 => conv_std_logic_vector(38, 8),
13248 => conv_std_logic_vector(38, 8),
13249 => conv_std_logic_vector(38, 8),
13250 => conv_std_logic_vector(38, 8),
13251 => conv_std_logic_vector(38, 8),
13252 => conv_std_logic_vector(39, 8),
13253 => conv_std_logic_vector(39, 8),
13254 => conv_std_logic_vector(39, 8),
13255 => conv_std_logic_vector(39, 8),
13256 => conv_std_logic_vector(39, 8),
13257 => conv_std_logic_vector(40, 8),
13258 => conv_std_logic_vector(40, 8),
13259 => conv_std_logic_vector(40, 8),
13260 => conv_std_logic_vector(40, 8),
13261 => conv_std_logic_vector(40, 8),
13262 => conv_std_logic_vector(41, 8),
13263 => conv_std_logic_vector(41, 8),
13264 => conv_std_logic_vector(41, 8),
13265 => conv_std_logic_vector(41, 8),
13266 => conv_std_logic_vector(41, 8),
13267 => conv_std_logic_vector(42, 8),
13268 => conv_std_logic_vector(42, 8),
13269 => conv_std_logic_vector(42, 8),
13270 => conv_std_logic_vector(42, 8),
13271 => conv_std_logic_vector(42, 8),
13272 => conv_std_logic_vector(43, 8),
13273 => conv_std_logic_vector(43, 8),
13274 => conv_std_logic_vector(43, 8),
13275 => conv_std_logic_vector(43, 8),
13276 => conv_std_logic_vector(43, 8),
13277 => conv_std_logic_vector(44, 8),
13278 => conv_std_logic_vector(44, 8),
13279 => conv_std_logic_vector(44, 8),
13280 => conv_std_logic_vector(44, 8),
13281 => conv_std_logic_vector(44, 8),
13282 => conv_std_logic_vector(45, 8),
13283 => conv_std_logic_vector(45, 8),
13284 => conv_std_logic_vector(45, 8),
13285 => conv_std_logic_vector(45, 8),
13286 => conv_std_logic_vector(45, 8),
13287 => conv_std_logic_vector(46, 8),
13288 => conv_std_logic_vector(46, 8),
13289 => conv_std_logic_vector(46, 8),
13290 => conv_std_logic_vector(46, 8),
13291 => conv_std_logic_vector(46, 8),
13292 => conv_std_logic_vector(47, 8),
13293 => conv_std_logic_vector(47, 8),
13294 => conv_std_logic_vector(47, 8),
13295 => conv_std_logic_vector(47, 8),
13296 => conv_std_logic_vector(47, 8),
13297 => conv_std_logic_vector(48, 8),
13298 => conv_std_logic_vector(48, 8),
13299 => conv_std_logic_vector(48, 8),
13300 => conv_std_logic_vector(48, 8),
13301 => conv_std_logic_vector(48, 8),
13302 => conv_std_logic_vector(49, 8),
13303 => conv_std_logic_vector(49, 8),
13304 => conv_std_logic_vector(49, 8),
13305 => conv_std_logic_vector(49, 8),
13306 => conv_std_logic_vector(49, 8),
13307 => conv_std_logic_vector(50, 8),
13308 => conv_std_logic_vector(50, 8),
13309 => conv_std_logic_vector(50, 8),
13310 => conv_std_logic_vector(50, 8),
13311 => conv_std_logic_vector(50, 8),
13312 => conv_std_logic_vector(0, 8),
13313 => conv_std_logic_vector(0, 8),
13314 => conv_std_logic_vector(0, 8),
13315 => conv_std_logic_vector(0, 8),
13316 => conv_std_logic_vector(0, 8),
13317 => conv_std_logic_vector(1, 8),
13318 => conv_std_logic_vector(1, 8),
13319 => conv_std_logic_vector(1, 8),
13320 => conv_std_logic_vector(1, 8),
13321 => conv_std_logic_vector(1, 8),
13322 => conv_std_logic_vector(2, 8),
13323 => conv_std_logic_vector(2, 8),
13324 => conv_std_logic_vector(2, 8),
13325 => conv_std_logic_vector(2, 8),
13326 => conv_std_logic_vector(2, 8),
13327 => conv_std_logic_vector(3, 8),
13328 => conv_std_logic_vector(3, 8),
13329 => conv_std_logic_vector(3, 8),
13330 => conv_std_logic_vector(3, 8),
13331 => conv_std_logic_vector(3, 8),
13332 => conv_std_logic_vector(4, 8),
13333 => conv_std_logic_vector(4, 8),
13334 => conv_std_logic_vector(4, 8),
13335 => conv_std_logic_vector(4, 8),
13336 => conv_std_logic_vector(4, 8),
13337 => conv_std_logic_vector(5, 8),
13338 => conv_std_logic_vector(5, 8),
13339 => conv_std_logic_vector(5, 8),
13340 => conv_std_logic_vector(5, 8),
13341 => conv_std_logic_vector(5, 8),
13342 => conv_std_logic_vector(6, 8),
13343 => conv_std_logic_vector(6, 8),
13344 => conv_std_logic_vector(6, 8),
13345 => conv_std_logic_vector(6, 8),
13346 => conv_std_logic_vector(6, 8),
13347 => conv_std_logic_vector(7, 8),
13348 => conv_std_logic_vector(7, 8),
13349 => conv_std_logic_vector(7, 8),
13350 => conv_std_logic_vector(7, 8),
13351 => conv_std_logic_vector(7, 8),
13352 => conv_std_logic_vector(8, 8),
13353 => conv_std_logic_vector(8, 8),
13354 => conv_std_logic_vector(8, 8),
13355 => conv_std_logic_vector(8, 8),
13356 => conv_std_logic_vector(8, 8),
13357 => conv_std_logic_vector(9, 8),
13358 => conv_std_logic_vector(9, 8),
13359 => conv_std_logic_vector(9, 8),
13360 => conv_std_logic_vector(9, 8),
13361 => conv_std_logic_vector(9, 8),
13362 => conv_std_logic_vector(10, 8),
13363 => conv_std_logic_vector(10, 8),
13364 => conv_std_logic_vector(10, 8),
13365 => conv_std_logic_vector(10, 8),
13366 => conv_std_logic_vector(10, 8),
13367 => conv_std_logic_vector(11, 8),
13368 => conv_std_logic_vector(11, 8),
13369 => conv_std_logic_vector(11, 8),
13370 => conv_std_logic_vector(11, 8),
13371 => conv_std_logic_vector(11, 8),
13372 => conv_std_logic_vector(12, 8),
13373 => conv_std_logic_vector(12, 8),
13374 => conv_std_logic_vector(12, 8),
13375 => conv_std_logic_vector(12, 8),
13376 => conv_std_logic_vector(13, 8),
13377 => conv_std_logic_vector(13, 8),
13378 => conv_std_logic_vector(13, 8),
13379 => conv_std_logic_vector(13, 8),
13380 => conv_std_logic_vector(13, 8),
13381 => conv_std_logic_vector(14, 8),
13382 => conv_std_logic_vector(14, 8),
13383 => conv_std_logic_vector(14, 8),
13384 => conv_std_logic_vector(14, 8),
13385 => conv_std_logic_vector(14, 8),
13386 => conv_std_logic_vector(15, 8),
13387 => conv_std_logic_vector(15, 8),
13388 => conv_std_logic_vector(15, 8),
13389 => conv_std_logic_vector(15, 8),
13390 => conv_std_logic_vector(15, 8),
13391 => conv_std_logic_vector(16, 8),
13392 => conv_std_logic_vector(16, 8),
13393 => conv_std_logic_vector(16, 8),
13394 => conv_std_logic_vector(16, 8),
13395 => conv_std_logic_vector(16, 8),
13396 => conv_std_logic_vector(17, 8),
13397 => conv_std_logic_vector(17, 8),
13398 => conv_std_logic_vector(17, 8),
13399 => conv_std_logic_vector(17, 8),
13400 => conv_std_logic_vector(17, 8),
13401 => conv_std_logic_vector(18, 8),
13402 => conv_std_logic_vector(18, 8),
13403 => conv_std_logic_vector(18, 8),
13404 => conv_std_logic_vector(18, 8),
13405 => conv_std_logic_vector(18, 8),
13406 => conv_std_logic_vector(19, 8),
13407 => conv_std_logic_vector(19, 8),
13408 => conv_std_logic_vector(19, 8),
13409 => conv_std_logic_vector(19, 8),
13410 => conv_std_logic_vector(19, 8),
13411 => conv_std_logic_vector(20, 8),
13412 => conv_std_logic_vector(20, 8),
13413 => conv_std_logic_vector(20, 8),
13414 => conv_std_logic_vector(20, 8),
13415 => conv_std_logic_vector(20, 8),
13416 => conv_std_logic_vector(21, 8),
13417 => conv_std_logic_vector(21, 8),
13418 => conv_std_logic_vector(21, 8),
13419 => conv_std_logic_vector(21, 8),
13420 => conv_std_logic_vector(21, 8),
13421 => conv_std_logic_vector(22, 8),
13422 => conv_std_logic_vector(22, 8),
13423 => conv_std_logic_vector(22, 8),
13424 => conv_std_logic_vector(22, 8),
13425 => conv_std_logic_vector(22, 8),
13426 => conv_std_logic_vector(23, 8),
13427 => conv_std_logic_vector(23, 8),
13428 => conv_std_logic_vector(23, 8),
13429 => conv_std_logic_vector(23, 8),
13430 => conv_std_logic_vector(23, 8),
13431 => conv_std_logic_vector(24, 8),
13432 => conv_std_logic_vector(24, 8),
13433 => conv_std_logic_vector(24, 8),
13434 => conv_std_logic_vector(24, 8),
13435 => conv_std_logic_vector(24, 8),
13436 => conv_std_logic_vector(25, 8),
13437 => conv_std_logic_vector(25, 8),
13438 => conv_std_logic_vector(25, 8),
13439 => conv_std_logic_vector(25, 8),
13440 => conv_std_logic_vector(26, 8),
13441 => conv_std_logic_vector(26, 8),
13442 => conv_std_logic_vector(26, 8),
13443 => conv_std_logic_vector(26, 8),
13444 => conv_std_logic_vector(26, 8),
13445 => conv_std_logic_vector(27, 8),
13446 => conv_std_logic_vector(27, 8),
13447 => conv_std_logic_vector(27, 8),
13448 => conv_std_logic_vector(27, 8),
13449 => conv_std_logic_vector(27, 8),
13450 => conv_std_logic_vector(28, 8),
13451 => conv_std_logic_vector(28, 8),
13452 => conv_std_logic_vector(28, 8),
13453 => conv_std_logic_vector(28, 8),
13454 => conv_std_logic_vector(28, 8),
13455 => conv_std_logic_vector(29, 8),
13456 => conv_std_logic_vector(29, 8),
13457 => conv_std_logic_vector(29, 8),
13458 => conv_std_logic_vector(29, 8),
13459 => conv_std_logic_vector(29, 8),
13460 => conv_std_logic_vector(30, 8),
13461 => conv_std_logic_vector(30, 8),
13462 => conv_std_logic_vector(30, 8),
13463 => conv_std_logic_vector(30, 8),
13464 => conv_std_logic_vector(30, 8),
13465 => conv_std_logic_vector(31, 8),
13466 => conv_std_logic_vector(31, 8),
13467 => conv_std_logic_vector(31, 8),
13468 => conv_std_logic_vector(31, 8),
13469 => conv_std_logic_vector(31, 8),
13470 => conv_std_logic_vector(32, 8),
13471 => conv_std_logic_vector(32, 8),
13472 => conv_std_logic_vector(32, 8),
13473 => conv_std_logic_vector(32, 8),
13474 => conv_std_logic_vector(32, 8),
13475 => conv_std_logic_vector(33, 8),
13476 => conv_std_logic_vector(33, 8),
13477 => conv_std_logic_vector(33, 8),
13478 => conv_std_logic_vector(33, 8),
13479 => conv_std_logic_vector(33, 8),
13480 => conv_std_logic_vector(34, 8),
13481 => conv_std_logic_vector(34, 8),
13482 => conv_std_logic_vector(34, 8),
13483 => conv_std_logic_vector(34, 8),
13484 => conv_std_logic_vector(34, 8),
13485 => conv_std_logic_vector(35, 8),
13486 => conv_std_logic_vector(35, 8),
13487 => conv_std_logic_vector(35, 8),
13488 => conv_std_logic_vector(35, 8),
13489 => conv_std_logic_vector(35, 8),
13490 => conv_std_logic_vector(36, 8),
13491 => conv_std_logic_vector(36, 8),
13492 => conv_std_logic_vector(36, 8),
13493 => conv_std_logic_vector(36, 8),
13494 => conv_std_logic_vector(36, 8),
13495 => conv_std_logic_vector(37, 8),
13496 => conv_std_logic_vector(37, 8),
13497 => conv_std_logic_vector(37, 8),
13498 => conv_std_logic_vector(37, 8),
13499 => conv_std_logic_vector(37, 8),
13500 => conv_std_logic_vector(38, 8),
13501 => conv_std_logic_vector(38, 8),
13502 => conv_std_logic_vector(38, 8),
13503 => conv_std_logic_vector(38, 8),
13504 => conv_std_logic_vector(39, 8),
13505 => conv_std_logic_vector(39, 8),
13506 => conv_std_logic_vector(39, 8),
13507 => conv_std_logic_vector(39, 8),
13508 => conv_std_logic_vector(39, 8),
13509 => conv_std_logic_vector(40, 8),
13510 => conv_std_logic_vector(40, 8),
13511 => conv_std_logic_vector(40, 8),
13512 => conv_std_logic_vector(40, 8),
13513 => conv_std_logic_vector(40, 8),
13514 => conv_std_logic_vector(41, 8),
13515 => conv_std_logic_vector(41, 8),
13516 => conv_std_logic_vector(41, 8),
13517 => conv_std_logic_vector(41, 8),
13518 => conv_std_logic_vector(41, 8),
13519 => conv_std_logic_vector(42, 8),
13520 => conv_std_logic_vector(42, 8),
13521 => conv_std_logic_vector(42, 8),
13522 => conv_std_logic_vector(42, 8),
13523 => conv_std_logic_vector(42, 8),
13524 => conv_std_logic_vector(43, 8),
13525 => conv_std_logic_vector(43, 8),
13526 => conv_std_logic_vector(43, 8),
13527 => conv_std_logic_vector(43, 8),
13528 => conv_std_logic_vector(43, 8),
13529 => conv_std_logic_vector(44, 8),
13530 => conv_std_logic_vector(44, 8),
13531 => conv_std_logic_vector(44, 8),
13532 => conv_std_logic_vector(44, 8),
13533 => conv_std_logic_vector(44, 8),
13534 => conv_std_logic_vector(45, 8),
13535 => conv_std_logic_vector(45, 8),
13536 => conv_std_logic_vector(45, 8),
13537 => conv_std_logic_vector(45, 8),
13538 => conv_std_logic_vector(45, 8),
13539 => conv_std_logic_vector(46, 8),
13540 => conv_std_logic_vector(46, 8),
13541 => conv_std_logic_vector(46, 8),
13542 => conv_std_logic_vector(46, 8),
13543 => conv_std_logic_vector(46, 8),
13544 => conv_std_logic_vector(47, 8),
13545 => conv_std_logic_vector(47, 8),
13546 => conv_std_logic_vector(47, 8),
13547 => conv_std_logic_vector(47, 8),
13548 => conv_std_logic_vector(47, 8),
13549 => conv_std_logic_vector(48, 8),
13550 => conv_std_logic_vector(48, 8),
13551 => conv_std_logic_vector(48, 8),
13552 => conv_std_logic_vector(48, 8),
13553 => conv_std_logic_vector(48, 8),
13554 => conv_std_logic_vector(49, 8),
13555 => conv_std_logic_vector(49, 8),
13556 => conv_std_logic_vector(49, 8),
13557 => conv_std_logic_vector(49, 8),
13558 => conv_std_logic_vector(49, 8),
13559 => conv_std_logic_vector(50, 8),
13560 => conv_std_logic_vector(50, 8),
13561 => conv_std_logic_vector(50, 8),
13562 => conv_std_logic_vector(50, 8),
13563 => conv_std_logic_vector(50, 8),
13564 => conv_std_logic_vector(51, 8),
13565 => conv_std_logic_vector(51, 8),
13566 => conv_std_logic_vector(51, 8),
13567 => conv_std_logic_vector(51, 8),
13568 => conv_std_logic_vector(0, 8),
13569 => conv_std_logic_vector(0, 8),
13570 => conv_std_logic_vector(0, 8),
13571 => conv_std_logic_vector(0, 8),
13572 => conv_std_logic_vector(0, 8),
13573 => conv_std_logic_vector(1, 8),
13574 => conv_std_logic_vector(1, 8),
13575 => conv_std_logic_vector(1, 8),
13576 => conv_std_logic_vector(1, 8),
13577 => conv_std_logic_vector(1, 8),
13578 => conv_std_logic_vector(2, 8),
13579 => conv_std_logic_vector(2, 8),
13580 => conv_std_logic_vector(2, 8),
13581 => conv_std_logic_vector(2, 8),
13582 => conv_std_logic_vector(2, 8),
13583 => conv_std_logic_vector(3, 8),
13584 => conv_std_logic_vector(3, 8),
13585 => conv_std_logic_vector(3, 8),
13586 => conv_std_logic_vector(3, 8),
13587 => conv_std_logic_vector(3, 8),
13588 => conv_std_logic_vector(4, 8),
13589 => conv_std_logic_vector(4, 8),
13590 => conv_std_logic_vector(4, 8),
13591 => conv_std_logic_vector(4, 8),
13592 => conv_std_logic_vector(4, 8),
13593 => conv_std_logic_vector(5, 8),
13594 => conv_std_logic_vector(5, 8),
13595 => conv_std_logic_vector(5, 8),
13596 => conv_std_logic_vector(5, 8),
13597 => conv_std_logic_vector(6, 8),
13598 => conv_std_logic_vector(6, 8),
13599 => conv_std_logic_vector(6, 8),
13600 => conv_std_logic_vector(6, 8),
13601 => conv_std_logic_vector(6, 8),
13602 => conv_std_logic_vector(7, 8),
13603 => conv_std_logic_vector(7, 8),
13604 => conv_std_logic_vector(7, 8),
13605 => conv_std_logic_vector(7, 8),
13606 => conv_std_logic_vector(7, 8),
13607 => conv_std_logic_vector(8, 8),
13608 => conv_std_logic_vector(8, 8),
13609 => conv_std_logic_vector(8, 8),
13610 => conv_std_logic_vector(8, 8),
13611 => conv_std_logic_vector(8, 8),
13612 => conv_std_logic_vector(9, 8),
13613 => conv_std_logic_vector(9, 8),
13614 => conv_std_logic_vector(9, 8),
13615 => conv_std_logic_vector(9, 8),
13616 => conv_std_logic_vector(9, 8),
13617 => conv_std_logic_vector(10, 8),
13618 => conv_std_logic_vector(10, 8),
13619 => conv_std_logic_vector(10, 8),
13620 => conv_std_logic_vector(10, 8),
13621 => conv_std_logic_vector(10, 8),
13622 => conv_std_logic_vector(11, 8),
13623 => conv_std_logic_vector(11, 8),
13624 => conv_std_logic_vector(11, 8),
13625 => conv_std_logic_vector(11, 8),
13626 => conv_std_logic_vector(12, 8),
13627 => conv_std_logic_vector(12, 8),
13628 => conv_std_logic_vector(12, 8),
13629 => conv_std_logic_vector(12, 8),
13630 => conv_std_logic_vector(12, 8),
13631 => conv_std_logic_vector(13, 8),
13632 => conv_std_logic_vector(13, 8),
13633 => conv_std_logic_vector(13, 8),
13634 => conv_std_logic_vector(13, 8),
13635 => conv_std_logic_vector(13, 8),
13636 => conv_std_logic_vector(14, 8),
13637 => conv_std_logic_vector(14, 8),
13638 => conv_std_logic_vector(14, 8),
13639 => conv_std_logic_vector(14, 8),
13640 => conv_std_logic_vector(14, 8),
13641 => conv_std_logic_vector(15, 8),
13642 => conv_std_logic_vector(15, 8),
13643 => conv_std_logic_vector(15, 8),
13644 => conv_std_logic_vector(15, 8),
13645 => conv_std_logic_vector(15, 8),
13646 => conv_std_logic_vector(16, 8),
13647 => conv_std_logic_vector(16, 8),
13648 => conv_std_logic_vector(16, 8),
13649 => conv_std_logic_vector(16, 8),
13650 => conv_std_logic_vector(16, 8),
13651 => conv_std_logic_vector(17, 8),
13652 => conv_std_logic_vector(17, 8),
13653 => conv_std_logic_vector(17, 8),
13654 => conv_std_logic_vector(17, 8),
13655 => conv_std_logic_vector(18, 8),
13656 => conv_std_logic_vector(18, 8),
13657 => conv_std_logic_vector(18, 8),
13658 => conv_std_logic_vector(18, 8),
13659 => conv_std_logic_vector(18, 8),
13660 => conv_std_logic_vector(19, 8),
13661 => conv_std_logic_vector(19, 8),
13662 => conv_std_logic_vector(19, 8),
13663 => conv_std_logic_vector(19, 8),
13664 => conv_std_logic_vector(19, 8),
13665 => conv_std_logic_vector(20, 8),
13666 => conv_std_logic_vector(20, 8),
13667 => conv_std_logic_vector(20, 8),
13668 => conv_std_logic_vector(20, 8),
13669 => conv_std_logic_vector(20, 8),
13670 => conv_std_logic_vector(21, 8),
13671 => conv_std_logic_vector(21, 8),
13672 => conv_std_logic_vector(21, 8),
13673 => conv_std_logic_vector(21, 8),
13674 => conv_std_logic_vector(21, 8),
13675 => conv_std_logic_vector(22, 8),
13676 => conv_std_logic_vector(22, 8),
13677 => conv_std_logic_vector(22, 8),
13678 => conv_std_logic_vector(22, 8),
13679 => conv_std_logic_vector(22, 8),
13680 => conv_std_logic_vector(23, 8),
13681 => conv_std_logic_vector(23, 8),
13682 => conv_std_logic_vector(23, 8),
13683 => conv_std_logic_vector(23, 8),
13684 => conv_std_logic_vector(24, 8),
13685 => conv_std_logic_vector(24, 8),
13686 => conv_std_logic_vector(24, 8),
13687 => conv_std_logic_vector(24, 8),
13688 => conv_std_logic_vector(24, 8),
13689 => conv_std_logic_vector(25, 8),
13690 => conv_std_logic_vector(25, 8),
13691 => conv_std_logic_vector(25, 8),
13692 => conv_std_logic_vector(25, 8),
13693 => conv_std_logic_vector(25, 8),
13694 => conv_std_logic_vector(26, 8),
13695 => conv_std_logic_vector(26, 8),
13696 => conv_std_logic_vector(26, 8),
13697 => conv_std_logic_vector(26, 8),
13698 => conv_std_logic_vector(26, 8),
13699 => conv_std_logic_vector(27, 8),
13700 => conv_std_logic_vector(27, 8),
13701 => conv_std_logic_vector(27, 8),
13702 => conv_std_logic_vector(27, 8),
13703 => conv_std_logic_vector(27, 8),
13704 => conv_std_logic_vector(28, 8),
13705 => conv_std_logic_vector(28, 8),
13706 => conv_std_logic_vector(28, 8),
13707 => conv_std_logic_vector(28, 8),
13708 => conv_std_logic_vector(28, 8),
13709 => conv_std_logic_vector(29, 8),
13710 => conv_std_logic_vector(29, 8),
13711 => conv_std_logic_vector(29, 8),
13712 => conv_std_logic_vector(29, 8),
13713 => conv_std_logic_vector(30, 8),
13714 => conv_std_logic_vector(30, 8),
13715 => conv_std_logic_vector(30, 8),
13716 => conv_std_logic_vector(30, 8),
13717 => conv_std_logic_vector(30, 8),
13718 => conv_std_logic_vector(31, 8),
13719 => conv_std_logic_vector(31, 8),
13720 => conv_std_logic_vector(31, 8),
13721 => conv_std_logic_vector(31, 8),
13722 => conv_std_logic_vector(31, 8),
13723 => conv_std_logic_vector(32, 8),
13724 => conv_std_logic_vector(32, 8),
13725 => conv_std_logic_vector(32, 8),
13726 => conv_std_logic_vector(32, 8),
13727 => conv_std_logic_vector(32, 8),
13728 => conv_std_logic_vector(33, 8),
13729 => conv_std_logic_vector(33, 8),
13730 => conv_std_logic_vector(33, 8),
13731 => conv_std_logic_vector(33, 8),
13732 => conv_std_logic_vector(33, 8),
13733 => conv_std_logic_vector(34, 8),
13734 => conv_std_logic_vector(34, 8),
13735 => conv_std_logic_vector(34, 8),
13736 => conv_std_logic_vector(34, 8),
13737 => conv_std_logic_vector(34, 8),
13738 => conv_std_logic_vector(35, 8),
13739 => conv_std_logic_vector(35, 8),
13740 => conv_std_logic_vector(35, 8),
13741 => conv_std_logic_vector(35, 8),
13742 => conv_std_logic_vector(36, 8),
13743 => conv_std_logic_vector(36, 8),
13744 => conv_std_logic_vector(36, 8),
13745 => conv_std_logic_vector(36, 8),
13746 => conv_std_logic_vector(36, 8),
13747 => conv_std_logic_vector(37, 8),
13748 => conv_std_logic_vector(37, 8),
13749 => conv_std_logic_vector(37, 8),
13750 => conv_std_logic_vector(37, 8),
13751 => conv_std_logic_vector(37, 8),
13752 => conv_std_logic_vector(38, 8),
13753 => conv_std_logic_vector(38, 8),
13754 => conv_std_logic_vector(38, 8),
13755 => conv_std_logic_vector(38, 8),
13756 => conv_std_logic_vector(38, 8),
13757 => conv_std_logic_vector(39, 8),
13758 => conv_std_logic_vector(39, 8),
13759 => conv_std_logic_vector(39, 8),
13760 => conv_std_logic_vector(39, 8),
13761 => conv_std_logic_vector(39, 8),
13762 => conv_std_logic_vector(40, 8),
13763 => conv_std_logic_vector(40, 8),
13764 => conv_std_logic_vector(40, 8),
13765 => conv_std_logic_vector(40, 8),
13766 => conv_std_logic_vector(40, 8),
13767 => conv_std_logic_vector(41, 8),
13768 => conv_std_logic_vector(41, 8),
13769 => conv_std_logic_vector(41, 8),
13770 => conv_std_logic_vector(41, 8),
13771 => conv_std_logic_vector(42, 8),
13772 => conv_std_logic_vector(42, 8),
13773 => conv_std_logic_vector(42, 8),
13774 => conv_std_logic_vector(42, 8),
13775 => conv_std_logic_vector(42, 8),
13776 => conv_std_logic_vector(43, 8),
13777 => conv_std_logic_vector(43, 8),
13778 => conv_std_logic_vector(43, 8),
13779 => conv_std_logic_vector(43, 8),
13780 => conv_std_logic_vector(43, 8),
13781 => conv_std_logic_vector(44, 8),
13782 => conv_std_logic_vector(44, 8),
13783 => conv_std_logic_vector(44, 8),
13784 => conv_std_logic_vector(44, 8),
13785 => conv_std_logic_vector(44, 8),
13786 => conv_std_logic_vector(45, 8),
13787 => conv_std_logic_vector(45, 8),
13788 => conv_std_logic_vector(45, 8),
13789 => conv_std_logic_vector(45, 8),
13790 => conv_std_logic_vector(45, 8),
13791 => conv_std_logic_vector(46, 8),
13792 => conv_std_logic_vector(46, 8),
13793 => conv_std_logic_vector(46, 8),
13794 => conv_std_logic_vector(46, 8),
13795 => conv_std_logic_vector(46, 8),
13796 => conv_std_logic_vector(47, 8),
13797 => conv_std_logic_vector(47, 8),
13798 => conv_std_logic_vector(47, 8),
13799 => conv_std_logic_vector(47, 8),
13800 => conv_std_logic_vector(48, 8),
13801 => conv_std_logic_vector(48, 8),
13802 => conv_std_logic_vector(48, 8),
13803 => conv_std_logic_vector(48, 8),
13804 => conv_std_logic_vector(48, 8),
13805 => conv_std_logic_vector(49, 8),
13806 => conv_std_logic_vector(49, 8),
13807 => conv_std_logic_vector(49, 8),
13808 => conv_std_logic_vector(49, 8),
13809 => conv_std_logic_vector(49, 8),
13810 => conv_std_logic_vector(50, 8),
13811 => conv_std_logic_vector(50, 8),
13812 => conv_std_logic_vector(50, 8),
13813 => conv_std_logic_vector(50, 8),
13814 => conv_std_logic_vector(50, 8),
13815 => conv_std_logic_vector(51, 8),
13816 => conv_std_logic_vector(51, 8),
13817 => conv_std_logic_vector(51, 8),
13818 => conv_std_logic_vector(51, 8),
13819 => conv_std_logic_vector(51, 8),
13820 => conv_std_logic_vector(52, 8),
13821 => conv_std_logic_vector(52, 8),
13822 => conv_std_logic_vector(52, 8),
13823 => conv_std_logic_vector(52, 8),
13824 => conv_std_logic_vector(0, 8),
13825 => conv_std_logic_vector(0, 8),
13826 => conv_std_logic_vector(0, 8),
13827 => conv_std_logic_vector(0, 8),
13828 => conv_std_logic_vector(0, 8),
13829 => conv_std_logic_vector(1, 8),
13830 => conv_std_logic_vector(1, 8),
13831 => conv_std_logic_vector(1, 8),
13832 => conv_std_logic_vector(1, 8),
13833 => conv_std_logic_vector(1, 8),
13834 => conv_std_logic_vector(2, 8),
13835 => conv_std_logic_vector(2, 8),
13836 => conv_std_logic_vector(2, 8),
13837 => conv_std_logic_vector(2, 8),
13838 => conv_std_logic_vector(2, 8),
13839 => conv_std_logic_vector(3, 8),
13840 => conv_std_logic_vector(3, 8),
13841 => conv_std_logic_vector(3, 8),
13842 => conv_std_logic_vector(3, 8),
13843 => conv_std_logic_vector(4, 8),
13844 => conv_std_logic_vector(4, 8),
13845 => conv_std_logic_vector(4, 8),
13846 => conv_std_logic_vector(4, 8),
13847 => conv_std_logic_vector(4, 8),
13848 => conv_std_logic_vector(5, 8),
13849 => conv_std_logic_vector(5, 8),
13850 => conv_std_logic_vector(5, 8),
13851 => conv_std_logic_vector(5, 8),
13852 => conv_std_logic_vector(5, 8),
13853 => conv_std_logic_vector(6, 8),
13854 => conv_std_logic_vector(6, 8),
13855 => conv_std_logic_vector(6, 8),
13856 => conv_std_logic_vector(6, 8),
13857 => conv_std_logic_vector(6, 8),
13858 => conv_std_logic_vector(7, 8),
13859 => conv_std_logic_vector(7, 8),
13860 => conv_std_logic_vector(7, 8),
13861 => conv_std_logic_vector(7, 8),
13862 => conv_std_logic_vector(8, 8),
13863 => conv_std_logic_vector(8, 8),
13864 => conv_std_logic_vector(8, 8),
13865 => conv_std_logic_vector(8, 8),
13866 => conv_std_logic_vector(8, 8),
13867 => conv_std_logic_vector(9, 8),
13868 => conv_std_logic_vector(9, 8),
13869 => conv_std_logic_vector(9, 8),
13870 => conv_std_logic_vector(9, 8),
13871 => conv_std_logic_vector(9, 8),
13872 => conv_std_logic_vector(10, 8),
13873 => conv_std_logic_vector(10, 8),
13874 => conv_std_logic_vector(10, 8),
13875 => conv_std_logic_vector(10, 8),
13876 => conv_std_logic_vector(10, 8),
13877 => conv_std_logic_vector(11, 8),
13878 => conv_std_logic_vector(11, 8),
13879 => conv_std_logic_vector(11, 8),
13880 => conv_std_logic_vector(11, 8),
13881 => conv_std_logic_vector(12, 8),
13882 => conv_std_logic_vector(12, 8),
13883 => conv_std_logic_vector(12, 8),
13884 => conv_std_logic_vector(12, 8),
13885 => conv_std_logic_vector(12, 8),
13886 => conv_std_logic_vector(13, 8),
13887 => conv_std_logic_vector(13, 8),
13888 => conv_std_logic_vector(13, 8),
13889 => conv_std_logic_vector(13, 8),
13890 => conv_std_logic_vector(13, 8),
13891 => conv_std_logic_vector(14, 8),
13892 => conv_std_logic_vector(14, 8),
13893 => conv_std_logic_vector(14, 8),
13894 => conv_std_logic_vector(14, 8),
13895 => conv_std_logic_vector(14, 8),
13896 => conv_std_logic_vector(15, 8),
13897 => conv_std_logic_vector(15, 8),
13898 => conv_std_logic_vector(15, 8),
13899 => conv_std_logic_vector(15, 8),
13900 => conv_std_logic_vector(16, 8),
13901 => conv_std_logic_vector(16, 8),
13902 => conv_std_logic_vector(16, 8),
13903 => conv_std_logic_vector(16, 8),
13904 => conv_std_logic_vector(16, 8),
13905 => conv_std_logic_vector(17, 8),
13906 => conv_std_logic_vector(17, 8),
13907 => conv_std_logic_vector(17, 8),
13908 => conv_std_logic_vector(17, 8),
13909 => conv_std_logic_vector(17, 8),
13910 => conv_std_logic_vector(18, 8),
13911 => conv_std_logic_vector(18, 8),
13912 => conv_std_logic_vector(18, 8),
13913 => conv_std_logic_vector(18, 8),
13914 => conv_std_logic_vector(18, 8),
13915 => conv_std_logic_vector(19, 8),
13916 => conv_std_logic_vector(19, 8),
13917 => conv_std_logic_vector(19, 8),
13918 => conv_std_logic_vector(19, 8),
13919 => conv_std_logic_vector(20, 8),
13920 => conv_std_logic_vector(20, 8),
13921 => conv_std_logic_vector(20, 8),
13922 => conv_std_logic_vector(20, 8),
13923 => conv_std_logic_vector(20, 8),
13924 => conv_std_logic_vector(21, 8),
13925 => conv_std_logic_vector(21, 8),
13926 => conv_std_logic_vector(21, 8),
13927 => conv_std_logic_vector(21, 8),
13928 => conv_std_logic_vector(21, 8),
13929 => conv_std_logic_vector(22, 8),
13930 => conv_std_logic_vector(22, 8),
13931 => conv_std_logic_vector(22, 8),
13932 => conv_std_logic_vector(22, 8),
13933 => conv_std_logic_vector(22, 8),
13934 => conv_std_logic_vector(23, 8),
13935 => conv_std_logic_vector(23, 8),
13936 => conv_std_logic_vector(23, 8),
13937 => conv_std_logic_vector(23, 8),
13938 => conv_std_logic_vector(24, 8),
13939 => conv_std_logic_vector(24, 8),
13940 => conv_std_logic_vector(24, 8),
13941 => conv_std_logic_vector(24, 8),
13942 => conv_std_logic_vector(24, 8),
13943 => conv_std_logic_vector(25, 8),
13944 => conv_std_logic_vector(25, 8),
13945 => conv_std_logic_vector(25, 8),
13946 => conv_std_logic_vector(25, 8),
13947 => conv_std_logic_vector(25, 8),
13948 => conv_std_logic_vector(26, 8),
13949 => conv_std_logic_vector(26, 8),
13950 => conv_std_logic_vector(26, 8),
13951 => conv_std_logic_vector(26, 8),
13952 => conv_std_logic_vector(27, 8),
13953 => conv_std_logic_vector(27, 8),
13954 => conv_std_logic_vector(27, 8),
13955 => conv_std_logic_vector(27, 8),
13956 => conv_std_logic_vector(27, 8),
13957 => conv_std_logic_vector(28, 8),
13958 => conv_std_logic_vector(28, 8),
13959 => conv_std_logic_vector(28, 8),
13960 => conv_std_logic_vector(28, 8),
13961 => conv_std_logic_vector(28, 8),
13962 => conv_std_logic_vector(29, 8),
13963 => conv_std_logic_vector(29, 8),
13964 => conv_std_logic_vector(29, 8),
13965 => conv_std_logic_vector(29, 8),
13966 => conv_std_logic_vector(29, 8),
13967 => conv_std_logic_vector(30, 8),
13968 => conv_std_logic_vector(30, 8),
13969 => conv_std_logic_vector(30, 8),
13970 => conv_std_logic_vector(30, 8),
13971 => conv_std_logic_vector(31, 8),
13972 => conv_std_logic_vector(31, 8),
13973 => conv_std_logic_vector(31, 8),
13974 => conv_std_logic_vector(31, 8),
13975 => conv_std_logic_vector(31, 8),
13976 => conv_std_logic_vector(32, 8),
13977 => conv_std_logic_vector(32, 8),
13978 => conv_std_logic_vector(32, 8),
13979 => conv_std_logic_vector(32, 8),
13980 => conv_std_logic_vector(32, 8),
13981 => conv_std_logic_vector(33, 8),
13982 => conv_std_logic_vector(33, 8),
13983 => conv_std_logic_vector(33, 8),
13984 => conv_std_logic_vector(33, 8),
13985 => conv_std_logic_vector(33, 8),
13986 => conv_std_logic_vector(34, 8),
13987 => conv_std_logic_vector(34, 8),
13988 => conv_std_logic_vector(34, 8),
13989 => conv_std_logic_vector(34, 8),
13990 => conv_std_logic_vector(35, 8),
13991 => conv_std_logic_vector(35, 8),
13992 => conv_std_logic_vector(35, 8),
13993 => conv_std_logic_vector(35, 8),
13994 => conv_std_logic_vector(35, 8),
13995 => conv_std_logic_vector(36, 8),
13996 => conv_std_logic_vector(36, 8),
13997 => conv_std_logic_vector(36, 8),
13998 => conv_std_logic_vector(36, 8),
13999 => conv_std_logic_vector(36, 8),
14000 => conv_std_logic_vector(37, 8),
14001 => conv_std_logic_vector(37, 8),
14002 => conv_std_logic_vector(37, 8),
14003 => conv_std_logic_vector(37, 8),
14004 => conv_std_logic_vector(37, 8),
14005 => conv_std_logic_vector(38, 8),
14006 => conv_std_logic_vector(38, 8),
14007 => conv_std_logic_vector(38, 8),
14008 => conv_std_logic_vector(38, 8),
14009 => conv_std_logic_vector(39, 8),
14010 => conv_std_logic_vector(39, 8),
14011 => conv_std_logic_vector(39, 8),
14012 => conv_std_logic_vector(39, 8),
14013 => conv_std_logic_vector(39, 8),
14014 => conv_std_logic_vector(40, 8),
14015 => conv_std_logic_vector(40, 8),
14016 => conv_std_logic_vector(40, 8),
14017 => conv_std_logic_vector(40, 8),
14018 => conv_std_logic_vector(40, 8),
14019 => conv_std_logic_vector(41, 8),
14020 => conv_std_logic_vector(41, 8),
14021 => conv_std_logic_vector(41, 8),
14022 => conv_std_logic_vector(41, 8),
14023 => conv_std_logic_vector(41, 8),
14024 => conv_std_logic_vector(42, 8),
14025 => conv_std_logic_vector(42, 8),
14026 => conv_std_logic_vector(42, 8),
14027 => conv_std_logic_vector(42, 8),
14028 => conv_std_logic_vector(43, 8),
14029 => conv_std_logic_vector(43, 8),
14030 => conv_std_logic_vector(43, 8),
14031 => conv_std_logic_vector(43, 8),
14032 => conv_std_logic_vector(43, 8),
14033 => conv_std_logic_vector(44, 8),
14034 => conv_std_logic_vector(44, 8),
14035 => conv_std_logic_vector(44, 8),
14036 => conv_std_logic_vector(44, 8),
14037 => conv_std_logic_vector(44, 8),
14038 => conv_std_logic_vector(45, 8),
14039 => conv_std_logic_vector(45, 8),
14040 => conv_std_logic_vector(45, 8),
14041 => conv_std_logic_vector(45, 8),
14042 => conv_std_logic_vector(45, 8),
14043 => conv_std_logic_vector(46, 8),
14044 => conv_std_logic_vector(46, 8),
14045 => conv_std_logic_vector(46, 8),
14046 => conv_std_logic_vector(46, 8),
14047 => conv_std_logic_vector(47, 8),
14048 => conv_std_logic_vector(47, 8),
14049 => conv_std_logic_vector(47, 8),
14050 => conv_std_logic_vector(47, 8),
14051 => conv_std_logic_vector(47, 8),
14052 => conv_std_logic_vector(48, 8),
14053 => conv_std_logic_vector(48, 8),
14054 => conv_std_logic_vector(48, 8),
14055 => conv_std_logic_vector(48, 8),
14056 => conv_std_logic_vector(48, 8),
14057 => conv_std_logic_vector(49, 8),
14058 => conv_std_logic_vector(49, 8),
14059 => conv_std_logic_vector(49, 8),
14060 => conv_std_logic_vector(49, 8),
14061 => conv_std_logic_vector(49, 8),
14062 => conv_std_logic_vector(50, 8),
14063 => conv_std_logic_vector(50, 8),
14064 => conv_std_logic_vector(50, 8),
14065 => conv_std_logic_vector(50, 8),
14066 => conv_std_logic_vector(51, 8),
14067 => conv_std_logic_vector(51, 8),
14068 => conv_std_logic_vector(51, 8),
14069 => conv_std_logic_vector(51, 8),
14070 => conv_std_logic_vector(51, 8),
14071 => conv_std_logic_vector(52, 8),
14072 => conv_std_logic_vector(52, 8),
14073 => conv_std_logic_vector(52, 8),
14074 => conv_std_logic_vector(52, 8),
14075 => conv_std_logic_vector(52, 8),
14076 => conv_std_logic_vector(53, 8),
14077 => conv_std_logic_vector(53, 8),
14078 => conv_std_logic_vector(53, 8),
14079 => conv_std_logic_vector(53, 8),
14080 => conv_std_logic_vector(0, 8),
14081 => conv_std_logic_vector(0, 8),
14082 => conv_std_logic_vector(0, 8),
14083 => conv_std_logic_vector(0, 8),
14084 => conv_std_logic_vector(0, 8),
14085 => conv_std_logic_vector(1, 8),
14086 => conv_std_logic_vector(1, 8),
14087 => conv_std_logic_vector(1, 8),
14088 => conv_std_logic_vector(1, 8),
14089 => conv_std_logic_vector(1, 8),
14090 => conv_std_logic_vector(2, 8),
14091 => conv_std_logic_vector(2, 8),
14092 => conv_std_logic_vector(2, 8),
14093 => conv_std_logic_vector(2, 8),
14094 => conv_std_logic_vector(3, 8),
14095 => conv_std_logic_vector(3, 8),
14096 => conv_std_logic_vector(3, 8),
14097 => conv_std_logic_vector(3, 8),
14098 => conv_std_logic_vector(3, 8),
14099 => conv_std_logic_vector(4, 8),
14100 => conv_std_logic_vector(4, 8),
14101 => conv_std_logic_vector(4, 8),
14102 => conv_std_logic_vector(4, 8),
14103 => conv_std_logic_vector(4, 8),
14104 => conv_std_logic_vector(5, 8),
14105 => conv_std_logic_vector(5, 8),
14106 => conv_std_logic_vector(5, 8),
14107 => conv_std_logic_vector(5, 8),
14108 => conv_std_logic_vector(6, 8),
14109 => conv_std_logic_vector(6, 8),
14110 => conv_std_logic_vector(6, 8),
14111 => conv_std_logic_vector(6, 8),
14112 => conv_std_logic_vector(6, 8),
14113 => conv_std_logic_vector(7, 8),
14114 => conv_std_logic_vector(7, 8),
14115 => conv_std_logic_vector(7, 8),
14116 => conv_std_logic_vector(7, 8),
14117 => conv_std_logic_vector(7, 8),
14118 => conv_std_logic_vector(8, 8),
14119 => conv_std_logic_vector(8, 8),
14120 => conv_std_logic_vector(8, 8),
14121 => conv_std_logic_vector(8, 8),
14122 => conv_std_logic_vector(9, 8),
14123 => conv_std_logic_vector(9, 8),
14124 => conv_std_logic_vector(9, 8),
14125 => conv_std_logic_vector(9, 8),
14126 => conv_std_logic_vector(9, 8),
14127 => conv_std_logic_vector(10, 8),
14128 => conv_std_logic_vector(10, 8),
14129 => conv_std_logic_vector(10, 8),
14130 => conv_std_logic_vector(10, 8),
14131 => conv_std_logic_vector(10, 8),
14132 => conv_std_logic_vector(11, 8),
14133 => conv_std_logic_vector(11, 8),
14134 => conv_std_logic_vector(11, 8),
14135 => conv_std_logic_vector(11, 8),
14136 => conv_std_logic_vector(12, 8),
14137 => conv_std_logic_vector(12, 8),
14138 => conv_std_logic_vector(12, 8),
14139 => conv_std_logic_vector(12, 8),
14140 => conv_std_logic_vector(12, 8),
14141 => conv_std_logic_vector(13, 8),
14142 => conv_std_logic_vector(13, 8),
14143 => conv_std_logic_vector(13, 8),
14144 => conv_std_logic_vector(13, 8),
14145 => conv_std_logic_vector(13, 8),
14146 => conv_std_logic_vector(14, 8),
14147 => conv_std_logic_vector(14, 8),
14148 => conv_std_logic_vector(14, 8),
14149 => conv_std_logic_vector(14, 8),
14150 => conv_std_logic_vector(15, 8),
14151 => conv_std_logic_vector(15, 8),
14152 => conv_std_logic_vector(15, 8),
14153 => conv_std_logic_vector(15, 8),
14154 => conv_std_logic_vector(15, 8),
14155 => conv_std_logic_vector(16, 8),
14156 => conv_std_logic_vector(16, 8),
14157 => conv_std_logic_vector(16, 8),
14158 => conv_std_logic_vector(16, 8),
14159 => conv_std_logic_vector(16, 8),
14160 => conv_std_logic_vector(17, 8),
14161 => conv_std_logic_vector(17, 8),
14162 => conv_std_logic_vector(17, 8),
14163 => conv_std_logic_vector(17, 8),
14164 => conv_std_logic_vector(18, 8),
14165 => conv_std_logic_vector(18, 8),
14166 => conv_std_logic_vector(18, 8),
14167 => conv_std_logic_vector(18, 8),
14168 => conv_std_logic_vector(18, 8),
14169 => conv_std_logic_vector(19, 8),
14170 => conv_std_logic_vector(19, 8),
14171 => conv_std_logic_vector(19, 8),
14172 => conv_std_logic_vector(19, 8),
14173 => conv_std_logic_vector(19, 8),
14174 => conv_std_logic_vector(20, 8),
14175 => conv_std_logic_vector(20, 8),
14176 => conv_std_logic_vector(20, 8),
14177 => conv_std_logic_vector(20, 8),
14178 => conv_std_logic_vector(21, 8),
14179 => conv_std_logic_vector(21, 8),
14180 => conv_std_logic_vector(21, 8),
14181 => conv_std_logic_vector(21, 8),
14182 => conv_std_logic_vector(21, 8),
14183 => conv_std_logic_vector(22, 8),
14184 => conv_std_logic_vector(22, 8),
14185 => conv_std_logic_vector(22, 8),
14186 => conv_std_logic_vector(22, 8),
14187 => conv_std_logic_vector(22, 8),
14188 => conv_std_logic_vector(23, 8),
14189 => conv_std_logic_vector(23, 8),
14190 => conv_std_logic_vector(23, 8),
14191 => conv_std_logic_vector(23, 8),
14192 => conv_std_logic_vector(24, 8),
14193 => conv_std_logic_vector(24, 8),
14194 => conv_std_logic_vector(24, 8),
14195 => conv_std_logic_vector(24, 8),
14196 => conv_std_logic_vector(24, 8),
14197 => conv_std_logic_vector(25, 8),
14198 => conv_std_logic_vector(25, 8),
14199 => conv_std_logic_vector(25, 8),
14200 => conv_std_logic_vector(25, 8),
14201 => conv_std_logic_vector(25, 8),
14202 => conv_std_logic_vector(26, 8),
14203 => conv_std_logic_vector(26, 8),
14204 => conv_std_logic_vector(26, 8),
14205 => conv_std_logic_vector(26, 8),
14206 => conv_std_logic_vector(27, 8),
14207 => conv_std_logic_vector(27, 8),
14208 => conv_std_logic_vector(27, 8),
14209 => conv_std_logic_vector(27, 8),
14210 => conv_std_logic_vector(27, 8),
14211 => conv_std_logic_vector(28, 8),
14212 => conv_std_logic_vector(28, 8),
14213 => conv_std_logic_vector(28, 8),
14214 => conv_std_logic_vector(28, 8),
14215 => conv_std_logic_vector(29, 8),
14216 => conv_std_logic_vector(29, 8),
14217 => conv_std_logic_vector(29, 8),
14218 => conv_std_logic_vector(29, 8),
14219 => conv_std_logic_vector(29, 8),
14220 => conv_std_logic_vector(30, 8),
14221 => conv_std_logic_vector(30, 8),
14222 => conv_std_logic_vector(30, 8),
14223 => conv_std_logic_vector(30, 8),
14224 => conv_std_logic_vector(30, 8),
14225 => conv_std_logic_vector(31, 8),
14226 => conv_std_logic_vector(31, 8),
14227 => conv_std_logic_vector(31, 8),
14228 => conv_std_logic_vector(31, 8),
14229 => conv_std_logic_vector(32, 8),
14230 => conv_std_logic_vector(32, 8),
14231 => conv_std_logic_vector(32, 8),
14232 => conv_std_logic_vector(32, 8),
14233 => conv_std_logic_vector(32, 8),
14234 => conv_std_logic_vector(33, 8),
14235 => conv_std_logic_vector(33, 8),
14236 => conv_std_logic_vector(33, 8),
14237 => conv_std_logic_vector(33, 8),
14238 => conv_std_logic_vector(33, 8),
14239 => conv_std_logic_vector(34, 8),
14240 => conv_std_logic_vector(34, 8),
14241 => conv_std_logic_vector(34, 8),
14242 => conv_std_logic_vector(34, 8),
14243 => conv_std_logic_vector(35, 8),
14244 => conv_std_logic_vector(35, 8),
14245 => conv_std_logic_vector(35, 8),
14246 => conv_std_logic_vector(35, 8),
14247 => conv_std_logic_vector(35, 8),
14248 => conv_std_logic_vector(36, 8),
14249 => conv_std_logic_vector(36, 8),
14250 => conv_std_logic_vector(36, 8),
14251 => conv_std_logic_vector(36, 8),
14252 => conv_std_logic_vector(36, 8),
14253 => conv_std_logic_vector(37, 8),
14254 => conv_std_logic_vector(37, 8),
14255 => conv_std_logic_vector(37, 8),
14256 => conv_std_logic_vector(37, 8),
14257 => conv_std_logic_vector(38, 8),
14258 => conv_std_logic_vector(38, 8),
14259 => conv_std_logic_vector(38, 8),
14260 => conv_std_logic_vector(38, 8),
14261 => conv_std_logic_vector(38, 8),
14262 => conv_std_logic_vector(39, 8),
14263 => conv_std_logic_vector(39, 8),
14264 => conv_std_logic_vector(39, 8),
14265 => conv_std_logic_vector(39, 8),
14266 => conv_std_logic_vector(39, 8),
14267 => conv_std_logic_vector(40, 8),
14268 => conv_std_logic_vector(40, 8),
14269 => conv_std_logic_vector(40, 8),
14270 => conv_std_logic_vector(40, 8),
14271 => conv_std_logic_vector(41, 8),
14272 => conv_std_logic_vector(41, 8),
14273 => conv_std_logic_vector(41, 8),
14274 => conv_std_logic_vector(41, 8),
14275 => conv_std_logic_vector(41, 8),
14276 => conv_std_logic_vector(42, 8),
14277 => conv_std_logic_vector(42, 8),
14278 => conv_std_logic_vector(42, 8),
14279 => conv_std_logic_vector(42, 8),
14280 => conv_std_logic_vector(42, 8),
14281 => conv_std_logic_vector(43, 8),
14282 => conv_std_logic_vector(43, 8),
14283 => conv_std_logic_vector(43, 8),
14284 => conv_std_logic_vector(43, 8),
14285 => conv_std_logic_vector(44, 8),
14286 => conv_std_logic_vector(44, 8),
14287 => conv_std_logic_vector(44, 8),
14288 => conv_std_logic_vector(44, 8),
14289 => conv_std_logic_vector(44, 8),
14290 => conv_std_logic_vector(45, 8),
14291 => conv_std_logic_vector(45, 8),
14292 => conv_std_logic_vector(45, 8),
14293 => conv_std_logic_vector(45, 8),
14294 => conv_std_logic_vector(45, 8),
14295 => conv_std_logic_vector(46, 8),
14296 => conv_std_logic_vector(46, 8),
14297 => conv_std_logic_vector(46, 8),
14298 => conv_std_logic_vector(46, 8),
14299 => conv_std_logic_vector(47, 8),
14300 => conv_std_logic_vector(47, 8),
14301 => conv_std_logic_vector(47, 8),
14302 => conv_std_logic_vector(47, 8),
14303 => conv_std_logic_vector(47, 8),
14304 => conv_std_logic_vector(48, 8),
14305 => conv_std_logic_vector(48, 8),
14306 => conv_std_logic_vector(48, 8),
14307 => conv_std_logic_vector(48, 8),
14308 => conv_std_logic_vector(48, 8),
14309 => conv_std_logic_vector(49, 8),
14310 => conv_std_logic_vector(49, 8),
14311 => conv_std_logic_vector(49, 8),
14312 => conv_std_logic_vector(49, 8),
14313 => conv_std_logic_vector(50, 8),
14314 => conv_std_logic_vector(50, 8),
14315 => conv_std_logic_vector(50, 8),
14316 => conv_std_logic_vector(50, 8),
14317 => conv_std_logic_vector(50, 8),
14318 => conv_std_logic_vector(51, 8),
14319 => conv_std_logic_vector(51, 8),
14320 => conv_std_logic_vector(51, 8),
14321 => conv_std_logic_vector(51, 8),
14322 => conv_std_logic_vector(51, 8),
14323 => conv_std_logic_vector(52, 8),
14324 => conv_std_logic_vector(52, 8),
14325 => conv_std_logic_vector(52, 8),
14326 => conv_std_logic_vector(52, 8),
14327 => conv_std_logic_vector(53, 8),
14328 => conv_std_logic_vector(53, 8),
14329 => conv_std_logic_vector(53, 8),
14330 => conv_std_logic_vector(53, 8),
14331 => conv_std_logic_vector(53, 8),
14332 => conv_std_logic_vector(54, 8),
14333 => conv_std_logic_vector(54, 8),
14334 => conv_std_logic_vector(54, 8),
14335 => conv_std_logic_vector(54, 8),
14336 => conv_std_logic_vector(0, 8),
14337 => conv_std_logic_vector(0, 8),
14338 => conv_std_logic_vector(0, 8),
14339 => conv_std_logic_vector(0, 8),
14340 => conv_std_logic_vector(0, 8),
14341 => conv_std_logic_vector(1, 8),
14342 => conv_std_logic_vector(1, 8),
14343 => conv_std_logic_vector(1, 8),
14344 => conv_std_logic_vector(1, 8),
14345 => conv_std_logic_vector(1, 8),
14346 => conv_std_logic_vector(2, 8),
14347 => conv_std_logic_vector(2, 8),
14348 => conv_std_logic_vector(2, 8),
14349 => conv_std_logic_vector(2, 8),
14350 => conv_std_logic_vector(3, 8),
14351 => conv_std_logic_vector(3, 8),
14352 => conv_std_logic_vector(3, 8),
14353 => conv_std_logic_vector(3, 8),
14354 => conv_std_logic_vector(3, 8),
14355 => conv_std_logic_vector(4, 8),
14356 => conv_std_logic_vector(4, 8),
14357 => conv_std_logic_vector(4, 8),
14358 => conv_std_logic_vector(4, 8),
14359 => conv_std_logic_vector(5, 8),
14360 => conv_std_logic_vector(5, 8),
14361 => conv_std_logic_vector(5, 8),
14362 => conv_std_logic_vector(5, 8),
14363 => conv_std_logic_vector(5, 8),
14364 => conv_std_logic_vector(6, 8),
14365 => conv_std_logic_vector(6, 8),
14366 => conv_std_logic_vector(6, 8),
14367 => conv_std_logic_vector(6, 8),
14368 => conv_std_logic_vector(7, 8),
14369 => conv_std_logic_vector(7, 8),
14370 => conv_std_logic_vector(7, 8),
14371 => conv_std_logic_vector(7, 8),
14372 => conv_std_logic_vector(7, 8),
14373 => conv_std_logic_vector(8, 8),
14374 => conv_std_logic_vector(8, 8),
14375 => conv_std_logic_vector(8, 8),
14376 => conv_std_logic_vector(8, 8),
14377 => conv_std_logic_vector(8, 8),
14378 => conv_std_logic_vector(9, 8),
14379 => conv_std_logic_vector(9, 8),
14380 => conv_std_logic_vector(9, 8),
14381 => conv_std_logic_vector(9, 8),
14382 => conv_std_logic_vector(10, 8),
14383 => conv_std_logic_vector(10, 8),
14384 => conv_std_logic_vector(10, 8),
14385 => conv_std_logic_vector(10, 8),
14386 => conv_std_logic_vector(10, 8),
14387 => conv_std_logic_vector(11, 8),
14388 => conv_std_logic_vector(11, 8),
14389 => conv_std_logic_vector(11, 8),
14390 => conv_std_logic_vector(11, 8),
14391 => conv_std_logic_vector(12, 8),
14392 => conv_std_logic_vector(12, 8),
14393 => conv_std_logic_vector(12, 8),
14394 => conv_std_logic_vector(12, 8),
14395 => conv_std_logic_vector(12, 8),
14396 => conv_std_logic_vector(13, 8),
14397 => conv_std_logic_vector(13, 8),
14398 => conv_std_logic_vector(13, 8),
14399 => conv_std_logic_vector(13, 8),
14400 => conv_std_logic_vector(14, 8),
14401 => conv_std_logic_vector(14, 8),
14402 => conv_std_logic_vector(14, 8),
14403 => conv_std_logic_vector(14, 8),
14404 => conv_std_logic_vector(14, 8),
14405 => conv_std_logic_vector(15, 8),
14406 => conv_std_logic_vector(15, 8),
14407 => conv_std_logic_vector(15, 8),
14408 => conv_std_logic_vector(15, 8),
14409 => conv_std_logic_vector(15, 8),
14410 => conv_std_logic_vector(16, 8),
14411 => conv_std_logic_vector(16, 8),
14412 => conv_std_logic_vector(16, 8),
14413 => conv_std_logic_vector(16, 8),
14414 => conv_std_logic_vector(17, 8),
14415 => conv_std_logic_vector(17, 8),
14416 => conv_std_logic_vector(17, 8),
14417 => conv_std_logic_vector(17, 8),
14418 => conv_std_logic_vector(17, 8),
14419 => conv_std_logic_vector(18, 8),
14420 => conv_std_logic_vector(18, 8),
14421 => conv_std_logic_vector(18, 8),
14422 => conv_std_logic_vector(18, 8),
14423 => conv_std_logic_vector(19, 8),
14424 => conv_std_logic_vector(19, 8),
14425 => conv_std_logic_vector(19, 8),
14426 => conv_std_logic_vector(19, 8),
14427 => conv_std_logic_vector(19, 8),
14428 => conv_std_logic_vector(20, 8),
14429 => conv_std_logic_vector(20, 8),
14430 => conv_std_logic_vector(20, 8),
14431 => conv_std_logic_vector(20, 8),
14432 => conv_std_logic_vector(21, 8),
14433 => conv_std_logic_vector(21, 8),
14434 => conv_std_logic_vector(21, 8),
14435 => conv_std_logic_vector(21, 8),
14436 => conv_std_logic_vector(21, 8),
14437 => conv_std_logic_vector(22, 8),
14438 => conv_std_logic_vector(22, 8),
14439 => conv_std_logic_vector(22, 8),
14440 => conv_std_logic_vector(22, 8),
14441 => conv_std_logic_vector(22, 8),
14442 => conv_std_logic_vector(23, 8),
14443 => conv_std_logic_vector(23, 8),
14444 => conv_std_logic_vector(23, 8),
14445 => conv_std_logic_vector(23, 8),
14446 => conv_std_logic_vector(24, 8),
14447 => conv_std_logic_vector(24, 8),
14448 => conv_std_logic_vector(24, 8),
14449 => conv_std_logic_vector(24, 8),
14450 => conv_std_logic_vector(24, 8),
14451 => conv_std_logic_vector(25, 8),
14452 => conv_std_logic_vector(25, 8),
14453 => conv_std_logic_vector(25, 8),
14454 => conv_std_logic_vector(25, 8),
14455 => conv_std_logic_vector(26, 8),
14456 => conv_std_logic_vector(26, 8),
14457 => conv_std_logic_vector(26, 8),
14458 => conv_std_logic_vector(26, 8),
14459 => conv_std_logic_vector(26, 8),
14460 => conv_std_logic_vector(27, 8),
14461 => conv_std_logic_vector(27, 8),
14462 => conv_std_logic_vector(27, 8),
14463 => conv_std_logic_vector(27, 8),
14464 => conv_std_logic_vector(28, 8),
14465 => conv_std_logic_vector(28, 8),
14466 => conv_std_logic_vector(28, 8),
14467 => conv_std_logic_vector(28, 8),
14468 => conv_std_logic_vector(28, 8),
14469 => conv_std_logic_vector(29, 8),
14470 => conv_std_logic_vector(29, 8),
14471 => conv_std_logic_vector(29, 8),
14472 => conv_std_logic_vector(29, 8),
14473 => conv_std_logic_vector(29, 8),
14474 => conv_std_logic_vector(30, 8),
14475 => conv_std_logic_vector(30, 8),
14476 => conv_std_logic_vector(30, 8),
14477 => conv_std_logic_vector(30, 8),
14478 => conv_std_logic_vector(31, 8),
14479 => conv_std_logic_vector(31, 8),
14480 => conv_std_logic_vector(31, 8),
14481 => conv_std_logic_vector(31, 8),
14482 => conv_std_logic_vector(31, 8),
14483 => conv_std_logic_vector(32, 8),
14484 => conv_std_logic_vector(32, 8),
14485 => conv_std_logic_vector(32, 8),
14486 => conv_std_logic_vector(32, 8),
14487 => conv_std_logic_vector(33, 8),
14488 => conv_std_logic_vector(33, 8),
14489 => conv_std_logic_vector(33, 8),
14490 => conv_std_logic_vector(33, 8),
14491 => conv_std_logic_vector(33, 8),
14492 => conv_std_logic_vector(34, 8),
14493 => conv_std_logic_vector(34, 8),
14494 => conv_std_logic_vector(34, 8),
14495 => conv_std_logic_vector(34, 8),
14496 => conv_std_logic_vector(35, 8),
14497 => conv_std_logic_vector(35, 8),
14498 => conv_std_logic_vector(35, 8),
14499 => conv_std_logic_vector(35, 8),
14500 => conv_std_logic_vector(35, 8),
14501 => conv_std_logic_vector(36, 8),
14502 => conv_std_logic_vector(36, 8),
14503 => conv_std_logic_vector(36, 8),
14504 => conv_std_logic_vector(36, 8),
14505 => conv_std_logic_vector(36, 8),
14506 => conv_std_logic_vector(37, 8),
14507 => conv_std_logic_vector(37, 8),
14508 => conv_std_logic_vector(37, 8),
14509 => conv_std_logic_vector(37, 8),
14510 => conv_std_logic_vector(38, 8),
14511 => conv_std_logic_vector(38, 8),
14512 => conv_std_logic_vector(38, 8),
14513 => conv_std_logic_vector(38, 8),
14514 => conv_std_logic_vector(38, 8),
14515 => conv_std_logic_vector(39, 8),
14516 => conv_std_logic_vector(39, 8),
14517 => conv_std_logic_vector(39, 8),
14518 => conv_std_logic_vector(39, 8),
14519 => conv_std_logic_vector(40, 8),
14520 => conv_std_logic_vector(40, 8),
14521 => conv_std_logic_vector(40, 8),
14522 => conv_std_logic_vector(40, 8),
14523 => conv_std_logic_vector(40, 8),
14524 => conv_std_logic_vector(41, 8),
14525 => conv_std_logic_vector(41, 8),
14526 => conv_std_logic_vector(41, 8),
14527 => conv_std_logic_vector(41, 8),
14528 => conv_std_logic_vector(42, 8),
14529 => conv_std_logic_vector(42, 8),
14530 => conv_std_logic_vector(42, 8),
14531 => conv_std_logic_vector(42, 8),
14532 => conv_std_logic_vector(42, 8),
14533 => conv_std_logic_vector(43, 8),
14534 => conv_std_logic_vector(43, 8),
14535 => conv_std_logic_vector(43, 8),
14536 => conv_std_logic_vector(43, 8),
14537 => conv_std_logic_vector(43, 8),
14538 => conv_std_logic_vector(44, 8),
14539 => conv_std_logic_vector(44, 8),
14540 => conv_std_logic_vector(44, 8),
14541 => conv_std_logic_vector(44, 8),
14542 => conv_std_logic_vector(45, 8),
14543 => conv_std_logic_vector(45, 8),
14544 => conv_std_logic_vector(45, 8),
14545 => conv_std_logic_vector(45, 8),
14546 => conv_std_logic_vector(45, 8),
14547 => conv_std_logic_vector(46, 8),
14548 => conv_std_logic_vector(46, 8),
14549 => conv_std_logic_vector(46, 8),
14550 => conv_std_logic_vector(46, 8),
14551 => conv_std_logic_vector(47, 8),
14552 => conv_std_logic_vector(47, 8),
14553 => conv_std_logic_vector(47, 8),
14554 => conv_std_logic_vector(47, 8),
14555 => conv_std_logic_vector(47, 8),
14556 => conv_std_logic_vector(48, 8),
14557 => conv_std_logic_vector(48, 8),
14558 => conv_std_logic_vector(48, 8),
14559 => conv_std_logic_vector(48, 8),
14560 => conv_std_logic_vector(49, 8),
14561 => conv_std_logic_vector(49, 8),
14562 => conv_std_logic_vector(49, 8),
14563 => conv_std_logic_vector(49, 8),
14564 => conv_std_logic_vector(49, 8),
14565 => conv_std_logic_vector(50, 8),
14566 => conv_std_logic_vector(50, 8),
14567 => conv_std_logic_vector(50, 8),
14568 => conv_std_logic_vector(50, 8),
14569 => conv_std_logic_vector(50, 8),
14570 => conv_std_logic_vector(51, 8),
14571 => conv_std_logic_vector(51, 8),
14572 => conv_std_logic_vector(51, 8),
14573 => conv_std_logic_vector(51, 8),
14574 => conv_std_logic_vector(52, 8),
14575 => conv_std_logic_vector(52, 8),
14576 => conv_std_logic_vector(52, 8),
14577 => conv_std_logic_vector(52, 8),
14578 => conv_std_logic_vector(52, 8),
14579 => conv_std_logic_vector(53, 8),
14580 => conv_std_logic_vector(53, 8),
14581 => conv_std_logic_vector(53, 8),
14582 => conv_std_logic_vector(53, 8),
14583 => conv_std_logic_vector(54, 8),
14584 => conv_std_logic_vector(54, 8),
14585 => conv_std_logic_vector(54, 8),
14586 => conv_std_logic_vector(54, 8),
14587 => conv_std_logic_vector(54, 8),
14588 => conv_std_logic_vector(55, 8),
14589 => conv_std_logic_vector(55, 8),
14590 => conv_std_logic_vector(55, 8),
14591 => conv_std_logic_vector(55, 8),
14592 => conv_std_logic_vector(0, 8),
14593 => conv_std_logic_vector(0, 8),
14594 => conv_std_logic_vector(0, 8),
14595 => conv_std_logic_vector(0, 8),
14596 => conv_std_logic_vector(0, 8),
14597 => conv_std_logic_vector(1, 8),
14598 => conv_std_logic_vector(1, 8),
14599 => conv_std_logic_vector(1, 8),
14600 => conv_std_logic_vector(1, 8),
14601 => conv_std_logic_vector(2, 8),
14602 => conv_std_logic_vector(2, 8),
14603 => conv_std_logic_vector(2, 8),
14604 => conv_std_logic_vector(2, 8),
14605 => conv_std_logic_vector(2, 8),
14606 => conv_std_logic_vector(3, 8),
14607 => conv_std_logic_vector(3, 8),
14608 => conv_std_logic_vector(3, 8),
14609 => conv_std_logic_vector(3, 8),
14610 => conv_std_logic_vector(4, 8),
14611 => conv_std_logic_vector(4, 8),
14612 => conv_std_logic_vector(4, 8),
14613 => conv_std_logic_vector(4, 8),
14614 => conv_std_logic_vector(4, 8),
14615 => conv_std_logic_vector(5, 8),
14616 => conv_std_logic_vector(5, 8),
14617 => conv_std_logic_vector(5, 8),
14618 => conv_std_logic_vector(5, 8),
14619 => conv_std_logic_vector(6, 8),
14620 => conv_std_logic_vector(6, 8),
14621 => conv_std_logic_vector(6, 8),
14622 => conv_std_logic_vector(6, 8),
14623 => conv_std_logic_vector(6, 8),
14624 => conv_std_logic_vector(7, 8),
14625 => conv_std_logic_vector(7, 8),
14626 => conv_std_logic_vector(7, 8),
14627 => conv_std_logic_vector(7, 8),
14628 => conv_std_logic_vector(8, 8),
14629 => conv_std_logic_vector(8, 8),
14630 => conv_std_logic_vector(8, 8),
14631 => conv_std_logic_vector(8, 8),
14632 => conv_std_logic_vector(8, 8),
14633 => conv_std_logic_vector(9, 8),
14634 => conv_std_logic_vector(9, 8),
14635 => conv_std_logic_vector(9, 8),
14636 => conv_std_logic_vector(9, 8),
14637 => conv_std_logic_vector(10, 8),
14638 => conv_std_logic_vector(10, 8),
14639 => conv_std_logic_vector(10, 8),
14640 => conv_std_logic_vector(10, 8),
14641 => conv_std_logic_vector(10, 8),
14642 => conv_std_logic_vector(11, 8),
14643 => conv_std_logic_vector(11, 8),
14644 => conv_std_logic_vector(11, 8),
14645 => conv_std_logic_vector(11, 8),
14646 => conv_std_logic_vector(12, 8),
14647 => conv_std_logic_vector(12, 8),
14648 => conv_std_logic_vector(12, 8),
14649 => conv_std_logic_vector(12, 8),
14650 => conv_std_logic_vector(12, 8),
14651 => conv_std_logic_vector(13, 8),
14652 => conv_std_logic_vector(13, 8),
14653 => conv_std_logic_vector(13, 8),
14654 => conv_std_logic_vector(13, 8),
14655 => conv_std_logic_vector(14, 8),
14656 => conv_std_logic_vector(14, 8),
14657 => conv_std_logic_vector(14, 8),
14658 => conv_std_logic_vector(14, 8),
14659 => conv_std_logic_vector(14, 8),
14660 => conv_std_logic_vector(15, 8),
14661 => conv_std_logic_vector(15, 8),
14662 => conv_std_logic_vector(15, 8),
14663 => conv_std_logic_vector(15, 8),
14664 => conv_std_logic_vector(16, 8),
14665 => conv_std_logic_vector(16, 8),
14666 => conv_std_logic_vector(16, 8),
14667 => conv_std_logic_vector(16, 8),
14668 => conv_std_logic_vector(16, 8),
14669 => conv_std_logic_vector(17, 8),
14670 => conv_std_logic_vector(17, 8),
14671 => conv_std_logic_vector(17, 8),
14672 => conv_std_logic_vector(17, 8),
14673 => conv_std_logic_vector(18, 8),
14674 => conv_std_logic_vector(18, 8),
14675 => conv_std_logic_vector(18, 8),
14676 => conv_std_logic_vector(18, 8),
14677 => conv_std_logic_vector(18, 8),
14678 => conv_std_logic_vector(19, 8),
14679 => conv_std_logic_vector(19, 8),
14680 => conv_std_logic_vector(19, 8),
14681 => conv_std_logic_vector(19, 8),
14682 => conv_std_logic_vector(20, 8),
14683 => conv_std_logic_vector(20, 8),
14684 => conv_std_logic_vector(20, 8),
14685 => conv_std_logic_vector(20, 8),
14686 => conv_std_logic_vector(20, 8),
14687 => conv_std_logic_vector(21, 8),
14688 => conv_std_logic_vector(21, 8),
14689 => conv_std_logic_vector(21, 8),
14690 => conv_std_logic_vector(21, 8),
14691 => conv_std_logic_vector(22, 8),
14692 => conv_std_logic_vector(22, 8),
14693 => conv_std_logic_vector(22, 8),
14694 => conv_std_logic_vector(22, 8),
14695 => conv_std_logic_vector(22, 8),
14696 => conv_std_logic_vector(23, 8),
14697 => conv_std_logic_vector(23, 8),
14698 => conv_std_logic_vector(23, 8),
14699 => conv_std_logic_vector(23, 8),
14700 => conv_std_logic_vector(24, 8),
14701 => conv_std_logic_vector(24, 8),
14702 => conv_std_logic_vector(24, 8),
14703 => conv_std_logic_vector(24, 8),
14704 => conv_std_logic_vector(24, 8),
14705 => conv_std_logic_vector(25, 8),
14706 => conv_std_logic_vector(25, 8),
14707 => conv_std_logic_vector(25, 8),
14708 => conv_std_logic_vector(25, 8),
14709 => conv_std_logic_vector(26, 8),
14710 => conv_std_logic_vector(26, 8),
14711 => conv_std_logic_vector(26, 8),
14712 => conv_std_logic_vector(26, 8),
14713 => conv_std_logic_vector(26, 8),
14714 => conv_std_logic_vector(27, 8),
14715 => conv_std_logic_vector(27, 8),
14716 => conv_std_logic_vector(27, 8),
14717 => conv_std_logic_vector(27, 8),
14718 => conv_std_logic_vector(28, 8),
14719 => conv_std_logic_vector(28, 8),
14720 => conv_std_logic_vector(28, 8),
14721 => conv_std_logic_vector(28, 8),
14722 => conv_std_logic_vector(28, 8),
14723 => conv_std_logic_vector(29, 8),
14724 => conv_std_logic_vector(29, 8),
14725 => conv_std_logic_vector(29, 8),
14726 => conv_std_logic_vector(29, 8),
14727 => conv_std_logic_vector(30, 8),
14728 => conv_std_logic_vector(30, 8),
14729 => conv_std_logic_vector(30, 8),
14730 => conv_std_logic_vector(30, 8),
14731 => conv_std_logic_vector(30, 8),
14732 => conv_std_logic_vector(31, 8),
14733 => conv_std_logic_vector(31, 8),
14734 => conv_std_logic_vector(31, 8),
14735 => conv_std_logic_vector(31, 8),
14736 => conv_std_logic_vector(32, 8),
14737 => conv_std_logic_vector(32, 8),
14738 => conv_std_logic_vector(32, 8),
14739 => conv_std_logic_vector(32, 8),
14740 => conv_std_logic_vector(32, 8),
14741 => conv_std_logic_vector(33, 8),
14742 => conv_std_logic_vector(33, 8),
14743 => conv_std_logic_vector(33, 8),
14744 => conv_std_logic_vector(33, 8),
14745 => conv_std_logic_vector(34, 8),
14746 => conv_std_logic_vector(34, 8),
14747 => conv_std_logic_vector(34, 8),
14748 => conv_std_logic_vector(34, 8),
14749 => conv_std_logic_vector(34, 8),
14750 => conv_std_logic_vector(35, 8),
14751 => conv_std_logic_vector(35, 8),
14752 => conv_std_logic_vector(35, 8),
14753 => conv_std_logic_vector(35, 8),
14754 => conv_std_logic_vector(36, 8),
14755 => conv_std_logic_vector(36, 8),
14756 => conv_std_logic_vector(36, 8),
14757 => conv_std_logic_vector(36, 8),
14758 => conv_std_logic_vector(36, 8),
14759 => conv_std_logic_vector(37, 8),
14760 => conv_std_logic_vector(37, 8),
14761 => conv_std_logic_vector(37, 8),
14762 => conv_std_logic_vector(37, 8),
14763 => conv_std_logic_vector(38, 8),
14764 => conv_std_logic_vector(38, 8),
14765 => conv_std_logic_vector(38, 8),
14766 => conv_std_logic_vector(38, 8),
14767 => conv_std_logic_vector(38, 8),
14768 => conv_std_logic_vector(39, 8),
14769 => conv_std_logic_vector(39, 8),
14770 => conv_std_logic_vector(39, 8),
14771 => conv_std_logic_vector(39, 8),
14772 => conv_std_logic_vector(40, 8),
14773 => conv_std_logic_vector(40, 8),
14774 => conv_std_logic_vector(40, 8),
14775 => conv_std_logic_vector(40, 8),
14776 => conv_std_logic_vector(40, 8),
14777 => conv_std_logic_vector(41, 8),
14778 => conv_std_logic_vector(41, 8),
14779 => conv_std_logic_vector(41, 8),
14780 => conv_std_logic_vector(41, 8),
14781 => conv_std_logic_vector(42, 8),
14782 => conv_std_logic_vector(42, 8),
14783 => conv_std_logic_vector(42, 8),
14784 => conv_std_logic_vector(42, 8),
14785 => conv_std_logic_vector(42, 8),
14786 => conv_std_logic_vector(43, 8),
14787 => conv_std_logic_vector(43, 8),
14788 => conv_std_logic_vector(43, 8),
14789 => conv_std_logic_vector(43, 8),
14790 => conv_std_logic_vector(44, 8),
14791 => conv_std_logic_vector(44, 8),
14792 => conv_std_logic_vector(44, 8),
14793 => conv_std_logic_vector(44, 8),
14794 => conv_std_logic_vector(44, 8),
14795 => conv_std_logic_vector(45, 8),
14796 => conv_std_logic_vector(45, 8),
14797 => conv_std_logic_vector(45, 8),
14798 => conv_std_logic_vector(45, 8),
14799 => conv_std_logic_vector(46, 8),
14800 => conv_std_logic_vector(46, 8),
14801 => conv_std_logic_vector(46, 8),
14802 => conv_std_logic_vector(46, 8),
14803 => conv_std_logic_vector(46, 8),
14804 => conv_std_logic_vector(47, 8),
14805 => conv_std_logic_vector(47, 8),
14806 => conv_std_logic_vector(47, 8),
14807 => conv_std_logic_vector(47, 8),
14808 => conv_std_logic_vector(48, 8),
14809 => conv_std_logic_vector(48, 8),
14810 => conv_std_logic_vector(48, 8),
14811 => conv_std_logic_vector(48, 8),
14812 => conv_std_logic_vector(48, 8),
14813 => conv_std_logic_vector(49, 8),
14814 => conv_std_logic_vector(49, 8),
14815 => conv_std_logic_vector(49, 8),
14816 => conv_std_logic_vector(49, 8),
14817 => conv_std_logic_vector(50, 8),
14818 => conv_std_logic_vector(50, 8),
14819 => conv_std_logic_vector(50, 8),
14820 => conv_std_logic_vector(50, 8),
14821 => conv_std_logic_vector(50, 8),
14822 => conv_std_logic_vector(51, 8),
14823 => conv_std_logic_vector(51, 8),
14824 => conv_std_logic_vector(51, 8),
14825 => conv_std_logic_vector(51, 8),
14826 => conv_std_logic_vector(52, 8),
14827 => conv_std_logic_vector(52, 8),
14828 => conv_std_logic_vector(52, 8),
14829 => conv_std_logic_vector(52, 8),
14830 => conv_std_logic_vector(52, 8),
14831 => conv_std_logic_vector(53, 8),
14832 => conv_std_logic_vector(53, 8),
14833 => conv_std_logic_vector(53, 8),
14834 => conv_std_logic_vector(53, 8),
14835 => conv_std_logic_vector(54, 8),
14836 => conv_std_logic_vector(54, 8),
14837 => conv_std_logic_vector(54, 8),
14838 => conv_std_logic_vector(54, 8),
14839 => conv_std_logic_vector(54, 8),
14840 => conv_std_logic_vector(55, 8),
14841 => conv_std_logic_vector(55, 8),
14842 => conv_std_logic_vector(55, 8),
14843 => conv_std_logic_vector(55, 8),
14844 => conv_std_logic_vector(56, 8),
14845 => conv_std_logic_vector(56, 8),
14846 => conv_std_logic_vector(56, 8),
14847 => conv_std_logic_vector(56, 8),
14848 => conv_std_logic_vector(0, 8),
14849 => conv_std_logic_vector(0, 8),
14850 => conv_std_logic_vector(0, 8),
14851 => conv_std_logic_vector(0, 8),
14852 => conv_std_logic_vector(0, 8),
14853 => conv_std_logic_vector(1, 8),
14854 => conv_std_logic_vector(1, 8),
14855 => conv_std_logic_vector(1, 8),
14856 => conv_std_logic_vector(1, 8),
14857 => conv_std_logic_vector(2, 8),
14858 => conv_std_logic_vector(2, 8),
14859 => conv_std_logic_vector(2, 8),
14860 => conv_std_logic_vector(2, 8),
14861 => conv_std_logic_vector(2, 8),
14862 => conv_std_logic_vector(3, 8),
14863 => conv_std_logic_vector(3, 8),
14864 => conv_std_logic_vector(3, 8),
14865 => conv_std_logic_vector(3, 8),
14866 => conv_std_logic_vector(4, 8),
14867 => conv_std_logic_vector(4, 8),
14868 => conv_std_logic_vector(4, 8),
14869 => conv_std_logic_vector(4, 8),
14870 => conv_std_logic_vector(4, 8),
14871 => conv_std_logic_vector(5, 8),
14872 => conv_std_logic_vector(5, 8),
14873 => conv_std_logic_vector(5, 8),
14874 => conv_std_logic_vector(5, 8),
14875 => conv_std_logic_vector(6, 8),
14876 => conv_std_logic_vector(6, 8),
14877 => conv_std_logic_vector(6, 8),
14878 => conv_std_logic_vector(6, 8),
14879 => conv_std_logic_vector(7, 8),
14880 => conv_std_logic_vector(7, 8),
14881 => conv_std_logic_vector(7, 8),
14882 => conv_std_logic_vector(7, 8),
14883 => conv_std_logic_vector(7, 8),
14884 => conv_std_logic_vector(8, 8),
14885 => conv_std_logic_vector(8, 8),
14886 => conv_std_logic_vector(8, 8),
14887 => conv_std_logic_vector(8, 8),
14888 => conv_std_logic_vector(9, 8),
14889 => conv_std_logic_vector(9, 8),
14890 => conv_std_logic_vector(9, 8),
14891 => conv_std_logic_vector(9, 8),
14892 => conv_std_logic_vector(9, 8),
14893 => conv_std_logic_vector(10, 8),
14894 => conv_std_logic_vector(10, 8),
14895 => conv_std_logic_vector(10, 8),
14896 => conv_std_logic_vector(10, 8),
14897 => conv_std_logic_vector(11, 8),
14898 => conv_std_logic_vector(11, 8),
14899 => conv_std_logic_vector(11, 8),
14900 => conv_std_logic_vector(11, 8),
14901 => conv_std_logic_vector(12, 8),
14902 => conv_std_logic_vector(12, 8),
14903 => conv_std_logic_vector(12, 8),
14904 => conv_std_logic_vector(12, 8),
14905 => conv_std_logic_vector(12, 8),
14906 => conv_std_logic_vector(13, 8),
14907 => conv_std_logic_vector(13, 8),
14908 => conv_std_logic_vector(13, 8),
14909 => conv_std_logic_vector(13, 8),
14910 => conv_std_logic_vector(14, 8),
14911 => conv_std_logic_vector(14, 8),
14912 => conv_std_logic_vector(14, 8),
14913 => conv_std_logic_vector(14, 8),
14914 => conv_std_logic_vector(14, 8),
14915 => conv_std_logic_vector(15, 8),
14916 => conv_std_logic_vector(15, 8),
14917 => conv_std_logic_vector(15, 8),
14918 => conv_std_logic_vector(15, 8),
14919 => conv_std_logic_vector(16, 8),
14920 => conv_std_logic_vector(16, 8),
14921 => conv_std_logic_vector(16, 8),
14922 => conv_std_logic_vector(16, 8),
14923 => conv_std_logic_vector(16, 8),
14924 => conv_std_logic_vector(17, 8),
14925 => conv_std_logic_vector(17, 8),
14926 => conv_std_logic_vector(17, 8),
14927 => conv_std_logic_vector(17, 8),
14928 => conv_std_logic_vector(18, 8),
14929 => conv_std_logic_vector(18, 8),
14930 => conv_std_logic_vector(18, 8),
14931 => conv_std_logic_vector(18, 8),
14932 => conv_std_logic_vector(19, 8),
14933 => conv_std_logic_vector(19, 8),
14934 => conv_std_logic_vector(19, 8),
14935 => conv_std_logic_vector(19, 8),
14936 => conv_std_logic_vector(19, 8),
14937 => conv_std_logic_vector(20, 8),
14938 => conv_std_logic_vector(20, 8),
14939 => conv_std_logic_vector(20, 8),
14940 => conv_std_logic_vector(20, 8),
14941 => conv_std_logic_vector(21, 8),
14942 => conv_std_logic_vector(21, 8),
14943 => conv_std_logic_vector(21, 8),
14944 => conv_std_logic_vector(21, 8),
14945 => conv_std_logic_vector(21, 8),
14946 => conv_std_logic_vector(22, 8),
14947 => conv_std_logic_vector(22, 8),
14948 => conv_std_logic_vector(22, 8),
14949 => conv_std_logic_vector(22, 8),
14950 => conv_std_logic_vector(23, 8),
14951 => conv_std_logic_vector(23, 8),
14952 => conv_std_logic_vector(23, 8),
14953 => conv_std_logic_vector(23, 8),
14954 => conv_std_logic_vector(24, 8),
14955 => conv_std_logic_vector(24, 8),
14956 => conv_std_logic_vector(24, 8),
14957 => conv_std_logic_vector(24, 8),
14958 => conv_std_logic_vector(24, 8),
14959 => conv_std_logic_vector(25, 8),
14960 => conv_std_logic_vector(25, 8),
14961 => conv_std_logic_vector(25, 8),
14962 => conv_std_logic_vector(25, 8),
14963 => conv_std_logic_vector(26, 8),
14964 => conv_std_logic_vector(26, 8),
14965 => conv_std_logic_vector(26, 8),
14966 => conv_std_logic_vector(26, 8),
14967 => conv_std_logic_vector(26, 8),
14968 => conv_std_logic_vector(27, 8),
14969 => conv_std_logic_vector(27, 8),
14970 => conv_std_logic_vector(27, 8),
14971 => conv_std_logic_vector(27, 8),
14972 => conv_std_logic_vector(28, 8),
14973 => conv_std_logic_vector(28, 8),
14974 => conv_std_logic_vector(28, 8),
14975 => conv_std_logic_vector(28, 8),
14976 => conv_std_logic_vector(29, 8),
14977 => conv_std_logic_vector(29, 8),
14978 => conv_std_logic_vector(29, 8),
14979 => conv_std_logic_vector(29, 8),
14980 => conv_std_logic_vector(29, 8),
14981 => conv_std_logic_vector(30, 8),
14982 => conv_std_logic_vector(30, 8),
14983 => conv_std_logic_vector(30, 8),
14984 => conv_std_logic_vector(30, 8),
14985 => conv_std_logic_vector(31, 8),
14986 => conv_std_logic_vector(31, 8),
14987 => conv_std_logic_vector(31, 8),
14988 => conv_std_logic_vector(31, 8),
14989 => conv_std_logic_vector(31, 8),
14990 => conv_std_logic_vector(32, 8),
14991 => conv_std_logic_vector(32, 8),
14992 => conv_std_logic_vector(32, 8),
14993 => conv_std_logic_vector(32, 8),
14994 => conv_std_logic_vector(33, 8),
14995 => conv_std_logic_vector(33, 8),
14996 => conv_std_logic_vector(33, 8),
14997 => conv_std_logic_vector(33, 8),
14998 => conv_std_logic_vector(33, 8),
14999 => conv_std_logic_vector(34, 8),
15000 => conv_std_logic_vector(34, 8),
15001 => conv_std_logic_vector(34, 8),
15002 => conv_std_logic_vector(34, 8),
15003 => conv_std_logic_vector(35, 8),
15004 => conv_std_logic_vector(35, 8),
15005 => conv_std_logic_vector(35, 8),
15006 => conv_std_logic_vector(35, 8),
15007 => conv_std_logic_vector(36, 8),
15008 => conv_std_logic_vector(36, 8),
15009 => conv_std_logic_vector(36, 8),
15010 => conv_std_logic_vector(36, 8),
15011 => conv_std_logic_vector(36, 8),
15012 => conv_std_logic_vector(37, 8),
15013 => conv_std_logic_vector(37, 8),
15014 => conv_std_logic_vector(37, 8),
15015 => conv_std_logic_vector(37, 8),
15016 => conv_std_logic_vector(38, 8),
15017 => conv_std_logic_vector(38, 8),
15018 => conv_std_logic_vector(38, 8),
15019 => conv_std_logic_vector(38, 8),
15020 => conv_std_logic_vector(38, 8),
15021 => conv_std_logic_vector(39, 8),
15022 => conv_std_logic_vector(39, 8),
15023 => conv_std_logic_vector(39, 8),
15024 => conv_std_logic_vector(39, 8),
15025 => conv_std_logic_vector(40, 8),
15026 => conv_std_logic_vector(40, 8),
15027 => conv_std_logic_vector(40, 8),
15028 => conv_std_logic_vector(40, 8),
15029 => conv_std_logic_vector(41, 8),
15030 => conv_std_logic_vector(41, 8),
15031 => conv_std_logic_vector(41, 8),
15032 => conv_std_logic_vector(41, 8),
15033 => conv_std_logic_vector(41, 8),
15034 => conv_std_logic_vector(42, 8),
15035 => conv_std_logic_vector(42, 8),
15036 => conv_std_logic_vector(42, 8),
15037 => conv_std_logic_vector(42, 8),
15038 => conv_std_logic_vector(43, 8),
15039 => conv_std_logic_vector(43, 8),
15040 => conv_std_logic_vector(43, 8),
15041 => conv_std_logic_vector(43, 8),
15042 => conv_std_logic_vector(43, 8),
15043 => conv_std_logic_vector(44, 8),
15044 => conv_std_logic_vector(44, 8),
15045 => conv_std_logic_vector(44, 8),
15046 => conv_std_logic_vector(44, 8),
15047 => conv_std_logic_vector(45, 8),
15048 => conv_std_logic_vector(45, 8),
15049 => conv_std_logic_vector(45, 8),
15050 => conv_std_logic_vector(45, 8),
15051 => conv_std_logic_vector(45, 8),
15052 => conv_std_logic_vector(46, 8),
15053 => conv_std_logic_vector(46, 8),
15054 => conv_std_logic_vector(46, 8),
15055 => conv_std_logic_vector(46, 8),
15056 => conv_std_logic_vector(47, 8),
15057 => conv_std_logic_vector(47, 8),
15058 => conv_std_logic_vector(47, 8),
15059 => conv_std_logic_vector(47, 8),
15060 => conv_std_logic_vector(48, 8),
15061 => conv_std_logic_vector(48, 8),
15062 => conv_std_logic_vector(48, 8),
15063 => conv_std_logic_vector(48, 8),
15064 => conv_std_logic_vector(48, 8),
15065 => conv_std_logic_vector(49, 8),
15066 => conv_std_logic_vector(49, 8),
15067 => conv_std_logic_vector(49, 8),
15068 => conv_std_logic_vector(49, 8),
15069 => conv_std_logic_vector(50, 8),
15070 => conv_std_logic_vector(50, 8),
15071 => conv_std_logic_vector(50, 8),
15072 => conv_std_logic_vector(50, 8),
15073 => conv_std_logic_vector(50, 8),
15074 => conv_std_logic_vector(51, 8),
15075 => conv_std_logic_vector(51, 8),
15076 => conv_std_logic_vector(51, 8),
15077 => conv_std_logic_vector(51, 8),
15078 => conv_std_logic_vector(52, 8),
15079 => conv_std_logic_vector(52, 8),
15080 => conv_std_logic_vector(52, 8),
15081 => conv_std_logic_vector(52, 8),
15082 => conv_std_logic_vector(53, 8),
15083 => conv_std_logic_vector(53, 8),
15084 => conv_std_logic_vector(53, 8),
15085 => conv_std_logic_vector(53, 8),
15086 => conv_std_logic_vector(53, 8),
15087 => conv_std_logic_vector(54, 8),
15088 => conv_std_logic_vector(54, 8),
15089 => conv_std_logic_vector(54, 8),
15090 => conv_std_logic_vector(54, 8),
15091 => conv_std_logic_vector(55, 8),
15092 => conv_std_logic_vector(55, 8),
15093 => conv_std_logic_vector(55, 8),
15094 => conv_std_logic_vector(55, 8),
15095 => conv_std_logic_vector(55, 8),
15096 => conv_std_logic_vector(56, 8),
15097 => conv_std_logic_vector(56, 8),
15098 => conv_std_logic_vector(56, 8),
15099 => conv_std_logic_vector(56, 8),
15100 => conv_std_logic_vector(57, 8),
15101 => conv_std_logic_vector(57, 8),
15102 => conv_std_logic_vector(57, 8),
15103 => conv_std_logic_vector(57, 8),
15104 => conv_std_logic_vector(0, 8),
15105 => conv_std_logic_vector(0, 8),
15106 => conv_std_logic_vector(0, 8),
15107 => conv_std_logic_vector(0, 8),
15108 => conv_std_logic_vector(0, 8),
15109 => conv_std_logic_vector(1, 8),
15110 => conv_std_logic_vector(1, 8),
15111 => conv_std_logic_vector(1, 8),
15112 => conv_std_logic_vector(1, 8),
15113 => conv_std_logic_vector(2, 8),
15114 => conv_std_logic_vector(2, 8),
15115 => conv_std_logic_vector(2, 8),
15116 => conv_std_logic_vector(2, 8),
15117 => conv_std_logic_vector(2, 8),
15118 => conv_std_logic_vector(3, 8),
15119 => conv_std_logic_vector(3, 8),
15120 => conv_std_logic_vector(3, 8),
15121 => conv_std_logic_vector(3, 8),
15122 => conv_std_logic_vector(4, 8),
15123 => conv_std_logic_vector(4, 8),
15124 => conv_std_logic_vector(4, 8),
15125 => conv_std_logic_vector(4, 8),
15126 => conv_std_logic_vector(5, 8),
15127 => conv_std_logic_vector(5, 8),
15128 => conv_std_logic_vector(5, 8),
15129 => conv_std_logic_vector(5, 8),
15130 => conv_std_logic_vector(5, 8),
15131 => conv_std_logic_vector(6, 8),
15132 => conv_std_logic_vector(6, 8),
15133 => conv_std_logic_vector(6, 8),
15134 => conv_std_logic_vector(6, 8),
15135 => conv_std_logic_vector(7, 8),
15136 => conv_std_logic_vector(7, 8),
15137 => conv_std_logic_vector(7, 8),
15138 => conv_std_logic_vector(7, 8),
15139 => conv_std_logic_vector(8, 8),
15140 => conv_std_logic_vector(8, 8),
15141 => conv_std_logic_vector(8, 8),
15142 => conv_std_logic_vector(8, 8),
15143 => conv_std_logic_vector(8, 8),
15144 => conv_std_logic_vector(9, 8),
15145 => conv_std_logic_vector(9, 8),
15146 => conv_std_logic_vector(9, 8),
15147 => conv_std_logic_vector(9, 8),
15148 => conv_std_logic_vector(10, 8),
15149 => conv_std_logic_vector(10, 8),
15150 => conv_std_logic_vector(10, 8),
15151 => conv_std_logic_vector(10, 8),
15152 => conv_std_logic_vector(11, 8),
15153 => conv_std_logic_vector(11, 8),
15154 => conv_std_logic_vector(11, 8),
15155 => conv_std_logic_vector(11, 8),
15156 => conv_std_logic_vector(11, 8),
15157 => conv_std_logic_vector(12, 8),
15158 => conv_std_logic_vector(12, 8),
15159 => conv_std_logic_vector(12, 8),
15160 => conv_std_logic_vector(12, 8),
15161 => conv_std_logic_vector(13, 8),
15162 => conv_std_logic_vector(13, 8),
15163 => conv_std_logic_vector(13, 8),
15164 => conv_std_logic_vector(13, 8),
15165 => conv_std_logic_vector(14, 8),
15166 => conv_std_logic_vector(14, 8),
15167 => conv_std_logic_vector(14, 8),
15168 => conv_std_logic_vector(14, 8),
15169 => conv_std_logic_vector(14, 8),
15170 => conv_std_logic_vector(15, 8),
15171 => conv_std_logic_vector(15, 8),
15172 => conv_std_logic_vector(15, 8),
15173 => conv_std_logic_vector(15, 8),
15174 => conv_std_logic_vector(16, 8),
15175 => conv_std_logic_vector(16, 8),
15176 => conv_std_logic_vector(16, 8),
15177 => conv_std_logic_vector(16, 8),
15178 => conv_std_logic_vector(17, 8),
15179 => conv_std_logic_vector(17, 8),
15180 => conv_std_logic_vector(17, 8),
15181 => conv_std_logic_vector(17, 8),
15182 => conv_std_logic_vector(17, 8),
15183 => conv_std_logic_vector(18, 8),
15184 => conv_std_logic_vector(18, 8),
15185 => conv_std_logic_vector(18, 8),
15186 => conv_std_logic_vector(18, 8),
15187 => conv_std_logic_vector(19, 8),
15188 => conv_std_logic_vector(19, 8),
15189 => conv_std_logic_vector(19, 8),
15190 => conv_std_logic_vector(19, 8),
15191 => conv_std_logic_vector(20, 8),
15192 => conv_std_logic_vector(20, 8),
15193 => conv_std_logic_vector(20, 8),
15194 => conv_std_logic_vector(20, 8),
15195 => conv_std_logic_vector(20, 8),
15196 => conv_std_logic_vector(21, 8),
15197 => conv_std_logic_vector(21, 8),
15198 => conv_std_logic_vector(21, 8),
15199 => conv_std_logic_vector(21, 8),
15200 => conv_std_logic_vector(22, 8),
15201 => conv_std_logic_vector(22, 8),
15202 => conv_std_logic_vector(22, 8),
15203 => conv_std_logic_vector(22, 8),
15204 => conv_std_logic_vector(23, 8),
15205 => conv_std_logic_vector(23, 8),
15206 => conv_std_logic_vector(23, 8),
15207 => conv_std_logic_vector(23, 8),
15208 => conv_std_logic_vector(23, 8),
15209 => conv_std_logic_vector(24, 8),
15210 => conv_std_logic_vector(24, 8),
15211 => conv_std_logic_vector(24, 8),
15212 => conv_std_logic_vector(24, 8),
15213 => conv_std_logic_vector(25, 8),
15214 => conv_std_logic_vector(25, 8),
15215 => conv_std_logic_vector(25, 8),
15216 => conv_std_logic_vector(25, 8),
15217 => conv_std_logic_vector(26, 8),
15218 => conv_std_logic_vector(26, 8),
15219 => conv_std_logic_vector(26, 8),
15220 => conv_std_logic_vector(26, 8),
15221 => conv_std_logic_vector(26, 8),
15222 => conv_std_logic_vector(27, 8),
15223 => conv_std_logic_vector(27, 8),
15224 => conv_std_logic_vector(27, 8),
15225 => conv_std_logic_vector(27, 8),
15226 => conv_std_logic_vector(28, 8),
15227 => conv_std_logic_vector(28, 8),
15228 => conv_std_logic_vector(28, 8),
15229 => conv_std_logic_vector(28, 8),
15230 => conv_std_logic_vector(29, 8),
15231 => conv_std_logic_vector(29, 8),
15232 => conv_std_logic_vector(29, 8),
15233 => conv_std_logic_vector(29, 8),
15234 => conv_std_logic_vector(29, 8),
15235 => conv_std_logic_vector(30, 8),
15236 => conv_std_logic_vector(30, 8),
15237 => conv_std_logic_vector(30, 8),
15238 => conv_std_logic_vector(30, 8),
15239 => conv_std_logic_vector(31, 8),
15240 => conv_std_logic_vector(31, 8),
15241 => conv_std_logic_vector(31, 8),
15242 => conv_std_logic_vector(31, 8),
15243 => conv_std_logic_vector(32, 8),
15244 => conv_std_logic_vector(32, 8),
15245 => conv_std_logic_vector(32, 8),
15246 => conv_std_logic_vector(32, 8),
15247 => conv_std_logic_vector(32, 8),
15248 => conv_std_logic_vector(33, 8),
15249 => conv_std_logic_vector(33, 8),
15250 => conv_std_logic_vector(33, 8),
15251 => conv_std_logic_vector(33, 8),
15252 => conv_std_logic_vector(34, 8),
15253 => conv_std_logic_vector(34, 8),
15254 => conv_std_logic_vector(34, 8),
15255 => conv_std_logic_vector(34, 8),
15256 => conv_std_logic_vector(35, 8),
15257 => conv_std_logic_vector(35, 8),
15258 => conv_std_logic_vector(35, 8),
15259 => conv_std_logic_vector(35, 8),
15260 => conv_std_logic_vector(35, 8),
15261 => conv_std_logic_vector(36, 8),
15262 => conv_std_logic_vector(36, 8),
15263 => conv_std_logic_vector(36, 8),
15264 => conv_std_logic_vector(36, 8),
15265 => conv_std_logic_vector(37, 8),
15266 => conv_std_logic_vector(37, 8),
15267 => conv_std_logic_vector(37, 8),
15268 => conv_std_logic_vector(37, 8),
15269 => conv_std_logic_vector(38, 8),
15270 => conv_std_logic_vector(38, 8),
15271 => conv_std_logic_vector(38, 8),
15272 => conv_std_logic_vector(38, 8),
15273 => conv_std_logic_vector(38, 8),
15274 => conv_std_logic_vector(39, 8),
15275 => conv_std_logic_vector(39, 8),
15276 => conv_std_logic_vector(39, 8),
15277 => conv_std_logic_vector(39, 8),
15278 => conv_std_logic_vector(40, 8),
15279 => conv_std_logic_vector(40, 8),
15280 => conv_std_logic_vector(40, 8),
15281 => conv_std_logic_vector(40, 8),
15282 => conv_std_logic_vector(41, 8),
15283 => conv_std_logic_vector(41, 8),
15284 => conv_std_logic_vector(41, 8),
15285 => conv_std_logic_vector(41, 8),
15286 => conv_std_logic_vector(41, 8),
15287 => conv_std_logic_vector(42, 8),
15288 => conv_std_logic_vector(42, 8),
15289 => conv_std_logic_vector(42, 8),
15290 => conv_std_logic_vector(42, 8),
15291 => conv_std_logic_vector(43, 8),
15292 => conv_std_logic_vector(43, 8),
15293 => conv_std_logic_vector(43, 8),
15294 => conv_std_logic_vector(43, 8),
15295 => conv_std_logic_vector(44, 8),
15296 => conv_std_logic_vector(44, 8),
15297 => conv_std_logic_vector(44, 8),
15298 => conv_std_logic_vector(44, 8),
15299 => conv_std_logic_vector(44, 8),
15300 => conv_std_logic_vector(45, 8),
15301 => conv_std_logic_vector(45, 8),
15302 => conv_std_logic_vector(45, 8),
15303 => conv_std_logic_vector(45, 8),
15304 => conv_std_logic_vector(46, 8),
15305 => conv_std_logic_vector(46, 8),
15306 => conv_std_logic_vector(46, 8),
15307 => conv_std_logic_vector(46, 8),
15308 => conv_std_logic_vector(47, 8),
15309 => conv_std_logic_vector(47, 8),
15310 => conv_std_logic_vector(47, 8),
15311 => conv_std_logic_vector(47, 8),
15312 => conv_std_logic_vector(47, 8),
15313 => conv_std_logic_vector(48, 8),
15314 => conv_std_logic_vector(48, 8),
15315 => conv_std_logic_vector(48, 8),
15316 => conv_std_logic_vector(48, 8),
15317 => conv_std_logic_vector(49, 8),
15318 => conv_std_logic_vector(49, 8),
15319 => conv_std_logic_vector(49, 8),
15320 => conv_std_logic_vector(49, 8),
15321 => conv_std_logic_vector(50, 8),
15322 => conv_std_logic_vector(50, 8),
15323 => conv_std_logic_vector(50, 8),
15324 => conv_std_logic_vector(50, 8),
15325 => conv_std_logic_vector(50, 8),
15326 => conv_std_logic_vector(51, 8),
15327 => conv_std_logic_vector(51, 8),
15328 => conv_std_logic_vector(51, 8),
15329 => conv_std_logic_vector(51, 8),
15330 => conv_std_logic_vector(52, 8),
15331 => conv_std_logic_vector(52, 8),
15332 => conv_std_logic_vector(52, 8),
15333 => conv_std_logic_vector(52, 8),
15334 => conv_std_logic_vector(53, 8),
15335 => conv_std_logic_vector(53, 8),
15336 => conv_std_logic_vector(53, 8),
15337 => conv_std_logic_vector(53, 8),
15338 => conv_std_logic_vector(53, 8),
15339 => conv_std_logic_vector(54, 8),
15340 => conv_std_logic_vector(54, 8),
15341 => conv_std_logic_vector(54, 8),
15342 => conv_std_logic_vector(54, 8),
15343 => conv_std_logic_vector(55, 8),
15344 => conv_std_logic_vector(55, 8),
15345 => conv_std_logic_vector(55, 8),
15346 => conv_std_logic_vector(55, 8),
15347 => conv_std_logic_vector(56, 8),
15348 => conv_std_logic_vector(56, 8),
15349 => conv_std_logic_vector(56, 8),
15350 => conv_std_logic_vector(56, 8),
15351 => conv_std_logic_vector(56, 8),
15352 => conv_std_logic_vector(57, 8),
15353 => conv_std_logic_vector(57, 8),
15354 => conv_std_logic_vector(57, 8),
15355 => conv_std_logic_vector(57, 8),
15356 => conv_std_logic_vector(58, 8),
15357 => conv_std_logic_vector(58, 8),
15358 => conv_std_logic_vector(58, 8),
15359 => conv_std_logic_vector(58, 8),
15360 => conv_std_logic_vector(0, 8),
15361 => conv_std_logic_vector(0, 8),
15362 => conv_std_logic_vector(0, 8),
15363 => conv_std_logic_vector(0, 8),
15364 => conv_std_logic_vector(0, 8),
15365 => conv_std_logic_vector(1, 8),
15366 => conv_std_logic_vector(1, 8),
15367 => conv_std_logic_vector(1, 8),
15368 => conv_std_logic_vector(1, 8),
15369 => conv_std_logic_vector(2, 8),
15370 => conv_std_logic_vector(2, 8),
15371 => conv_std_logic_vector(2, 8),
15372 => conv_std_logic_vector(2, 8),
15373 => conv_std_logic_vector(3, 8),
15374 => conv_std_logic_vector(3, 8),
15375 => conv_std_logic_vector(3, 8),
15376 => conv_std_logic_vector(3, 8),
15377 => conv_std_logic_vector(3, 8),
15378 => conv_std_logic_vector(4, 8),
15379 => conv_std_logic_vector(4, 8),
15380 => conv_std_logic_vector(4, 8),
15381 => conv_std_logic_vector(4, 8),
15382 => conv_std_logic_vector(5, 8),
15383 => conv_std_logic_vector(5, 8),
15384 => conv_std_logic_vector(5, 8),
15385 => conv_std_logic_vector(5, 8),
15386 => conv_std_logic_vector(6, 8),
15387 => conv_std_logic_vector(6, 8),
15388 => conv_std_logic_vector(6, 8),
15389 => conv_std_logic_vector(6, 8),
15390 => conv_std_logic_vector(7, 8),
15391 => conv_std_logic_vector(7, 8),
15392 => conv_std_logic_vector(7, 8),
15393 => conv_std_logic_vector(7, 8),
15394 => conv_std_logic_vector(7, 8),
15395 => conv_std_logic_vector(8, 8),
15396 => conv_std_logic_vector(8, 8),
15397 => conv_std_logic_vector(8, 8),
15398 => conv_std_logic_vector(8, 8),
15399 => conv_std_logic_vector(9, 8),
15400 => conv_std_logic_vector(9, 8),
15401 => conv_std_logic_vector(9, 8),
15402 => conv_std_logic_vector(9, 8),
15403 => conv_std_logic_vector(10, 8),
15404 => conv_std_logic_vector(10, 8),
15405 => conv_std_logic_vector(10, 8),
15406 => conv_std_logic_vector(10, 8),
15407 => conv_std_logic_vector(11, 8),
15408 => conv_std_logic_vector(11, 8),
15409 => conv_std_logic_vector(11, 8),
15410 => conv_std_logic_vector(11, 8),
15411 => conv_std_logic_vector(11, 8),
15412 => conv_std_logic_vector(12, 8),
15413 => conv_std_logic_vector(12, 8),
15414 => conv_std_logic_vector(12, 8),
15415 => conv_std_logic_vector(12, 8),
15416 => conv_std_logic_vector(13, 8),
15417 => conv_std_logic_vector(13, 8),
15418 => conv_std_logic_vector(13, 8),
15419 => conv_std_logic_vector(13, 8),
15420 => conv_std_logic_vector(14, 8),
15421 => conv_std_logic_vector(14, 8),
15422 => conv_std_logic_vector(14, 8),
15423 => conv_std_logic_vector(14, 8),
15424 => conv_std_logic_vector(15, 8),
15425 => conv_std_logic_vector(15, 8),
15426 => conv_std_logic_vector(15, 8),
15427 => conv_std_logic_vector(15, 8),
15428 => conv_std_logic_vector(15, 8),
15429 => conv_std_logic_vector(16, 8),
15430 => conv_std_logic_vector(16, 8),
15431 => conv_std_logic_vector(16, 8),
15432 => conv_std_logic_vector(16, 8),
15433 => conv_std_logic_vector(17, 8),
15434 => conv_std_logic_vector(17, 8),
15435 => conv_std_logic_vector(17, 8),
15436 => conv_std_logic_vector(17, 8),
15437 => conv_std_logic_vector(18, 8),
15438 => conv_std_logic_vector(18, 8),
15439 => conv_std_logic_vector(18, 8),
15440 => conv_std_logic_vector(18, 8),
15441 => conv_std_logic_vector(18, 8),
15442 => conv_std_logic_vector(19, 8),
15443 => conv_std_logic_vector(19, 8),
15444 => conv_std_logic_vector(19, 8),
15445 => conv_std_logic_vector(19, 8),
15446 => conv_std_logic_vector(20, 8),
15447 => conv_std_logic_vector(20, 8),
15448 => conv_std_logic_vector(20, 8),
15449 => conv_std_logic_vector(20, 8),
15450 => conv_std_logic_vector(21, 8),
15451 => conv_std_logic_vector(21, 8),
15452 => conv_std_logic_vector(21, 8),
15453 => conv_std_logic_vector(21, 8),
15454 => conv_std_logic_vector(22, 8),
15455 => conv_std_logic_vector(22, 8),
15456 => conv_std_logic_vector(22, 8),
15457 => conv_std_logic_vector(22, 8),
15458 => conv_std_logic_vector(22, 8),
15459 => conv_std_logic_vector(23, 8),
15460 => conv_std_logic_vector(23, 8),
15461 => conv_std_logic_vector(23, 8),
15462 => conv_std_logic_vector(23, 8),
15463 => conv_std_logic_vector(24, 8),
15464 => conv_std_logic_vector(24, 8),
15465 => conv_std_logic_vector(24, 8),
15466 => conv_std_logic_vector(24, 8),
15467 => conv_std_logic_vector(25, 8),
15468 => conv_std_logic_vector(25, 8),
15469 => conv_std_logic_vector(25, 8),
15470 => conv_std_logic_vector(25, 8),
15471 => conv_std_logic_vector(26, 8),
15472 => conv_std_logic_vector(26, 8),
15473 => conv_std_logic_vector(26, 8),
15474 => conv_std_logic_vector(26, 8),
15475 => conv_std_logic_vector(26, 8),
15476 => conv_std_logic_vector(27, 8),
15477 => conv_std_logic_vector(27, 8),
15478 => conv_std_logic_vector(27, 8),
15479 => conv_std_logic_vector(27, 8),
15480 => conv_std_logic_vector(28, 8),
15481 => conv_std_logic_vector(28, 8),
15482 => conv_std_logic_vector(28, 8),
15483 => conv_std_logic_vector(28, 8),
15484 => conv_std_logic_vector(29, 8),
15485 => conv_std_logic_vector(29, 8),
15486 => conv_std_logic_vector(29, 8),
15487 => conv_std_logic_vector(29, 8),
15488 => conv_std_logic_vector(30, 8),
15489 => conv_std_logic_vector(30, 8),
15490 => conv_std_logic_vector(30, 8),
15491 => conv_std_logic_vector(30, 8),
15492 => conv_std_logic_vector(30, 8),
15493 => conv_std_logic_vector(31, 8),
15494 => conv_std_logic_vector(31, 8),
15495 => conv_std_logic_vector(31, 8),
15496 => conv_std_logic_vector(31, 8),
15497 => conv_std_logic_vector(32, 8),
15498 => conv_std_logic_vector(32, 8),
15499 => conv_std_logic_vector(32, 8),
15500 => conv_std_logic_vector(32, 8),
15501 => conv_std_logic_vector(33, 8),
15502 => conv_std_logic_vector(33, 8),
15503 => conv_std_logic_vector(33, 8),
15504 => conv_std_logic_vector(33, 8),
15505 => conv_std_logic_vector(33, 8),
15506 => conv_std_logic_vector(34, 8),
15507 => conv_std_logic_vector(34, 8),
15508 => conv_std_logic_vector(34, 8),
15509 => conv_std_logic_vector(34, 8),
15510 => conv_std_logic_vector(35, 8),
15511 => conv_std_logic_vector(35, 8),
15512 => conv_std_logic_vector(35, 8),
15513 => conv_std_logic_vector(35, 8),
15514 => conv_std_logic_vector(36, 8),
15515 => conv_std_logic_vector(36, 8),
15516 => conv_std_logic_vector(36, 8),
15517 => conv_std_logic_vector(36, 8),
15518 => conv_std_logic_vector(37, 8),
15519 => conv_std_logic_vector(37, 8),
15520 => conv_std_logic_vector(37, 8),
15521 => conv_std_logic_vector(37, 8),
15522 => conv_std_logic_vector(37, 8),
15523 => conv_std_logic_vector(38, 8),
15524 => conv_std_logic_vector(38, 8),
15525 => conv_std_logic_vector(38, 8),
15526 => conv_std_logic_vector(38, 8),
15527 => conv_std_logic_vector(39, 8),
15528 => conv_std_logic_vector(39, 8),
15529 => conv_std_logic_vector(39, 8),
15530 => conv_std_logic_vector(39, 8),
15531 => conv_std_logic_vector(40, 8),
15532 => conv_std_logic_vector(40, 8),
15533 => conv_std_logic_vector(40, 8),
15534 => conv_std_logic_vector(40, 8),
15535 => conv_std_logic_vector(41, 8),
15536 => conv_std_logic_vector(41, 8),
15537 => conv_std_logic_vector(41, 8),
15538 => conv_std_logic_vector(41, 8),
15539 => conv_std_logic_vector(41, 8),
15540 => conv_std_logic_vector(42, 8),
15541 => conv_std_logic_vector(42, 8),
15542 => conv_std_logic_vector(42, 8),
15543 => conv_std_logic_vector(42, 8),
15544 => conv_std_logic_vector(43, 8),
15545 => conv_std_logic_vector(43, 8),
15546 => conv_std_logic_vector(43, 8),
15547 => conv_std_logic_vector(43, 8),
15548 => conv_std_logic_vector(44, 8),
15549 => conv_std_logic_vector(44, 8),
15550 => conv_std_logic_vector(44, 8),
15551 => conv_std_logic_vector(44, 8),
15552 => conv_std_logic_vector(45, 8),
15553 => conv_std_logic_vector(45, 8),
15554 => conv_std_logic_vector(45, 8),
15555 => conv_std_logic_vector(45, 8),
15556 => conv_std_logic_vector(45, 8),
15557 => conv_std_logic_vector(46, 8),
15558 => conv_std_logic_vector(46, 8),
15559 => conv_std_logic_vector(46, 8),
15560 => conv_std_logic_vector(46, 8),
15561 => conv_std_logic_vector(47, 8),
15562 => conv_std_logic_vector(47, 8),
15563 => conv_std_logic_vector(47, 8),
15564 => conv_std_logic_vector(47, 8),
15565 => conv_std_logic_vector(48, 8),
15566 => conv_std_logic_vector(48, 8),
15567 => conv_std_logic_vector(48, 8),
15568 => conv_std_logic_vector(48, 8),
15569 => conv_std_logic_vector(48, 8),
15570 => conv_std_logic_vector(49, 8),
15571 => conv_std_logic_vector(49, 8),
15572 => conv_std_logic_vector(49, 8),
15573 => conv_std_logic_vector(49, 8),
15574 => conv_std_logic_vector(50, 8),
15575 => conv_std_logic_vector(50, 8),
15576 => conv_std_logic_vector(50, 8),
15577 => conv_std_logic_vector(50, 8),
15578 => conv_std_logic_vector(51, 8),
15579 => conv_std_logic_vector(51, 8),
15580 => conv_std_logic_vector(51, 8),
15581 => conv_std_logic_vector(51, 8),
15582 => conv_std_logic_vector(52, 8),
15583 => conv_std_logic_vector(52, 8),
15584 => conv_std_logic_vector(52, 8),
15585 => conv_std_logic_vector(52, 8),
15586 => conv_std_logic_vector(52, 8),
15587 => conv_std_logic_vector(53, 8),
15588 => conv_std_logic_vector(53, 8),
15589 => conv_std_logic_vector(53, 8),
15590 => conv_std_logic_vector(53, 8),
15591 => conv_std_logic_vector(54, 8),
15592 => conv_std_logic_vector(54, 8),
15593 => conv_std_logic_vector(54, 8),
15594 => conv_std_logic_vector(54, 8),
15595 => conv_std_logic_vector(55, 8),
15596 => conv_std_logic_vector(55, 8),
15597 => conv_std_logic_vector(55, 8),
15598 => conv_std_logic_vector(55, 8),
15599 => conv_std_logic_vector(56, 8),
15600 => conv_std_logic_vector(56, 8),
15601 => conv_std_logic_vector(56, 8),
15602 => conv_std_logic_vector(56, 8),
15603 => conv_std_logic_vector(56, 8),
15604 => conv_std_logic_vector(57, 8),
15605 => conv_std_logic_vector(57, 8),
15606 => conv_std_logic_vector(57, 8),
15607 => conv_std_logic_vector(57, 8),
15608 => conv_std_logic_vector(58, 8),
15609 => conv_std_logic_vector(58, 8),
15610 => conv_std_logic_vector(58, 8),
15611 => conv_std_logic_vector(58, 8),
15612 => conv_std_logic_vector(59, 8),
15613 => conv_std_logic_vector(59, 8),
15614 => conv_std_logic_vector(59, 8),
15615 => conv_std_logic_vector(59, 8),
15616 => conv_std_logic_vector(0, 8),
15617 => conv_std_logic_vector(0, 8),
15618 => conv_std_logic_vector(0, 8),
15619 => conv_std_logic_vector(0, 8),
15620 => conv_std_logic_vector(0, 8),
15621 => conv_std_logic_vector(1, 8),
15622 => conv_std_logic_vector(1, 8),
15623 => conv_std_logic_vector(1, 8),
15624 => conv_std_logic_vector(1, 8),
15625 => conv_std_logic_vector(2, 8),
15626 => conv_std_logic_vector(2, 8),
15627 => conv_std_logic_vector(2, 8),
15628 => conv_std_logic_vector(2, 8),
15629 => conv_std_logic_vector(3, 8),
15630 => conv_std_logic_vector(3, 8),
15631 => conv_std_logic_vector(3, 8),
15632 => conv_std_logic_vector(3, 8),
15633 => conv_std_logic_vector(4, 8),
15634 => conv_std_logic_vector(4, 8),
15635 => conv_std_logic_vector(4, 8),
15636 => conv_std_logic_vector(4, 8),
15637 => conv_std_logic_vector(5, 8),
15638 => conv_std_logic_vector(5, 8),
15639 => conv_std_logic_vector(5, 8),
15640 => conv_std_logic_vector(5, 8),
15641 => conv_std_logic_vector(5, 8),
15642 => conv_std_logic_vector(6, 8),
15643 => conv_std_logic_vector(6, 8),
15644 => conv_std_logic_vector(6, 8),
15645 => conv_std_logic_vector(6, 8),
15646 => conv_std_logic_vector(7, 8),
15647 => conv_std_logic_vector(7, 8),
15648 => conv_std_logic_vector(7, 8),
15649 => conv_std_logic_vector(7, 8),
15650 => conv_std_logic_vector(8, 8),
15651 => conv_std_logic_vector(8, 8),
15652 => conv_std_logic_vector(8, 8),
15653 => conv_std_logic_vector(8, 8),
15654 => conv_std_logic_vector(9, 8),
15655 => conv_std_logic_vector(9, 8),
15656 => conv_std_logic_vector(9, 8),
15657 => conv_std_logic_vector(9, 8),
15658 => conv_std_logic_vector(10, 8),
15659 => conv_std_logic_vector(10, 8),
15660 => conv_std_logic_vector(10, 8),
15661 => conv_std_logic_vector(10, 8),
15662 => conv_std_logic_vector(10, 8),
15663 => conv_std_logic_vector(11, 8),
15664 => conv_std_logic_vector(11, 8),
15665 => conv_std_logic_vector(11, 8),
15666 => conv_std_logic_vector(11, 8),
15667 => conv_std_logic_vector(12, 8),
15668 => conv_std_logic_vector(12, 8),
15669 => conv_std_logic_vector(12, 8),
15670 => conv_std_logic_vector(12, 8),
15671 => conv_std_logic_vector(13, 8),
15672 => conv_std_logic_vector(13, 8),
15673 => conv_std_logic_vector(13, 8),
15674 => conv_std_logic_vector(13, 8),
15675 => conv_std_logic_vector(14, 8),
15676 => conv_std_logic_vector(14, 8),
15677 => conv_std_logic_vector(14, 8),
15678 => conv_std_logic_vector(14, 8),
15679 => conv_std_logic_vector(15, 8),
15680 => conv_std_logic_vector(15, 8),
15681 => conv_std_logic_vector(15, 8),
15682 => conv_std_logic_vector(15, 8),
15683 => conv_std_logic_vector(15, 8),
15684 => conv_std_logic_vector(16, 8),
15685 => conv_std_logic_vector(16, 8),
15686 => conv_std_logic_vector(16, 8),
15687 => conv_std_logic_vector(16, 8),
15688 => conv_std_logic_vector(17, 8),
15689 => conv_std_logic_vector(17, 8),
15690 => conv_std_logic_vector(17, 8),
15691 => conv_std_logic_vector(17, 8),
15692 => conv_std_logic_vector(18, 8),
15693 => conv_std_logic_vector(18, 8),
15694 => conv_std_logic_vector(18, 8),
15695 => conv_std_logic_vector(18, 8),
15696 => conv_std_logic_vector(19, 8),
15697 => conv_std_logic_vector(19, 8),
15698 => conv_std_logic_vector(19, 8),
15699 => conv_std_logic_vector(19, 8),
15700 => conv_std_logic_vector(20, 8),
15701 => conv_std_logic_vector(20, 8),
15702 => conv_std_logic_vector(20, 8),
15703 => conv_std_logic_vector(20, 8),
15704 => conv_std_logic_vector(20, 8),
15705 => conv_std_logic_vector(21, 8),
15706 => conv_std_logic_vector(21, 8),
15707 => conv_std_logic_vector(21, 8),
15708 => conv_std_logic_vector(21, 8),
15709 => conv_std_logic_vector(22, 8),
15710 => conv_std_logic_vector(22, 8),
15711 => conv_std_logic_vector(22, 8),
15712 => conv_std_logic_vector(22, 8),
15713 => conv_std_logic_vector(23, 8),
15714 => conv_std_logic_vector(23, 8),
15715 => conv_std_logic_vector(23, 8),
15716 => conv_std_logic_vector(23, 8),
15717 => conv_std_logic_vector(24, 8),
15718 => conv_std_logic_vector(24, 8),
15719 => conv_std_logic_vector(24, 8),
15720 => conv_std_logic_vector(24, 8),
15721 => conv_std_logic_vector(25, 8),
15722 => conv_std_logic_vector(25, 8),
15723 => conv_std_logic_vector(25, 8),
15724 => conv_std_logic_vector(25, 8),
15725 => conv_std_logic_vector(25, 8),
15726 => conv_std_logic_vector(26, 8),
15727 => conv_std_logic_vector(26, 8),
15728 => conv_std_logic_vector(26, 8),
15729 => conv_std_logic_vector(26, 8),
15730 => conv_std_logic_vector(27, 8),
15731 => conv_std_logic_vector(27, 8),
15732 => conv_std_logic_vector(27, 8),
15733 => conv_std_logic_vector(27, 8),
15734 => conv_std_logic_vector(28, 8),
15735 => conv_std_logic_vector(28, 8),
15736 => conv_std_logic_vector(28, 8),
15737 => conv_std_logic_vector(28, 8),
15738 => conv_std_logic_vector(29, 8),
15739 => conv_std_logic_vector(29, 8),
15740 => conv_std_logic_vector(29, 8),
15741 => conv_std_logic_vector(29, 8),
15742 => conv_std_logic_vector(30, 8),
15743 => conv_std_logic_vector(30, 8),
15744 => conv_std_logic_vector(30, 8),
15745 => conv_std_logic_vector(30, 8),
15746 => conv_std_logic_vector(30, 8),
15747 => conv_std_logic_vector(31, 8),
15748 => conv_std_logic_vector(31, 8),
15749 => conv_std_logic_vector(31, 8),
15750 => conv_std_logic_vector(31, 8),
15751 => conv_std_logic_vector(32, 8),
15752 => conv_std_logic_vector(32, 8),
15753 => conv_std_logic_vector(32, 8),
15754 => conv_std_logic_vector(32, 8),
15755 => conv_std_logic_vector(33, 8),
15756 => conv_std_logic_vector(33, 8),
15757 => conv_std_logic_vector(33, 8),
15758 => conv_std_logic_vector(33, 8),
15759 => conv_std_logic_vector(34, 8),
15760 => conv_std_logic_vector(34, 8),
15761 => conv_std_logic_vector(34, 8),
15762 => conv_std_logic_vector(34, 8),
15763 => conv_std_logic_vector(35, 8),
15764 => conv_std_logic_vector(35, 8),
15765 => conv_std_logic_vector(35, 8),
15766 => conv_std_logic_vector(35, 8),
15767 => conv_std_logic_vector(35, 8),
15768 => conv_std_logic_vector(36, 8),
15769 => conv_std_logic_vector(36, 8),
15770 => conv_std_logic_vector(36, 8),
15771 => conv_std_logic_vector(36, 8),
15772 => conv_std_logic_vector(37, 8),
15773 => conv_std_logic_vector(37, 8),
15774 => conv_std_logic_vector(37, 8),
15775 => conv_std_logic_vector(37, 8),
15776 => conv_std_logic_vector(38, 8),
15777 => conv_std_logic_vector(38, 8),
15778 => conv_std_logic_vector(38, 8),
15779 => conv_std_logic_vector(38, 8),
15780 => conv_std_logic_vector(39, 8),
15781 => conv_std_logic_vector(39, 8),
15782 => conv_std_logic_vector(39, 8),
15783 => conv_std_logic_vector(39, 8),
15784 => conv_std_logic_vector(40, 8),
15785 => conv_std_logic_vector(40, 8),
15786 => conv_std_logic_vector(40, 8),
15787 => conv_std_logic_vector(40, 8),
15788 => conv_std_logic_vector(40, 8),
15789 => conv_std_logic_vector(41, 8),
15790 => conv_std_logic_vector(41, 8),
15791 => conv_std_logic_vector(41, 8),
15792 => conv_std_logic_vector(41, 8),
15793 => conv_std_logic_vector(42, 8),
15794 => conv_std_logic_vector(42, 8),
15795 => conv_std_logic_vector(42, 8),
15796 => conv_std_logic_vector(42, 8),
15797 => conv_std_logic_vector(43, 8),
15798 => conv_std_logic_vector(43, 8),
15799 => conv_std_logic_vector(43, 8),
15800 => conv_std_logic_vector(43, 8),
15801 => conv_std_logic_vector(44, 8),
15802 => conv_std_logic_vector(44, 8),
15803 => conv_std_logic_vector(44, 8),
15804 => conv_std_logic_vector(44, 8),
15805 => conv_std_logic_vector(45, 8),
15806 => conv_std_logic_vector(45, 8),
15807 => conv_std_logic_vector(45, 8),
15808 => conv_std_logic_vector(45, 8),
15809 => conv_std_logic_vector(45, 8),
15810 => conv_std_logic_vector(46, 8),
15811 => conv_std_logic_vector(46, 8),
15812 => conv_std_logic_vector(46, 8),
15813 => conv_std_logic_vector(46, 8),
15814 => conv_std_logic_vector(47, 8),
15815 => conv_std_logic_vector(47, 8),
15816 => conv_std_logic_vector(47, 8),
15817 => conv_std_logic_vector(47, 8),
15818 => conv_std_logic_vector(48, 8),
15819 => conv_std_logic_vector(48, 8),
15820 => conv_std_logic_vector(48, 8),
15821 => conv_std_logic_vector(48, 8),
15822 => conv_std_logic_vector(49, 8),
15823 => conv_std_logic_vector(49, 8),
15824 => conv_std_logic_vector(49, 8),
15825 => conv_std_logic_vector(49, 8),
15826 => conv_std_logic_vector(50, 8),
15827 => conv_std_logic_vector(50, 8),
15828 => conv_std_logic_vector(50, 8),
15829 => conv_std_logic_vector(50, 8),
15830 => conv_std_logic_vector(50, 8),
15831 => conv_std_logic_vector(51, 8),
15832 => conv_std_logic_vector(51, 8),
15833 => conv_std_logic_vector(51, 8),
15834 => conv_std_logic_vector(51, 8),
15835 => conv_std_logic_vector(52, 8),
15836 => conv_std_logic_vector(52, 8),
15837 => conv_std_logic_vector(52, 8),
15838 => conv_std_logic_vector(52, 8),
15839 => conv_std_logic_vector(53, 8),
15840 => conv_std_logic_vector(53, 8),
15841 => conv_std_logic_vector(53, 8),
15842 => conv_std_logic_vector(53, 8),
15843 => conv_std_logic_vector(54, 8),
15844 => conv_std_logic_vector(54, 8),
15845 => conv_std_logic_vector(54, 8),
15846 => conv_std_logic_vector(54, 8),
15847 => conv_std_logic_vector(55, 8),
15848 => conv_std_logic_vector(55, 8),
15849 => conv_std_logic_vector(55, 8),
15850 => conv_std_logic_vector(55, 8),
15851 => conv_std_logic_vector(55, 8),
15852 => conv_std_logic_vector(56, 8),
15853 => conv_std_logic_vector(56, 8),
15854 => conv_std_logic_vector(56, 8),
15855 => conv_std_logic_vector(56, 8),
15856 => conv_std_logic_vector(57, 8),
15857 => conv_std_logic_vector(57, 8),
15858 => conv_std_logic_vector(57, 8),
15859 => conv_std_logic_vector(57, 8),
15860 => conv_std_logic_vector(58, 8),
15861 => conv_std_logic_vector(58, 8),
15862 => conv_std_logic_vector(58, 8),
15863 => conv_std_logic_vector(58, 8),
15864 => conv_std_logic_vector(59, 8),
15865 => conv_std_logic_vector(59, 8),
15866 => conv_std_logic_vector(59, 8),
15867 => conv_std_logic_vector(59, 8),
15868 => conv_std_logic_vector(60, 8),
15869 => conv_std_logic_vector(60, 8),
15870 => conv_std_logic_vector(60, 8),
15871 => conv_std_logic_vector(60, 8),
15872 => conv_std_logic_vector(0, 8),
15873 => conv_std_logic_vector(0, 8),
15874 => conv_std_logic_vector(0, 8),
15875 => conv_std_logic_vector(0, 8),
15876 => conv_std_logic_vector(0, 8),
15877 => conv_std_logic_vector(1, 8),
15878 => conv_std_logic_vector(1, 8),
15879 => conv_std_logic_vector(1, 8),
15880 => conv_std_logic_vector(1, 8),
15881 => conv_std_logic_vector(2, 8),
15882 => conv_std_logic_vector(2, 8),
15883 => conv_std_logic_vector(2, 8),
15884 => conv_std_logic_vector(2, 8),
15885 => conv_std_logic_vector(3, 8),
15886 => conv_std_logic_vector(3, 8),
15887 => conv_std_logic_vector(3, 8),
15888 => conv_std_logic_vector(3, 8),
15889 => conv_std_logic_vector(4, 8),
15890 => conv_std_logic_vector(4, 8),
15891 => conv_std_logic_vector(4, 8),
15892 => conv_std_logic_vector(4, 8),
15893 => conv_std_logic_vector(5, 8),
15894 => conv_std_logic_vector(5, 8),
15895 => conv_std_logic_vector(5, 8),
15896 => conv_std_logic_vector(5, 8),
15897 => conv_std_logic_vector(6, 8),
15898 => conv_std_logic_vector(6, 8),
15899 => conv_std_logic_vector(6, 8),
15900 => conv_std_logic_vector(6, 8),
15901 => conv_std_logic_vector(7, 8),
15902 => conv_std_logic_vector(7, 8),
15903 => conv_std_logic_vector(7, 8),
15904 => conv_std_logic_vector(7, 8),
15905 => conv_std_logic_vector(7, 8),
15906 => conv_std_logic_vector(8, 8),
15907 => conv_std_logic_vector(8, 8),
15908 => conv_std_logic_vector(8, 8),
15909 => conv_std_logic_vector(8, 8),
15910 => conv_std_logic_vector(9, 8),
15911 => conv_std_logic_vector(9, 8),
15912 => conv_std_logic_vector(9, 8),
15913 => conv_std_logic_vector(9, 8),
15914 => conv_std_logic_vector(10, 8),
15915 => conv_std_logic_vector(10, 8),
15916 => conv_std_logic_vector(10, 8),
15917 => conv_std_logic_vector(10, 8),
15918 => conv_std_logic_vector(11, 8),
15919 => conv_std_logic_vector(11, 8),
15920 => conv_std_logic_vector(11, 8),
15921 => conv_std_logic_vector(11, 8),
15922 => conv_std_logic_vector(12, 8),
15923 => conv_std_logic_vector(12, 8),
15924 => conv_std_logic_vector(12, 8),
15925 => conv_std_logic_vector(12, 8),
15926 => conv_std_logic_vector(13, 8),
15927 => conv_std_logic_vector(13, 8),
15928 => conv_std_logic_vector(13, 8),
15929 => conv_std_logic_vector(13, 8),
15930 => conv_std_logic_vector(14, 8),
15931 => conv_std_logic_vector(14, 8),
15932 => conv_std_logic_vector(14, 8),
15933 => conv_std_logic_vector(14, 8),
15934 => conv_std_logic_vector(15, 8),
15935 => conv_std_logic_vector(15, 8),
15936 => conv_std_logic_vector(15, 8),
15937 => conv_std_logic_vector(15, 8),
15938 => conv_std_logic_vector(15, 8),
15939 => conv_std_logic_vector(16, 8),
15940 => conv_std_logic_vector(16, 8),
15941 => conv_std_logic_vector(16, 8),
15942 => conv_std_logic_vector(16, 8),
15943 => conv_std_logic_vector(17, 8),
15944 => conv_std_logic_vector(17, 8),
15945 => conv_std_logic_vector(17, 8),
15946 => conv_std_logic_vector(17, 8),
15947 => conv_std_logic_vector(18, 8),
15948 => conv_std_logic_vector(18, 8),
15949 => conv_std_logic_vector(18, 8),
15950 => conv_std_logic_vector(18, 8),
15951 => conv_std_logic_vector(19, 8),
15952 => conv_std_logic_vector(19, 8),
15953 => conv_std_logic_vector(19, 8),
15954 => conv_std_logic_vector(19, 8),
15955 => conv_std_logic_vector(20, 8),
15956 => conv_std_logic_vector(20, 8),
15957 => conv_std_logic_vector(20, 8),
15958 => conv_std_logic_vector(20, 8),
15959 => conv_std_logic_vector(21, 8),
15960 => conv_std_logic_vector(21, 8),
15961 => conv_std_logic_vector(21, 8),
15962 => conv_std_logic_vector(21, 8),
15963 => conv_std_logic_vector(22, 8),
15964 => conv_std_logic_vector(22, 8),
15965 => conv_std_logic_vector(22, 8),
15966 => conv_std_logic_vector(22, 8),
15967 => conv_std_logic_vector(23, 8),
15968 => conv_std_logic_vector(23, 8),
15969 => conv_std_logic_vector(23, 8),
15970 => conv_std_logic_vector(23, 8),
15971 => conv_std_logic_vector(23, 8),
15972 => conv_std_logic_vector(24, 8),
15973 => conv_std_logic_vector(24, 8),
15974 => conv_std_logic_vector(24, 8),
15975 => conv_std_logic_vector(24, 8),
15976 => conv_std_logic_vector(25, 8),
15977 => conv_std_logic_vector(25, 8),
15978 => conv_std_logic_vector(25, 8),
15979 => conv_std_logic_vector(25, 8),
15980 => conv_std_logic_vector(26, 8),
15981 => conv_std_logic_vector(26, 8),
15982 => conv_std_logic_vector(26, 8),
15983 => conv_std_logic_vector(26, 8),
15984 => conv_std_logic_vector(27, 8),
15985 => conv_std_logic_vector(27, 8),
15986 => conv_std_logic_vector(27, 8),
15987 => conv_std_logic_vector(27, 8),
15988 => conv_std_logic_vector(28, 8),
15989 => conv_std_logic_vector(28, 8),
15990 => conv_std_logic_vector(28, 8),
15991 => conv_std_logic_vector(28, 8),
15992 => conv_std_logic_vector(29, 8),
15993 => conv_std_logic_vector(29, 8),
15994 => conv_std_logic_vector(29, 8),
15995 => conv_std_logic_vector(29, 8),
15996 => conv_std_logic_vector(30, 8),
15997 => conv_std_logic_vector(30, 8),
15998 => conv_std_logic_vector(30, 8),
15999 => conv_std_logic_vector(30, 8),
16000 => conv_std_logic_vector(31, 8),
16001 => conv_std_logic_vector(31, 8),
16002 => conv_std_logic_vector(31, 8),
16003 => conv_std_logic_vector(31, 8),
16004 => conv_std_logic_vector(31, 8),
16005 => conv_std_logic_vector(32, 8),
16006 => conv_std_logic_vector(32, 8),
16007 => conv_std_logic_vector(32, 8),
16008 => conv_std_logic_vector(32, 8),
16009 => conv_std_logic_vector(33, 8),
16010 => conv_std_logic_vector(33, 8),
16011 => conv_std_logic_vector(33, 8),
16012 => conv_std_logic_vector(33, 8),
16013 => conv_std_logic_vector(34, 8),
16014 => conv_std_logic_vector(34, 8),
16015 => conv_std_logic_vector(34, 8),
16016 => conv_std_logic_vector(34, 8),
16017 => conv_std_logic_vector(35, 8),
16018 => conv_std_logic_vector(35, 8),
16019 => conv_std_logic_vector(35, 8),
16020 => conv_std_logic_vector(35, 8),
16021 => conv_std_logic_vector(36, 8),
16022 => conv_std_logic_vector(36, 8),
16023 => conv_std_logic_vector(36, 8),
16024 => conv_std_logic_vector(36, 8),
16025 => conv_std_logic_vector(37, 8),
16026 => conv_std_logic_vector(37, 8),
16027 => conv_std_logic_vector(37, 8),
16028 => conv_std_logic_vector(37, 8),
16029 => conv_std_logic_vector(38, 8),
16030 => conv_std_logic_vector(38, 8),
16031 => conv_std_logic_vector(38, 8),
16032 => conv_std_logic_vector(38, 8),
16033 => conv_std_logic_vector(38, 8),
16034 => conv_std_logic_vector(39, 8),
16035 => conv_std_logic_vector(39, 8),
16036 => conv_std_logic_vector(39, 8),
16037 => conv_std_logic_vector(39, 8),
16038 => conv_std_logic_vector(40, 8),
16039 => conv_std_logic_vector(40, 8),
16040 => conv_std_logic_vector(40, 8),
16041 => conv_std_logic_vector(40, 8),
16042 => conv_std_logic_vector(41, 8),
16043 => conv_std_logic_vector(41, 8),
16044 => conv_std_logic_vector(41, 8),
16045 => conv_std_logic_vector(41, 8),
16046 => conv_std_logic_vector(42, 8),
16047 => conv_std_logic_vector(42, 8),
16048 => conv_std_logic_vector(42, 8),
16049 => conv_std_logic_vector(42, 8),
16050 => conv_std_logic_vector(43, 8),
16051 => conv_std_logic_vector(43, 8),
16052 => conv_std_logic_vector(43, 8),
16053 => conv_std_logic_vector(43, 8),
16054 => conv_std_logic_vector(44, 8),
16055 => conv_std_logic_vector(44, 8),
16056 => conv_std_logic_vector(44, 8),
16057 => conv_std_logic_vector(44, 8),
16058 => conv_std_logic_vector(45, 8),
16059 => conv_std_logic_vector(45, 8),
16060 => conv_std_logic_vector(45, 8),
16061 => conv_std_logic_vector(45, 8),
16062 => conv_std_logic_vector(46, 8),
16063 => conv_std_logic_vector(46, 8),
16064 => conv_std_logic_vector(46, 8),
16065 => conv_std_logic_vector(46, 8),
16066 => conv_std_logic_vector(46, 8),
16067 => conv_std_logic_vector(47, 8),
16068 => conv_std_logic_vector(47, 8),
16069 => conv_std_logic_vector(47, 8),
16070 => conv_std_logic_vector(47, 8),
16071 => conv_std_logic_vector(48, 8),
16072 => conv_std_logic_vector(48, 8),
16073 => conv_std_logic_vector(48, 8),
16074 => conv_std_logic_vector(48, 8),
16075 => conv_std_logic_vector(49, 8),
16076 => conv_std_logic_vector(49, 8),
16077 => conv_std_logic_vector(49, 8),
16078 => conv_std_logic_vector(49, 8),
16079 => conv_std_logic_vector(50, 8),
16080 => conv_std_logic_vector(50, 8),
16081 => conv_std_logic_vector(50, 8),
16082 => conv_std_logic_vector(50, 8),
16083 => conv_std_logic_vector(51, 8),
16084 => conv_std_logic_vector(51, 8),
16085 => conv_std_logic_vector(51, 8),
16086 => conv_std_logic_vector(51, 8),
16087 => conv_std_logic_vector(52, 8),
16088 => conv_std_logic_vector(52, 8),
16089 => conv_std_logic_vector(52, 8),
16090 => conv_std_logic_vector(52, 8),
16091 => conv_std_logic_vector(53, 8),
16092 => conv_std_logic_vector(53, 8),
16093 => conv_std_logic_vector(53, 8),
16094 => conv_std_logic_vector(53, 8),
16095 => conv_std_logic_vector(54, 8),
16096 => conv_std_logic_vector(54, 8),
16097 => conv_std_logic_vector(54, 8),
16098 => conv_std_logic_vector(54, 8),
16099 => conv_std_logic_vector(54, 8),
16100 => conv_std_logic_vector(55, 8),
16101 => conv_std_logic_vector(55, 8),
16102 => conv_std_logic_vector(55, 8),
16103 => conv_std_logic_vector(55, 8),
16104 => conv_std_logic_vector(56, 8),
16105 => conv_std_logic_vector(56, 8),
16106 => conv_std_logic_vector(56, 8),
16107 => conv_std_logic_vector(56, 8),
16108 => conv_std_logic_vector(57, 8),
16109 => conv_std_logic_vector(57, 8),
16110 => conv_std_logic_vector(57, 8),
16111 => conv_std_logic_vector(57, 8),
16112 => conv_std_logic_vector(58, 8),
16113 => conv_std_logic_vector(58, 8),
16114 => conv_std_logic_vector(58, 8),
16115 => conv_std_logic_vector(58, 8),
16116 => conv_std_logic_vector(59, 8),
16117 => conv_std_logic_vector(59, 8),
16118 => conv_std_logic_vector(59, 8),
16119 => conv_std_logic_vector(59, 8),
16120 => conv_std_logic_vector(60, 8),
16121 => conv_std_logic_vector(60, 8),
16122 => conv_std_logic_vector(60, 8),
16123 => conv_std_logic_vector(60, 8),
16124 => conv_std_logic_vector(61, 8),
16125 => conv_std_logic_vector(61, 8),
16126 => conv_std_logic_vector(61, 8),
16127 => conv_std_logic_vector(61, 8),
16128 => conv_std_logic_vector(0, 8),
16129 => conv_std_logic_vector(0, 8),
16130 => conv_std_logic_vector(0, 8),
16131 => conv_std_logic_vector(0, 8),
16132 => conv_std_logic_vector(0, 8),
16133 => conv_std_logic_vector(1, 8),
16134 => conv_std_logic_vector(1, 8),
16135 => conv_std_logic_vector(1, 8),
16136 => conv_std_logic_vector(1, 8),
16137 => conv_std_logic_vector(2, 8),
16138 => conv_std_logic_vector(2, 8),
16139 => conv_std_logic_vector(2, 8),
16140 => conv_std_logic_vector(2, 8),
16141 => conv_std_logic_vector(3, 8),
16142 => conv_std_logic_vector(3, 8),
16143 => conv_std_logic_vector(3, 8),
16144 => conv_std_logic_vector(3, 8),
16145 => conv_std_logic_vector(4, 8),
16146 => conv_std_logic_vector(4, 8),
16147 => conv_std_logic_vector(4, 8),
16148 => conv_std_logic_vector(4, 8),
16149 => conv_std_logic_vector(5, 8),
16150 => conv_std_logic_vector(5, 8),
16151 => conv_std_logic_vector(5, 8),
16152 => conv_std_logic_vector(5, 8),
16153 => conv_std_logic_vector(6, 8),
16154 => conv_std_logic_vector(6, 8),
16155 => conv_std_logic_vector(6, 8),
16156 => conv_std_logic_vector(6, 8),
16157 => conv_std_logic_vector(7, 8),
16158 => conv_std_logic_vector(7, 8),
16159 => conv_std_logic_vector(7, 8),
16160 => conv_std_logic_vector(7, 8),
16161 => conv_std_logic_vector(8, 8),
16162 => conv_std_logic_vector(8, 8),
16163 => conv_std_logic_vector(8, 8),
16164 => conv_std_logic_vector(8, 8),
16165 => conv_std_logic_vector(9, 8),
16166 => conv_std_logic_vector(9, 8),
16167 => conv_std_logic_vector(9, 8),
16168 => conv_std_logic_vector(9, 8),
16169 => conv_std_logic_vector(10, 8),
16170 => conv_std_logic_vector(10, 8),
16171 => conv_std_logic_vector(10, 8),
16172 => conv_std_logic_vector(10, 8),
16173 => conv_std_logic_vector(11, 8),
16174 => conv_std_logic_vector(11, 8),
16175 => conv_std_logic_vector(11, 8),
16176 => conv_std_logic_vector(11, 8),
16177 => conv_std_logic_vector(12, 8),
16178 => conv_std_logic_vector(12, 8),
16179 => conv_std_logic_vector(12, 8),
16180 => conv_std_logic_vector(12, 8),
16181 => conv_std_logic_vector(13, 8),
16182 => conv_std_logic_vector(13, 8),
16183 => conv_std_logic_vector(13, 8),
16184 => conv_std_logic_vector(13, 8),
16185 => conv_std_logic_vector(14, 8),
16186 => conv_std_logic_vector(14, 8),
16187 => conv_std_logic_vector(14, 8),
16188 => conv_std_logic_vector(14, 8),
16189 => conv_std_logic_vector(15, 8),
16190 => conv_std_logic_vector(15, 8),
16191 => conv_std_logic_vector(15, 8),
16192 => conv_std_logic_vector(15, 8),
16193 => conv_std_logic_vector(15, 8),
16194 => conv_std_logic_vector(16, 8),
16195 => conv_std_logic_vector(16, 8),
16196 => conv_std_logic_vector(16, 8),
16197 => conv_std_logic_vector(16, 8),
16198 => conv_std_logic_vector(17, 8),
16199 => conv_std_logic_vector(17, 8),
16200 => conv_std_logic_vector(17, 8),
16201 => conv_std_logic_vector(17, 8),
16202 => conv_std_logic_vector(18, 8),
16203 => conv_std_logic_vector(18, 8),
16204 => conv_std_logic_vector(18, 8),
16205 => conv_std_logic_vector(18, 8),
16206 => conv_std_logic_vector(19, 8),
16207 => conv_std_logic_vector(19, 8),
16208 => conv_std_logic_vector(19, 8),
16209 => conv_std_logic_vector(19, 8),
16210 => conv_std_logic_vector(20, 8),
16211 => conv_std_logic_vector(20, 8),
16212 => conv_std_logic_vector(20, 8),
16213 => conv_std_logic_vector(20, 8),
16214 => conv_std_logic_vector(21, 8),
16215 => conv_std_logic_vector(21, 8),
16216 => conv_std_logic_vector(21, 8),
16217 => conv_std_logic_vector(21, 8),
16218 => conv_std_logic_vector(22, 8),
16219 => conv_std_logic_vector(22, 8),
16220 => conv_std_logic_vector(22, 8),
16221 => conv_std_logic_vector(22, 8),
16222 => conv_std_logic_vector(23, 8),
16223 => conv_std_logic_vector(23, 8),
16224 => conv_std_logic_vector(23, 8),
16225 => conv_std_logic_vector(23, 8),
16226 => conv_std_logic_vector(24, 8),
16227 => conv_std_logic_vector(24, 8),
16228 => conv_std_logic_vector(24, 8),
16229 => conv_std_logic_vector(24, 8),
16230 => conv_std_logic_vector(25, 8),
16231 => conv_std_logic_vector(25, 8),
16232 => conv_std_logic_vector(25, 8),
16233 => conv_std_logic_vector(25, 8),
16234 => conv_std_logic_vector(26, 8),
16235 => conv_std_logic_vector(26, 8),
16236 => conv_std_logic_vector(26, 8),
16237 => conv_std_logic_vector(26, 8),
16238 => conv_std_logic_vector(27, 8),
16239 => conv_std_logic_vector(27, 8),
16240 => conv_std_logic_vector(27, 8),
16241 => conv_std_logic_vector(27, 8),
16242 => conv_std_logic_vector(28, 8),
16243 => conv_std_logic_vector(28, 8),
16244 => conv_std_logic_vector(28, 8),
16245 => conv_std_logic_vector(28, 8),
16246 => conv_std_logic_vector(29, 8),
16247 => conv_std_logic_vector(29, 8),
16248 => conv_std_logic_vector(29, 8),
16249 => conv_std_logic_vector(29, 8),
16250 => conv_std_logic_vector(30, 8),
16251 => conv_std_logic_vector(30, 8),
16252 => conv_std_logic_vector(30, 8),
16253 => conv_std_logic_vector(30, 8),
16254 => conv_std_logic_vector(31, 8),
16255 => conv_std_logic_vector(31, 8),
16256 => conv_std_logic_vector(31, 8),
16257 => conv_std_logic_vector(31, 8),
16258 => conv_std_logic_vector(31, 8),
16259 => conv_std_logic_vector(32, 8),
16260 => conv_std_logic_vector(32, 8),
16261 => conv_std_logic_vector(32, 8),
16262 => conv_std_logic_vector(32, 8),
16263 => conv_std_logic_vector(33, 8),
16264 => conv_std_logic_vector(33, 8),
16265 => conv_std_logic_vector(33, 8),
16266 => conv_std_logic_vector(33, 8),
16267 => conv_std_logic_vector(34, 8),
16268 => conv_std_logic_vector(34, 8),
16269 => conv_std_logic_vector(34, 8),
16270 => conv_std_logic_vector(34, 8),
16271 => conv_std_logic_vector(35, 8),
16272 => conv_std_logic_vector(35, 8),
16273 => conv_std_logic_vector(35, 8),
16274 => conv_std_logic_vector(35, 8),
16275 => conv_std_logic_vector(36, 8),
16276 => conv_std_logic_vector(36, 8),
16277 => conv_std_logic_vector(36, 8),
16278 => conv_std_logic_vector(36, 8),
16279 => conv_std_logic_vector(37, 8),
16280 => conv_std_logic_vector(37, 8),
16281 => conv_std_logic_vector(37, 8),
16282 => conv_std_logic_vector(37, 8),
16283 => conv_std_logic_vector(38, 8),
16284 => conv_std_logic_vector(38, 8),
16285 => conv_std_logic_vector(38, 8),
16286 => conv_std_logic_vector(38, 8),
16287 => conv_std_logic_vector(39, 8),
16288 => conv_std_logic_vector(39, 8),
16289 => conv_std_logic_vector(39, 8),
16290 => conv_std_logic_vector(39, 8),
16291 => conv_std_logic_vector(40, 8),
16292 => conv_std_logic_vector(40, 8),
16293 => conv_std_logic_vector(40, 8),
16294 => conv_std_logic_vector(40, 8),
16295 => conv_std_logic_vector(41, 8),
16296 => conv_std_logic_vector(41, 8),
16297 => conv_std_logic_vector(41, 8),
16298 => conv_std_logic_vector(41, 8),
16299 => conv_std_logic_vector(42, 8),
16300 => conv_std_logic_vector(42, 8),
16301 => conv_std_logic_vector(42, 8),
16302 => conv_std_logic_vector(42, 8),
16303 => conv_std_logic_vector(43, 8),
16304 => conv_std_logic_vector(43, 8),
16305 => conv_std_logic_vector(43, 8),
16306 => conv_std_logic_vector(43, 8),
16307 => conv_std_logic_vector(44, 8),
16308 => conv_std_logic_vector(44, 8),
16309 => conv_std_logic_vector(44, 8),
16310 => conv_std_logic_vector(44, 8),
16311 => conv_std_logic_vector(45, 8),
16312 => conv_std_logic_vector(45, 8),
16313 => conv_std_logic_vector(45, 8),
16314 => conv_std_logic_vector(45, 8),
16315 => conv_std_logic_vector(46, 8),
16316 => conv_std_logic_vector(46, 8),
16317 => conv_std_logic_vector(46, 8),
16318 => conv_std_logic_vector(46, 8),
16319 => conv_std_logic_vector(47, 8),
16320 => conv_std_logic_vector(47, 8),
16321 => conv_std_logic_vector(47, 8),
16322 => conv_std_logic_vector(47, 8),
16323 => conv_std_logic_vector(47, 8),
16324 => conv_std_logic_vector(48, 8),
16325 => conv_std_logic_vector(48, 8),
16326 => conv_std_logic_vector(48, 8),
16327 => conv_std_logic_vector(48, 8),
16328 => conv_std_logic_vector(49, 8),
16329 => conv_std_logic_vector(49, 8),
16330 => conv_std_logic_vector(49, 8),
16331 => conv_std_logic_vector(49, 8),
16332 => conv_std_logic_vector(50, 8),
16333 => conv_std_logic_vector(50, 8),
16334 => conv_std_logic_vector(50, 8),
16335 => conv_std_logic_vector(50, 8),
16336 => conv_std_logic_vector(51, 8),
16337 => conv_std_logic_vector(51, 8),
16338 => conv_std_logic_vector(51, 8),
16339 => conv_std_logic_vector(51, 8),
16340 => conv_std_logic_vector(52, 8),
16341 => conv_std_logic_vector(52, 8),
16342 => conv_std_logic_vector(52, 8),
16343 => conv_std_logic_vector(52, 8),
16344 => conv_std_logic_vector(53, 8),
16345 => conv_std_logic_vector(53, 8),
16346 => conv_std_logic_vector(53, 8),
16347 => conv_std_logic_vector(53, 8),
16348 => conv_std_logic_vector(54, 8),
16349 => conv_std_logic_vector(54, 8),
16350 => conv_std_logic_vector(54, 8),
16351 => conv_std_logic_vector(54, 8),
16352 => conv_std_logic_vector(55, 8),
16353 => conv_std_logic_vector(55, 8),
16354 => conv_std_logic_vector(55, 8),
16355 => conv_std_logic_vector(55, 8),
16356 => conv_std_logic_vector(56, 8),
16357 => conv_std_logic_vector(56, 8),
16358 => conv_std_logic_vector(56, 8),
16359 => conv_std_logic_vector(56, 8),
16360 => conv_std_logic_vector(57, 8),
16361 => conv_std_logic_vector(57, 8),
16362 => conv_std_logic_vector(57, 8),
16363 => conv_std_logic_vector(57, 8),
16364 => conv_std_logic_vector(58, 8),
16365 => conv_std_logic_vector(58, 8),
16366 => conv_std_logic_vector(58, 8),
16367 => conv_std_logic_vector(58, 8),
16368 => conv_std_logic_vector(59, 8),
16369 => conv_std_logic_vector(59, 8),
16370 => conv_std_logic_vector(59, 8),
16371 => conv_std_logic_vector(59, 8),
16372 => conv_std_logic_vector(60, 8),
16373 => conv_std_logic_vector(60, 8),
16374 => conv_std_logic_vector(60, 8),
16375 => conv_std_logic_vector(60, 8),
16376 => conv_std_logic_vector(61, 8),
16377 => conv_std_logic_vector(61, 8),
16378 => conv_std_logic_vector(61, 8),
16379 => conv_std_logic_vector(61, 8),
16380 => conv_std_logic_vector(62, 8),
16381 => conv_std_logic_vector(62, 8),
16382 => conv_std_logic_vector(62, 8),
16383 => conv_std_logic_vector(62, 8),
16384 => conv_std_logic_vector(0, 8),
16385 => conv_std_logic_vector(0, 8),
16386 => conv_std_logic_vector(0, 8),
16387 => conv_std_logic_vector(0, 8),
16388 => conv_std_logic_vector(1, 8),
16389 => conv_std_logic_vector(1, 8),
16390 => conv_std_logic_vector(1, 8),
16391 => conv_std_logic_vector(1, 8),
16392 => conv_std_logic_vector(2, 8),
16393 => conv_std_logic_vector(2, 8),
16394 => conv_std_logic_vector(2, 8),
16395 => conv_std_logic_vector(2, 8),
16396 => conv_std_logic_vector(3, 8),
16397 => conv_std_logic_vector(3, 8),
16398 => conv_std_logic_vector(3, 8),
16399 => conv_std_logic_vector(3, 8),
16400 => conv_std_logic_vector(4, 8),
16401 => conv_std_logic_vector(4, 8),
16402 => conv_std_logic_vector(4, 8),
16403 => conv_std_logic_vector(4, 8),
16404 => conv_std_logic_vector(5, 8),
16405 => conv_std_logic_vector(5, 8),
16406 => conv_std_logic_vector(5, 8),
16407 => conv_std_logic_vector(5, 8),
16408 => conv_std_logic_vector(6, 8),
16409 => conv_std_logic_vector(6, 8),
16410 => conv_std_logic_vector(6, 8),
16411 => conv_std_logic_vector(6, 8),
16412 => conv_std_logic_vector(7, 8),
16413 => conv_std_logic_vector(7, 8),
16414 => conv_std_logic_vector(7, 8),
16415 => conv_std_logic_vector(7, 8),
16416 => conv_std_logic_vector(8, 8),
16417 => conv_std_logic_vector(8, 8),
16418 => conv_std_logic_vector(8, 8),
16419 => conv_std_logic_vector(8, 8),
16420 => conv_std_logic_vector(9, 8),
16421 => conv_std_logic_vector(9, 8),
16422 => conv_std_logic_vector(9, 8),
16423 => conv_std_logic_vector(9, 8),
16424 => conv_std_logic_vector(10, 8),
16425 => conv_std_logic_vector(10, 8),
16426 => conv_std_logic_vector(10, 8),
16427 => conv_std_logic_vector(10, 8),
16428 => conv_std_logic_vector(11, 8),
16429 => conv_std_logic_vector(11, 8),
16430 => conv_std_logic_vector(11, 8),
16431 => conv_std_logic_vector(11, 8),
16432 => conv_std_logic_vector(12, 8),
16433 => conv_std_logic_vector(12, 8),
16434 => conv_std_logic_vector(12, 8),
16435 => conv_std_logic_vector(12, 8),
16436 => conv_std_logic_vector(13, 8),
16437 => conv_std_logic_vector(13, 8),
16438 => conv_std_logic_vector(13, 8),
16439 => conv_std_logic_vector(13, 8),
16440 => conv_std_logic_vector(14, 8),
16441 => conv_std_logic_vector(14, 8),
16442 => conv_std_logic_vector(14, 8),
16443 => conv_std_logic_vector(14, 8),
16444 => conv_std_logic_vector(15, 8),
16445 => conv_std_logic_vector(15, 8),
16446 => conv_std_logic_vector(15, 8),
16447 => conv_std_logic_vector(15, 8),
16448 => conv_std_logic_vector(16, 8),
16449 => conv_std_logic_vector(16, 8),
16450 => conv_std_logic_vector(16, 8),
16451 => conv_std_logic_vector(16, 8),
16452 => conv_std_logic_vector(17, 8),
16453 => conv_std_logic_vector(17, 8),
16454 => conv_std_logic_vector(17, 8),
16455 => conv_std_logic_vector(17, 8),
16456 => conv_std_logic_vector(18, 8),
16457 => conv_std_logic_vector(18, 8),
16458 => conv_std_logic_vector(18, 8),
16459 => conv_std_logic_vector(18, 8),
16460 => conv_std_logic_vector(19, 8),
16461 => conv_std_logic_vector(19, 8),
16462 => conv_std_logic_vector(19, 8),
16463 => conv_std_logic_vector(19, 8),
16464 => conv_std_logic_vector(20, 8),
16465 => conv_std_logic_vector(20, 8),
16466 => conv_std_logic_vector(20, 8),
16467 => conv_std_logic_vector(20, 8),
16468 => conv_std_logic_vector(21, 8),
16469 => conv_std_logic_vector(21, 8),
16470 => conv_std_logic_vector(21, 8),
16471 => conv_std_logic_vector(21, 8),
16472 => conv_std_logic_vector(22, 8),
16473 => conv_std_logic_vector(22, 8),
16474 => conv_std_logic_vector(22, 8),
16475 => conv_std_logic_vector(22, 8),
16476 => conv_std_logic_vector(23, 8),
16477 => conv_std_logic_vector(23, 8),
16478 => conv_std_logic_vector(23, 8),
16479 => conv_std_logic_vector(23, 8),
16480 => conv_std_logic_vector(24, 8),
16481 => conv_std_logic_vector(24, 8),
16482 => conv_std_logic_vector(24, 8),
16483 => conv_std_logic_vector(24, 8),
16484 => conv_std_logic_vector(25, 8),
16485 => conv_std_logic_vector(25, 8),
16486 => conv_std_logic_vector(25, 8),
16487 => conv_std_logic_vector(25, 8),
16488 => conv_std_logic_vector(26, 8),
16489 => conv_std_logic_vector(26, 8),
16490 => conv_std_logic_vector(26, 8),
16491 => conv_std_logic_vector(26, 8),
16492 => conv_std_logic_vector(27, 8),
16493 => conv_std_logic_vector(27, 8),
16494 => conv_std_logic_vector(27, 8),
16495 => conv_std_logic_vector(27, 8),
16496 => conv_std_logic_vector(28, 8),
16497 => conv_std_logic_vector(28, 8),
16498 => conv_std_logic_vector(28, 8),
16499 => conv_std_logic_vector(28, 8),
16500 => conv_std_logic_vector(29, 8),
16501 => conv_std_logic_vector(29, 8),
16502 => conv_std_logic_vector(29, 8),
16503 => conv_std_logic_vector(29, 8),
16504 => conv_std_logic_vector(30, 8),
16505 => conv_std_logic_vector(30, 8),
16506 => conv_std_logic_vector(30, 8),
16507 => conv_std_logic_vector(30, 8),
16508 => conv_std_logic_vector(31, 8),
16509 => conv_std_logic_vector(31, 8),
16510 => conv_std_logic_vector(31, 8),
16511 => conv_std_logic_vector(31, 8),
16512 => conv_std_logic_vector(32, 8),
16513 => conv_std_logic_vector(32, 8),
16514 => conv_std_logic_vector(32, 8),
16515 => conv_std_logic_vector(32, 8),
16516 => conv_std_logic_vector(33, 8),
16517 => conv_std_logic_vector(33, 8),
16518 => conv_std_logic_vector(33, 8),
16519 => conv_std_logic_vector(33, 8),
16520 => conv_std_logic_vector(34, 8),
16521 => conv_std_logic_vector(34, 8),
16522 => conv_std_logic_vector(34, 8),
16523 => conv_std_logic_vector(34, 8),
16524 => conv_std_logic_vector(35, 8),
16525 => conv_std_logic_vector(35, 8),
16526 => conv_std_logic_vector(35, 8),
16527 => conv_std_logic_vector(35, 8),
16528 => conv_std_logic_vector(36, 8),
16529 => conv_std_logic_vector(36, 8),
16530 => conv_std_logic_vector(36, 8),
16531 => conv_std_logic_vector(36, 8),
16532 => conv_std_logic_vector(37, 8),
16533 => conv_std_logic_vector(37, 8),
16534 => conv_std_logic_vector(37, 8),
16535 => conv_std_logic_vector(37, 8),
16536 => conv_std_logic_vector(38, 8),
16537 => conv_std_logic_vector(38, 8),
16538 => conv_std_logic_vector(38, 8),
16539 => conv_std_logic_vector(38, 8),
16540 => conv_std_logic_vector(39, 8),
16541 => conv_std_logic_vector(39, 8),
16542 => conv_std_logic_vector(39, 8),
16543 => conv_std_logic_vector(39, 8),
16544 => conv_std_logic_vector(40, 8),
16545 => conv_std_logic_vector(40, 8),
16546 => conv_std_logic_vector(40, 8),
16547 => conv_std_logic_vector(40, 8),
16548 => conv_std_logic_vector(41, 8),
16549 => conv_std_logic_vector(41, 8),
16550 => conv_std_logic_vector(41, 8),
16551 => conv_std_logic_vector(41, 8),
16552 => conv_std_logic_vector(42, 8),
16553 => conv_std_logic_vector(42, 8),
16554 => conv_std_logic_vector(42, 8),
16555 => conv_std_logic_vector(42, 8),
16556 => conv_std_logic_vector(43, 8),
16557 => conv_std_logic_vector(43, 8),
16558 => conv_std_logic_vector(43, 8),
16559 => conv_std_logic_vector(43, 8),
16560 => conv_std_logic_vector(44, 8),
16561 => conv_std_logic_vector(44, 8),
16562 => conv_std_logic_vector(44, 8),
16563 => conv_std_logic_vector(44, 8),
16564 => conv_std_logic_vector(45, 8),
16565 => conv_std_logic_vector(45, 8),
16566 => conv_std_logic_vector(45, 8),
16567 => conv_std_logic_vector(45, 8),
16568 => conv_std_logic_vector(46, 8),
16569 => conv_std_logic_vector(46, 8),
16570 => conv_std_logic_vector(46, 8),
16571 => conv_std_logic_vector(46, 8),
16572 => conv_std_logic_vector(47, 8),
16573 => conv_std_logic_vector(47, 8),
16574 => conv_std_logic_vector(47, 8),
16575 => conv_std_logic_vector(47, 8),
16576 => conv_std_logic_vector(48, 8),
16577 => conv_std_logic_vector(48, 8),
16578 => conv_std_logic_vector(48, 8),
16579 => conv_std_logic_vector(48, 8),
16580 => conv_std_logic_vector(49, 8),
16581 => conv_std_logic_vector(49, 8),
16582 => conv_std_logic_vector(49, 8),
16583 => conv_std_logic_vector(49, 8),
16584 => conv_std_logic_vector(50, 8),
16585 => conv_std_logic_vector(50, 8),
16586 => conv_std_logic_vector(50, 8),
16587 => conv_std_logic_vector(50, 8),
16588 => conv_std_logic_vector(51, 8),
16589 => conv_std_logic_vector(51, 8),
16590 => conv_std_logic_vector(51, 8),
16591 => conv_std_logic_vector(51, 8),
16592 => conv_std_logic_vector(52, 8),
16593 => conv_std_logic_vector(52, 8),
16594 => conv_std_logic_vector(52, 8),
16595 => conv_std_logic_vector(52, 8),
16596 => conv_std_logic_vector(53, 8),
16597 => conv_std_logic_vector(53, 8),
16598 => conv_std_logic_vector(53, 8),
16599 => conv_std_logic_vector(53, 8),
16600 => conv_std_logic_vector(54, 8),
16601 => conv_std_logic_vector(54, 8),
16602 => conv_std_logic_vector(54, 8),
16603 => conv_std_logic_vector(54, 8),
16604 => conv_std_logic_vector(55, 8),
16605 => conv_std_logic_vector(55, 8),
16606 => conv_std_logic_vector(55, 8),
16607 => conv_std_logic_vector(55, 8),
16608 => conv_std_logic_vector(56, 8),
16609 => conv_std_logic_vector(56, 8),
16610 => conv_std_logic_vector(56, 8),
16611 => conv_std_logic_vector(56, 8),
16612 => conv_std_logic_vector(57, 8),
16613 => conv_std_logic_vector(57, 8),
16614 => conv_std_logic_vector(57, 8),
16615 => conv_std_logic_vector(57, 8),
16616 => conv_std_logic_vector(58, 8),
16617 => conv_std_logic_vector(58, 8),
16618 => conv_std_logic_vector(58, 8),
16619 => conv_std_logic_vector(58, 8),
16620 => conv_std_logic_vector(59, 8),
16621 => conv_std_logic_vector(59, 8),
16622 => conv_std_logic_vector(59, 8),
16623 => conv_std_logic_vector(59, 8),
16624 => conv_std_logic_vector(60, 8),
16625 => conv_std_logic_vector(60, 8),
16626 => conv_std_logic_vector(60, 8),
16627 => conv_std_logic_vector(60, 8),
16628 => conv_std_logic_vector(61, 8),
16629 => conv_std_logic_vector(61, 8),
16630 => conv_std_logic_vector(61, 8),
16631 => conv_std_logic_vector(61, 8),
16632 => conv_std_logic_vector(62, 8),
16633 => conv_std_logic_vector(62, 8),
16634 => conv_std_logic_vector(62, 8),
16635 => conv_std_logic_vector(62, 8),
16636 => conv_std_logic_vector(63, 8),
16637 => conv_std_logic_vector(63, 8),
16638 => conv_std_logic_vector(63, 8),
16639 => conv_std_logic_vector(63, 8),
16640 => conv_std_logic_vector(0, 8),
16641 => conv_std_logic_vector(0, 8),
16642 => conv_std_logic_vector(0, 8),
16643 => conv_std_logic_vector(0, 8),
16644 => conv_std_logic_vector(1, 8),
16645 => conv_std_logic_vector(1, 8),
16646 => conv_std_logic_vector(1, 8),
16647 => conv_std_logic_vector(1, 8),
16648 => conv_std_logic_vector(2, 8),
16649 => conv_std_logic_vector(2, 8),
16650 => conv_std_logic_vector(2, 8),
16651 => conv_std_logic_vector(2, 8),
16652 => conv_std_logic_vector(3, 8),
16653 => conv_std_logic_vector(3, 8),
16654 => conv_std_logic_vector(3, 8),
16655 => conv_std_logic_vector(3, 8),
16656 => conv_std_logic_vector(4, 8),
16657 => conv_std_logic_vector(4, 8),
16658 => conv_std_logic_vector(4, 8),
16659 => conv_std_logic_vector(4, 8),
16660 => conv_std_logic_vector(5, 8),
16661 => conv_std_logic_vector(5, 8),
16662 => conv_std_logic_vector(5, 8),
16663 => conv_std_logic_vector(5, 8),
16664 => conv_std_logic_vector(6, 8),
16665 => conv_std_logic_vector(6, 8),
16666 => conv_std_logic_vector(6, 8),
16667 => conv_std_logic_vector(6, 8),
16668 => conv_std_logic_vector(7, 8),
16669 => conv_std_logic_vector(7, 8),
16670 => conv_std_logic_vector(7, 8),
16671 => conv_std_logic_vector(7, 8),
16672 => conv_std_logic_vector(8, 8),
16673 => conv_std_logic_vector(8, 8),
16674 => conv_std_logic_vector(8, 8),
16675 => conv_std_logic_vector(8, 8),
16676 => conv_std_logic_vector(9, 8),
16677 => conv_std_logic_vector(9, 8),
16678 => conv_std_logic_vector(9, 8),
16679 => conv_std_logic_vector(9, 8),
16680 => conv_std_logic_vector(10, 8),
16681 => conv_std_logic_vector(10, 8),
16682 => conv_std_logic_vector(10, 8),
16683 => conv_std_logic_vector(10, 8),
16684 => conv_std_logic_vector(11, 8),
16685 => conv_std_logic_vector(11, 8),
16686 => conv_std_logic_vector(11, 8),
16687 => conv_std_logic_vector(11, 8),
16688 => conv_std_logic_vector(12, 8),
16689 => conv_std_logic_vector(12, 8),
16690 => conv_std_logic_vector(12, 8),
16691 => conv_std_logic_vector(12, 8),
16692 => conv_std_logic_vector(13, 8),
16693 => conv_std_logic_vector(13, 8),
16694 => conv_std_logic_vector(13, 8),
16695 => conv_std_logic_vector(13, 8),
16696 => conv_std_logic_vector(14, 8),
16697 => conv_std_logic_vector(14, 8),
16698 => conv_std_logic_vector(14, 8),
16699 => conv_std_logic_vector(14, 8),
16700 => conv_std_logic_vector(15, 8),
16701 => conv_std_logic_vector(15, 8),
16702 => conv_std_logic_vector(15, 8),
16703 => conv_std_logic_vector(15, 8),
16704 => conv_std_logic_vector(16, 8),
16705 => conv_std_logic_vector(16, 8),
16706 => conv_std_logic_vector(16, 8),
16707 => conv_std_logic_vector(17, 8),
16708 => conv_std_logic_vector(17, 8),
16709 => conv_std_logic_vector(17, 8),
16710 => conv_std_logic_vector(17, 8),
16711 => conv_std_logic_vector(18, 8),
16712 => conv_std_logic_vector(18, 8),
16713 => conv_std_logic_vector(18, 8),
16714 => conv_std_logic_vector(18, 8),
16715 => conv_std_logic_vector(19, 8),
16716 => conv_std_logic_vector(19, 8),
16717 => conv_std_logic_vector(19, 8),
16718 => conv_std_logic_vector(19, 8),
16719 => conv_std_logic_vector(20, 8),
16720 => conv_std_logic_vector(20, 8),
16721 => conv_std_logic_vector(20, 8),
16722 => conv_std_logic_vector(20, 8),
16723 => conv_std_logic_vector(21, 8),
16724 => conv_std_logic_vector(21, 8),
16725 => conv_std_logic_vector(21, 8),
16726 => conv_std_logic_vector(21, 8),
16727 => conv_std_logic_vector(22, 8),
16728 => conv_std_logic_vector(22, 8),
16729 => conv_std_logic_vector(22, 8),
16730 => conv_std_logic_vector(22, 8),
16731 => conv_std_logic_vector(23, 8),
16732 => conv_std_logic_vector(23, 8),
16733 => conv_std_logic_vector(23, 8),
16734 => conv_std_logic_vector(23, 8),
16735 => conv_std_logic_vector(24, 8),
16736 => conv_std_logic_vector(24, 8),
16737 => conv_std_logic_vector(24, 8),
16738 => conv_std_logic_vector(24, 8),
16739 => conv_std_logic_vector(25, 8),
16740 => conv_std_logic_vector(25, 8),
16741 => conv_std_logic_vector(25, 8),
16742 => conv_std_logic_vector(25, 8),
16743 => conv_std_logic_vector(26, 8),
16744 => conv_std_logic_vector(26, 8),
16745 => conv_std_logic_vector(26, 8),
16746 => conv_std_logic_vector(26, 8),
16747 => conv_std_logic_vector(27, 8),
16748 => conv_std_logic_vector(27, 8),
16749 => conv_std_logic_vector(27, 8),
16750 => conv_std_logic_vector(27, 8),
16751 => conv_std_logic_vector(28, 8),
16752 => conv_std_logic_vector(28, 8),
16753 => conv_std_logic_vector(28, 8),
16754 => conv_std_logic_vector(28, 8),
16755 => conv_std_logic_vector(29, 8),
16756 => conv_std_logic_vector(29, 8),
16757 => conv_std_logic_vector(29, 8),
16758 => conv_std_logic_vector(29, 8),
16759 => conv_std_logic_vector(30, 8),
16760 => conv_std_logic_vector(30, 8),
16761 => conv_std_logic_vector(30, 8),
16762 => conv_std_logic_vector(30, 8),
16763 => conv_std_logic_vector(31, 8),
16764 => conv_std_logic_vector(31, 8),
16765 => conv_std_logic_vector(31, 8),
16766 => conv_std_logic_vector(31, 8),
16767 => conv_std_logic_vector(32, 8),
16768 => conv_std_logic_vector(32, 8),
16769 => conv_std_logic_vector(32, 8),
16770 => conv_std_logic_vector(33, 8),
16771 => conv_std_logic_vector(33, 8),
16772 => conv_std_logic_vector(33, 8),
16773 => conv_std_logic_vector(33, 8),
16774 => conv_std_logic_vector(34, 8),
16775 => conv_std_logic_vector(34, 8),
16776 => conv_std_logic_vector(34, 8),
16777 => conv_std_logic_vector(34, 8),
16778 => conv_std_logic_vector(35, 8),
16779 => conv_std_logic_vector(35, 8),
16780 => conv_std_logic_vector(35, 8),
16781 => conv_std_logic_vector(35, 8),
16782 => conv_std_logic_vector(36, 8),
16783 => conv_std_logic_vector(36, 8),
16784 => conv_std_logic_vector(36, 8),
16785 => conv_std_logic_vector(36, 8),
16786 => conv_std_logic_vector(37, 8),
16787 => conv_std_logic_vector(37, 8),
16788 => conv_std_logic_vector(37, 8),
16789 => conv_std_logic_vector(37, 8),
16790 => conv_std_logic_vector(38, 8),
16791 => conv_std_logic_vector(38, 8),
16792 => conv_std_logic_vector(38, 8),
16793 => conv_std_logic_vector(38, 8),
16794 => conv_std_logic_vector(39, 8),
16795 => conv_std_logic_vector(39, 8),
16796 => conv_std_logic_vector(39, 8),
16797 => conv_std_logic_vector(39, 8),
16798 => conv_std_logic_vector(40, 8),
16799 => conv_std_logic_vector(40, 8),
16800 => conv_std_logic_vector(40, 8),
16801 => conv_std_logic_vector(40, 8),
16802 => conv_std_logic_vector(41, 8),
16803 => conv_std_logic_vector(41, 8),
16804 => conv_std_logic_vector(41, 8),
16805 => conv_std_logic_vector(41, 8),
16806 => conv_std_logic_vector(42, 8),
16807 => conv_std_logic_vector(42, 8),
16808 => conv_std_logic_vector(42, 8),
16809 => conv_std_logic_vector(42, 8),
16810 => conv_std_logic_vector(43, 8),
16811 => conv_std_logic_vector(43, 8),
16812 => conv_std_logic_vector(43, 8),
16813 => conv_std_logic_vector(43, 8),
16814 => conv_std_logic_vector(44, 8),
16815 => conv_std_logic_vector(44, 8),
16816 => conv_std_logic_vector(44, 8),
16817 => conv_std_logic_vector(44, 8),
16818 => conv_std_logic_vector(45, 8),
16819 => conv_std_logic_vector(45, 8),
16820 => conv_std_logic_vector(45, 8),
16821 => conv_std_logic_vector(45, 8),
16822 => conv_std_logic_vector(46, 8),
16823 => conv_std_logic_vector(46, 8),
16824 => conv_std_logic_vector(46, 8),
16825 => conv_std_logic_vector(46, 8),
16826 => conv_std_logic_vector(47, 8),
16827 => conv_std_logic_vector(47, 8),
16828 => conv_std_logic_vector(47, 8),
16829 => conv_std_logic_vector(47, 8),
16830 => conv_std_logic_vector(48, 8),
16831 => conv_std_logic_vector(48, 8),
16832 => conv_std_logic_vector(48, 8),
16833 => conv_std_logic_vector(49, 8),
16834 => conv_std_logic_vector(49, 8),
16835 => conv_std_logic_vector(49, 8),
16836 => conv_std_logic_vector(49, 8),
16837 => conv_std_logic_vector(50, 8),
16838 => conv_std_logic_vector(50, 8),
16839 => conv_std_logic_vector(50, 8),
16840 => conv_std_logic_vector(50, 8),
16841 => conv_std_logic_vector(51, 8),
16842 => conv_std_logic_vector(51, 8),
16843 => conv_std_logic_vector(51, 8),
16844 => conv_std_logic_vector(51, 8),
16845 => conv_std_logic_vector(52, 8),
16846 => conv_std_logic_vector(52, 8),
16847 => conv_std_logic_vector(52, 8),
16848 => conv_std_logic_vector(52, 8),
16849 => conv_std_logic_vector(53, 8),
16850 => conv_std_logic_vector(53, 8),
16851 => conv_std_logic_vector(53, 8),
16852 => conv_std_logic_vector(53, 8),
16853 => conv_std_logic_vector(54, 8),
16854 => conv_std_logic_vector(54, 8),
16855 => conv_std_logic_vector(54, 8),
16856 => conv_std_logic_vector(54, 8),
16857 => conv_std_logic_vector(55, 8),
16858 => conv_std_logic_vector(55, 8),
16859 => conv_std_logic_vector(55, 8),
16860 => conv_std_logic_vector(55, 8),
16861 => conv_std_logic_vector(56, 8),
16862 => conv_std_logic_vector(56, 8),
16863 => conv_std_logic_vector(56, 8),
16864 => conv_std_logic_vector(56, 8),
16865 => conv_std_logic_vector(57, 8),
16866 => conv_std_logic_vector(57, 8),
16867 => conv_std_logic_vector(57, 8),
16868 => conv_std_logic_vector(57, 8),
16869 => conv_std_logic_vector(58, 8),
16870 => conv_std_logic_vector(58, 8),
16871 => conv_std_logic_vector(58, 8),
16872 => conv_std_logic_vector(58, 8),
16873 => conv_std_logic_vector(59, 8),
16874 => conv_std_logic_vector(59, 8),
16875 => conv_std_logic_vector(59, 8),
16876 => conv_std_logic_vector(59, 8),
16877 => conv_std_logic_vector(60, 8),
16878 => conv_std_logic_vector(60, 8),
16879 => conv_std_logic_vector(60, 8),
16880 => conv_std_logic_vector(60, 8),
16881 => conv_std_logic_vector(61, 8),
16882 => conv_std_logic_vector(61, 8),
16883 => conv_std_logic_vector(61, 8),
16884 => conv_std_logic_vector(61, 8),
16885 => conv_std_logic_vector(62, 8),
16886 => conv_std_logic_vector(62, 8),
16887 => conv_std_logic_vector(62, 8),
16888 => conv_std_logic_vector(62, 8),
16889 => conv_std_logic_vector(63, 8),
16890 => conv_std_logic_vector(63, 8),
16891 => conv_std_logic_vector(63, 8),
16892 => conv_std_logic_vector(63, 8),
16893 => conv_std_logic_vector(64, 8),
16894 => conv_std_logic_vector(64, 8),
16895 => conv_std_logic_vector(64, 8),
16896 => conv_std_logic_vector(0, 8),
16897 => conv_std_logic_vector(0, 8),
16898 => conv_std_logic_vector(0, 8),
16899 => conv_std_logic_vector(0, 8),
16900 => conv_std_logic_vector(1, 8),
16901 => conv_std_logic_vector(1, 8),
16902 => conv_std_logic_vector(1, 8),
16903 => conv_std_logic_vector(1, 8),
16904 => conv_std_logic_vector(2, 8),
16905 => conv_std_logic_vector(2, 8),
16906 => conv_std_logic_vector(2, 8),
16907 => conv_std_logic_vector(2, 8),
16908 => conv_std_logic_vector(3, 8),
16909 => conv_std_logic_vector(3, 8),
16910 => conv_std_logic_vector(3, 8),
16911 => conv_std_logic_vector(3, 8),
16912 => conv_std_logic_vector(4, 8),
16913 => conv_std_logic_vector(4, 8),
16914 => conv_std_logic_vector(4, 8),
16915 => conv_std_logic_vector(4, 8),
16916 => conv_std_logic_vector(5, 8),
16917 => conv_std_logic_vector(5, 8),
16918 => conv_std_logic_vector(5, 8),
16919 => conv_std_logic_vector(5, 8),
16920 => conv_std_logic_vector(6, 8),
16921 => conv_std_logic_vector(6, 8),
16922 => conv_std_logic_vector(6, 8),
16923 => conv_std_logic_vector(6, 8),
16924 => conv_std_logic_vector(7, 8),
16925 => conv_std_logic_vector(7, 8),
16926 => conv_std_logic_vector(7, 8),
16927 => conv_std_logic_vector(7, 8),
16928 => conv_std_logic_vector(8, 8),
16929 => conv_std_logic_vector(8, 8),
16930 => conv_std_logic_vector(8, 8),
16931 => conv_std_logic_vector(9, 8),
16932 => conv_std_logic_vector(9, 8),
16933 => conv_std_logic_vector(9, 8),
16934 => conv_std_logic_vector(9, 8),
16935 => conv_std_logic_vector(10, 8),
16936 => conv_std_logic_vector(10, 8),
16937 => conv_std_logic_vector(10, 8),
16938 => conv_std_logic_vector(10, 8),
16939 => conv_std_logic_vector(11, 8),
16940 => conv_std_logic_vector(11, 8),
16941 => conv_std_logic_vector(11, 8),
16942 => conv_std_logic_vector(11, 8),
16943 => conv_std_logic_vector(12, 8),
16944 => conv_std_logic_vector(12, 8),
16945 => conv_std_logic_vector(12, 8),
16946 => conv_std_logic_vector(12, 8),
16947 => conv_std_logic_vector(13, 8),
16948 => conv_std_logic_vector(13, 8),
16949 => conv_std_logic_vector(13, 8),
16950 => conv_std_logic_vector(13, 8),
16951 => conv_std_logic_vector(14, 8),
16952 => conv_std_logic_vector(14, 8),
16953 => conv_std_logic_vector(14, 8),
16954 => conv_std_logic_vector(14, 8),
16955 => conv_std_logic_vector(15, 8),
16956 => conv_std_logic_vector(15, 8),
16957 => conv_std_logic_vector(15, 8),
16958 => conv_std_logic_vector(15, 8),
16959 => conv_std_logic_vector(16, 8),
16960 => conv_std_logic_vector(16, 8),
16961 => conv_std_logic_vector(16, 8),
16962 => conv_std_logic_vector(17, 8),
16963 => conv_std_logic_vector(17, 8),
16964 => conv_std_logic_vector(17, 8),
16965 => conv_std_logic_vector(17, 8),
16966 => conv_std_logic_vector(18, 8),
16967 => conv_std_logic_vector(18, 8),
16968 => conv_std_logic_vector(18, 8),
16969 => conv_std_logic_vector(18, 8),
16970 => conv_std_logic_vector(19, 8),
16971 => conv_std_logic_vector(19, 8),
16972 => conv_std_logic_vector(19, 8),
16973 => conv_std_logic_vector(19, 8),
16974 => conv_std_logic_vector(20, 8),
16975 => conv_std_logic_vector(20, 8),
16976 => conv_std_logic_vector(20, 8),
16977 => conv_std_logic_vector(20, 8),
16978 => conv_std_logic_vector(21, 8),
16979 => conv_std_logic_vector(21, 8),
16980 => conv_std_logic_vector(21, 8),
16981 => conv_std_logic_vector(21, 8),
16982 => conv_std_logic_vector(22, 8),
16983 => conv_std_logic_vector(22, 8),
16984 => conv_std_logic_vector(22, 8),
16985 => conv_std_logic_vector(22, 8),
16986 => conv_std_logic_vector(23, 8),
16987 => conv_std_logic_vector(23, 8),
16988 => conv_std_logic_vector(23, 8),
16989 => conv_std_logic_vector(23, 8),
16990 => conv_std_logic_vector(24, 8),
16991 => conv_std_logic_vector(24, 8),
16992 => conv_std_logic_vector(24, 8),
16993 => conv_std_logic_vector(25, 8),
16994 => conv_std_logic_vector(25, 8),
16995 => conv_std_logic_vector(25, 8),
16996 => conv_std_logic_vector(25, 8),
16997 => conv_std_logic_vector(26, 8),
16998 => conv_std_logic_vector(26, 8),
16999 => conv_std_logic_vector(26, 8),
17000 => conv_std_logic_vector(26, 8),
17001 => conv_std_logic_vector(27, 8),
17002 => conv_std_logic_vector(27, 8),
17003 => conv_std_logic_vector(27, 8),
17004 => conv_std_logic_vector(27, 8),
17005 => conv_std_logic_vector(28, 8),
17006 => conv_std_logic_vector(28, 8),
17007 => conv_std_logic_vector(28, 8),
17008 => conv_std_logic_vector(28, 8),
17009 => conv_std_logic_vector(29, 8),
17010 => conv_std_logic_vector(29, 8),
17011 => conv_std_logic_vector(29, 8),
17012 => conv_std_logic_vector(29, 8),
17013 => conv_std_logic_vector(30, 8),
17014 => conv_std_logic_vector(30, 8),
17015 => conv_std_logic_vector(30, 8),
17016 => conv_std_logic_vector(30, 8),
17017 => conv_std_logic_vector(31, 8),
17018 => conv_std_logic_vector(31, 8),
17019 => conv_std_logic_vector(31, 8),
17020 => conv_std_logic_vector(31, 8),
17021 => conv_std_logic_vector(32, 8),
17022 => conv_std_logic_vector(32, 8),
17023 => conv_std_logic_vector(32, 8),
17024 => conv_std_logic_vector(33, 8),
17025 => conv_std_logic_vector(33, 8),
17026 => conv_std_logic_vector(33, 8),
17027 => conv_std_logic_vector(33, 8),
17028 => conv_std_logic_vector(34, 8),
17029 => conv_std_logic_vector(34, 8),
17030 => conv_std_logic_vector(34, 8),
17031 => conv_std_logic_vector(34, 8),
17032 => conv_std_logic_vector(35, 8),
17033 => conv_std_logic_vector(35, 8),
17034 => conv_std_logic_vector(35, 8),
17035 => conv_std_logic_vector(35, 8),
17036 => conv_std_logic_vector(36, 8),
17037 => conv_std_logic_vector(36, 8),
17038 => conv_std_logic_vector(36, 8),
17039 => conv_std_logic_vector(36, 8),
17040 => conv_std_logic_vector(37, 8),
17041 => conv_std_logic_vector(37, 8),
17042 => conv_std_logic_vector(37, 8),
17043 => conv_std_logic_vector(37, 8),
17044 => conv_std_logic_vector(38, 8),
17045 => conv_std_logic_vector(38, 8),
17046 => conv_std_logic_vector(38, 8),
17047 => conv_std_logic_vector(38, 8),
17048 => conv_std_logic_vector(39, 8),
17049 => conv_std_logic_vector(39, 8),
17050 => conv_std_logic_vector(39, 8),
17051 => conv_std_logic_vector(39, 8),
17052 => conv_std_logic_vector(40, 8),
17053 => conv_std_logic_vector(40, 8),
17054 => conv_std_logic_vector(40, 8),
17055 => conv_std_logic_vector(40, 8),
17056 => conv_std_logic_vector(41, 8),
17057 => conv_std_logic_vector(41, 8),
17058 => conv_std_logic_vector(41, 8),
17059 => conv_std_logic_vector(42, 8),
17060 => conv_std_logic_vector(42, 8),
17061 => conv_std_logic_vector(42, 8),
17062 => conv_std_logic_vector(42, 8),
17063 => conv_std_logic_vector(43, 8),
17064 => conv_std_logic_vector(43, 8),
17065 => conv_std_logic_vector(43, 8),
17066 => conv_std_logic_vector(43, 8),
17067 => conv_std_logic_vector(44, 8),
17068 => conv_std_logic_vector(44, 8),
17069 => conv_std_logic_vector(44, 8),
17070 => conv_std_logic_vector(44, 8),
17071 => conv_std_logic_vector(45, 8),
17072 => conv_std_logic_vector(45, 8),
17073 => conv_std_logic_vector(45, 8),
17074 => conv_std_logic_vector(45, 8),
17075 => conv_std_logic_vector(46, 8),
17076 => conv_std_logic_vector(46, 8),
17077 => conv_std_logic_vector(46, 8),
17078 => conv_std_logic_vector(46, 8),
17079 => conv_std_logic_vector(47, 8),
17080 => conv_std_logic_vector(47, 8),
17081 => conv_std_logic_vector(47, 8),
17082 => conv_std_logic_vector(47, 8),
17083 => conv_std_logic_vector(48, 8),
17084 => conv_std_logic_vector(48, 8),
17085 => conv_std_logic_vector(48, 8),
17086 => conv_std_logic_vector(48, 8),
17087 => conv_std_logic_vector(49, 8),
17088 => conv_std_logic_vector(49, 8),
17089 => conv_std_logic_vector(49, 8),
17090 => conv_std_logic_vector(50, 8),
17091 => conv_std_logic_vector(50, 8),
17092 => conv_std_logic_vector(50, 8),
17093 => conv_std_logic_vector(50, 8),
17094 => conv_std_logic_vector(51, 8),
17095 => conv_std_logic_vector(51, 8),
17096 => conv_std_logic_vector(51, 8),
17097 => conv_std_logic_vector(51, 8),
17098 => conv_std_logic_vector(52, 8),
17099 => conv_std_logic_vector(52, 8),
17100 => conv_std_logic_vector(52, 8),
17101 => conv_std_logic_vector(52, 8),
17102 => conv_std_logic_vector(53, 8),
17103 => conv_std_logic_vector(53, 8),
17104 => conv_std_logic_vector(53, 8),
17105 => conv_std_logic_vector(53, 8),
17106 => conv_std_logic_vector(54, 8),
17107 => conv_std_logic_vector(54, 8),
17108 => conv_std_logic_vector(54, 8),
17109 => conv_std_logic_vector(54, 8),
17110 => conv_std_logic_vector(55, 8),
17111 => conv_std_logic_vector(55, 8),
17112 => conv_std_logic_vector(55, 8),
17113 => conv_std_logic_vector(55, 8),
17114 => conv_std_logic_vector(56, 8),
17115 => conv_std_logic_vector(56, 8),
17116 => conv_std_logic_vector(56, 8),
17117 => conv_std_logic_vector(56, 8),
17118 => conv_std_logic_vector(57, 8),
17119 => conv_std_logic_vector(57, 8),
17120 => conv_std_logic_vector(57, 8),
17121 => conv_std_logic_vector(58, 8),
17122 => conv_std_logic_vector(58, 8),
17123 => conv_std_logic_vector(58, 8),
17124 => conv_std_logic_vector(58, 8),
17125 => conv_std_logic_vector(59, 8),
17126 => conv_std_logic_vector(59, 8),
17127 => conv_std_logic_vector(59, 8),
17128 => conv_std_logic_vector(59, 8),
17129 => conv_std_logic_vector(60, 8),
17130 => conv_std_logic_vector(60, 8),
17131 => conv_std_logic_vector(60, 8),
17132 => conv_std_logic_vector(60, 8),
17133 => conv_std_logic_vector(61, 8),
17134 => conv_std_logic_vector(61, 8),
17135 => conv_std_logic_vector(61, 8),
17136 => conv_std_logic_vector(61, 8),
17137 => conv_std_logic_vector(62, 8),
17138 => conv_std_logic_vector(62, 8),
17139 => conv_std_logic_vector(62, 8),
17140 => conv_std_logic_vector(62, 8),
17141 => conv_std_logic_vector(63, 8),
17142 => conv_std_logic_vector(63, 8),
17143 => conv_std_logic_vector(63, 8),
17144 => conv_std_logic_vector(63, 8),
17145 => conv_std_logic_vector(64, 8),
17146 => conv_std_logic_vector(64, 8),
17147 => conv_std_logic_vector(64, 8),
17148 => conv_std_logic_vector(64, 8),
17149 => conv_std_logic_vector(65, 8),
17150 => conv_std_logic_vector(65, 8),
17151 => conv_std_logic_vector(65, 8),
17152 => conv_std_logic_vector(0, 8),
17153 => conv_std_logic_vector(0, 8),
17154 => conv_std_logic_vector(0, 8),
17155 => conv_std_logic_vector(0, 8),
17156 => conv_std_logic_vector(1, 8),
17157 => conv_std_logic_vector(1, 8),
17158 => conv_std_logic_vector(1, 8),
17159 => conv_std_logic_vector(1, 8),
17160 => conv_std_logic_vector(2, 8),
17161 => conv_std_logic_vector(2, 8),
17162 => conv_std_logic_vector(2, 8),
17163 => conv_std_logic_vector(2, 8),
17164 => conv_std_logic_vector(3, 8),
17165 => conv_std_logic_vector(3, 8),
17166 => conv_std_logic_vector(3, 8),
17167 => conv_std_logic_vector(3, 8),
17168 => conv_std_logic_vector(4, 8),
17169 => conv_std_logic_vector(4, 8),
17170 => conv_std_logic_vector(4, 8),
17171 => conv_std_logic_vector(4, 8),
17172 => conv_std_logic_vector(5, 8),
17173 => conv_std_logic_vector(5, 8),
17174 => conv_std_logic_vector(5, 8),
17175 => conv_std_logic_vector(6, 8),
17176 => conv_std_logic_vector(6, 8),
17177 => conv_std_logic_vector(6, 8),
17178 => conv_std_logic_vector(6, 8),
17179 => conv_std_logic_vector(7, 8),
17180 => conv_std_logic_vector(7, 8),
17181 => conv_std_logic_vector(7, 8),
17182 => conv_std_logic_vector(7, 8),
17183 => conv_std_logic_vector(8, 8),
17184 => conv_std_logic_vector(8, 8),
17185 => conv_std_logic_vector(8, 8),
17186 => conv_std_logic_vector(8, 8),
17187 => conv_std_logic_vector(9, 8),
17188 => conv_std_logic_vector(9, 8),
17189 => conv_std_logic_vector(9, 8),
17190 => conv_std_logic_vector(9, 8),
17191 => conv_std_logic_vector(10, 8),
17192 => conv_std_logic_vector(10, 8),
17193 => conv_std_logic_vector(10, 8),
17194 => conv_std_logic_vector(10, 8),
17195 => conv_std_logic_vector(11, 8),
17196 => conv_std_logic_vector(11, 8),
17197 => conv_std_logic_vector(11, 8),
17198 => conv_std_logic_vector(12, 8),
17199 => conv_std_logic_vector(12, 8),
17200 => conv_std_logic_vector(12, 8),
17201 => conv_std_logic_vector(12, 8),
17202 => conv_std_logic_vector(13, 8),
17203 => conv_std_logic_vector(13, 8),
17204 => conv_std_logic_vector(13, 8),
17205 => conv_std_logic_vector(13, 8),
17206 => conv_std_logic_vector(14, 8),
17207 => conv_std_logic_vector(14, 8),
17208 => conv_std_logic_vector(14, 8),
17209 => conv_std_logic_vector(14, 8),
17210 => conv_std_logic_vector(15, 8),
17211 => conv_std_logic_vector(15, 8),
17212 => conv_std_logic_vector(15, 8),
17213 => conv_std_logic_vector(15, 8),
17214 => conv_std_logic_vector(16, 8),
17215 => conv_std_logic_vector(16, 8),
17216 => conv_std_logic_vector(16, 8),
17217 => conv_std_logic_vector(17, 8),
17218 => conv_std_logic_vector(17, 8),
17219 => conv_std_logic_vector(17, 8),
17220 => conv_std_logic_vector(17, 8),
17221 => conv_std_logic_vector(18, 8),
17222 => conv_std_logic_vector(18, 8),
17223 => conv_std_logic_vector(18, 8),
17224 => conv_std_logic_vector(18, 8),
17225 => conv_std_logic_vector(19, 8),
17226 => conv_std_logic_vector(19, 8),
17227 => conv_std_logic_vector(19, 8),
17228 => conv_std_logic_vector(19, 8),
17229 => conv_std_logic_vector(20, 8),
17230 => conv_std_logic_vector(20, 8),
17231 => conv_std_logic_vector(20, 8),
17232 => conv_std_logic_vector(20, 8),
17233 => conv_std_logic_vector(21, 8),
17234 => conv_std_logic_vector(21, 8),
17235 => conv_std_logic_vector(21, 8),
17236 => conv_std_logic_vector(21, 8),
17237 => conv_std_logic_vector(22, 8),
17238 => conv_std_logic_vector(22, 8),
17239 => conv_std_logic_vector(22, 8),
17240 => conv_std_logic_vector(23, 8),
17241 => conv_std_logic_vector(23, 8),
17242 => conv_std_logic_vector(23, 8),
17243 => conv_std_logic_vector(23, 8),
17244 => conv_std_logic_vector(24, 8),
17245 => conv_std_logic_vector(24, 8),
17246 => conv_std_logic_vector(24, 8),
17247 => conv_std_logic_vector(24, 8),
17248 => conv_std_logic_vector(25, 8),
17249 => conv_std_logic_vector(25, 8),
17250 => conv_std_logic_vector(25, 8),
17251 => conv_std_logic_vector(25, 8),
17252 => conv_std_logic_vector(26, 8),
17253 => conv_std_logic_vector(26, 8),
17254 => conv_std_logic_vector(26, 8),
17255 => conv_std_logic_vector(26, 8),
17256 => conv_std_logic_vector(27, 8),
17257 => conv_std_logic_vector(27, 8),
17258 => conv_std_logic_vector(27, 8),
17259 => conv_std_logic_vector(28, 8),
17260 => conv_std_logic_vector(28, 8),
17261 => conv_std_logic_vector(28, 8),
17262 => conv_std_logic_vector(28, 8),
17263 => conv_std_logic_vector(29, 8),
17264 => conv_std_logic_vector(29, 8),
17265 => conv_std_logic_vector(29, 8),
17266 => conv_std_logic_vector(29, 8),
17267 => conv_std_logic_vector(30, 8),
17268 => conv_std_logic_vector(30, 8),
17269 => conv_std_logic_vector(30, 8),
17270 => conv_std_logic_vector(30, 8),
17271 => conv_std_logic_vector(31, 8),
17272 => conv_std_logic_vector(31, 8),
17273 => conv_std_logic_vector(31, 8),
17274 => conv_std_logic_vector(31, 8),
17275 => conv_std_logic_vector(32, 8),
17276 => conv_std_logic_vector(32, 8),
17277 => conv_std_logic_vector(32, 8),
17278 => conv_std_logic_vector(32, 8),
17279 => conv_std_logic_vector(33, 8),
17280 => conv_std_logic_vector(33, 8),
17281 => conv_std_logic_vector(33, 8),
17282 => conv_std_logic_vector(34, 8),
17283 => conv_std_logic_vector(34, 8),
17284 => conv_std_logic_vector(34, 8),
17285 => conv_std_logic_vector(34, 8),
17286 => conv_std_logic_vector(35, 8),
17287 => conv_std_logic_vector(35, 8),
17288 => conv_std_logic_vector(35, 8),
17289 => conv_std_logic_vector(35, 8),
17290 => conv_std_logic_vector(36, 8),
17291 => conv_std_logic_vector(36, 8),
17292 => conv_std_logic_vector(36, 8),
17293 => conv_std_logic_vector(36, 8),
17294 => conv_std_logic_vector(37, 8),
17295 => conv_std_logic_vector(37, 8),
17296 => conv_std_logic_vector(37, 8),
17297 => conv_std_logic_vector(37, 8),
17298 => conv_std_logic_vector(38, 8),
17299 => conv_std_logic_vector(38, 8),
17300 => conv_std_logic_vector(38, 8),
17301 => conv_std_logic_vector(38, 8),
17302 => conv_std_logic_vector(39, 8),
17303 => conv_std_logic_vector(39, 8),
17304 => conv_std_logic_vector(39, 8),
17305 => conv_std_logic_vector(40, 8),
17306 => conv_std_logic_vector(40, 8),
17307 => conv_std_logic_vector(40, 8),
17308 => conv_std_logic_vector(40, 8),
17309 => conv_std_logic_vector(41, 8),
17310 => conv_std_logic_vector(41, 8),
17311 => conv_std_logic_vector(41, 8),
17312 => conv_std_logic_vector(41, 8),
17313 => conv_std_logic_vector(42, 8),
17314 => conv_std_logic_vector(42, 8),
17315 => conv_std_logic_vector(42, 8),
17316 => conv_std_logic_vector(42, 8),
17317 => conv_std_logic_vector(43, 8),
17318 => conv_std_logic_vector(43, 8),
17319 => conv_std_logic_vector(43, 8),
17320 => conv_std_logic_vector(43, 8),
17321 => conv_std_logic_vector(44, 8),
17322 => conv_std_logic_vector(44, 8),
17323 => conv_std_logic_vector(44, 8),
17324 => conv_std_logic_vector(45, 8),
17325 => conv_std_logic_vector(45, 8),
17326 => conv_std_logic_vector(45, 8),
17327 => conv_std_logic_vector(45, 8),
17328 => conv_std_logic_vector(46, 8),
17329 => conv_std_logic_vector(46, 8),
17330 => conv_std_logic_vector(46, 8),
17331 => conv_std_logic_vector(46, 8),
17332 => conv_std_logic_vector(47, 8),
17333 => conv_std_logic_vector(47, 8),
17334 => conv_std_logic_vector(47, 8),
17335 => conv_std_logic_vector(47, 8),
17336 => conv_std_logic_vector(48, 8),
17337 => conv_std_logic_vector(48, 8),
17338 => conv_std_logic_vector(48, 8),
17339 => conv_std_logic_vector(48, 8),
17340 => conv_std_logic_vector(49, 8),
17341 => conv_std_logic_vector(49, 8),
17342 => conv_std_logic_vector(49, 8),
17343 => conv_std_logic_vector(49, 8),
17344 => conv_std_logic_vector(50, 8),
17345 => conv_std_logic_vector(50, 8),
17346 => conv_std_logic_vector(50, 8),
17347 => conv_std_logic_vector(51, 8),
17348 => conv_std_logic_vector(51, 8),
17349 => conv_std_logic_vector(51, 8),
17350 => conv_std_logic_vector(51, 8),
17351 => conv_std_logic_vector(52, 8),
17352 => conv_std_logic_vector(52, 8),
17353 => conv_std_logic_vector(52, 8),
17354 => conv_std_logic_vector(52, 8),
17355 => conv_std_logic_vector(53, 8),
17356 => conv_std_logic_vector(53, 8),
17357 => conv_std_logic_vector(53, 8),
17358 => conv_std_logic_vector(53, 8),
17359 => conv_std_logic_vector(54, 8),
17360 => conv_std_logic_vector(54, 8),
17361 => conv_std_logic_vector(54, 8),
17362 => conv_std_logic_vector(54, 8),
17363 => conv_std_logic_vector(55, 8),
17364 => conv_std_logic_vector(55, 8),
17365 => conv_std_logic_vector(55, 8),
17366 => conv_std_logic_vector(56, 8),
17367 => conv_std_logic_vector(56, 8),
17368 => conv_std_logic_vector(56, 8),
17369 => conv_std_logic_vector(56, 8),
17370 => conv_std_logic_vector(57, 8),
17371 => conv_std_logic_vector(57, 8),
17372 => conv_std_logic_vector(57, 8),
17373 => conv_std_logic_vector(57, 8),
17374 => conv_std_logic_vector(58, 8),
17375 => conv_std_logic_vector(58, 8),
17376 => conv_std_logic_vector(58, 8),
17377 => conv_std_logic_vector(58, 8),
17378 => conv_std_logic_vector(59, 8),
17379 => conv_std_logic_vector(59, 8),
17380 => conv_std_logic_vector(59, 8),
17381 => conv_std_logic_vector(59, 8),
17382 => conv_std_logic_vector(60, 8),
17383 => conv_std_logic_vector(60, 8),
17384 => conv_std_logic_vector(60, 8),
17385 => conv_std_logic_vector(60, 8),
17386 => conv_std_logic_vector(61, 8),
17387 => conv_std_logic_vector(61, 8),
17388 => conv_std_logic_vector(61, 8),
17389 => conv_std_logic_vector(62, 8),
17390 => conv_std_logic_vector(62, 8),
17391 => conv_std_logic_vector(62, 8),
17392 => conv_std_logic_vector(62, 8),
17393 => conv_std_logic_vector(63, 8),
17394 => conv_std_logic_vector(63, 8),
17395 => conv_std_logic_vector(63, 8),
17396 => conv_std_logic_vector(63, 8),
17397 => conv_std_logic_vector(64, 8),
17398 => conv_std_logic_vector(64, 8),
17399 => conv_std_logic_vector(64, 8),
17400 => conv_std_logic_vector(64, 8),
17401 => conv_std_logic_vector(65, 8),
17402 => conv_std_logic_vector(65, 8),
17403 => conv_std_logic_vector(65, 8),
17404 => conv_std_logic_vector(65, 8),
17405 => conv_std_logic_vector(66, 8),
17406 => conv_std_logic_vector(66, 8),
17407 => conv_std_logic_vector(66, 8),
17408 => conv_std_logic_vector(0, 8),
17409 => conv_std_logic_vector(0, 8),
17410 => conv_std_logic_vector(0, 8),
17411 => conv_std_logic_vector(0, 8),
17412 => conv_std_logic_vector(1, 8),
17413 => conv_std_logic_vector(1, 8),
17414 => conv_std_logic_vector(1, 8),
17415 => conv_std_logic_vector(1, 8),
17416 => conv_std_logic_vector(2, 8),
17417 => conv_std_logic_vector(2, 8),
17418 => conv_std_logic_vector(2, 8),
17419 => conv_std_logic_vector(2, 8),
17420 => conv_std_logic_vector(3, 8),
17421 => conv_std_logic_vector(3, 8),
17422 => conv_std_logic_vector(3, 8),
17423 => conv_std_logic_vector(3, 8),
17424 => conv_std_logic_vector(4, 8),
17425 => conv_std_logic_vector(4, 8),
17426 => conv_std_logic_vector(4, 8),
17427 => conv_std_logic_vector(5, 8),
17428 => conv_std_logic_vector(5, 8),
17429 => conv_std_logic_vector(5, 8),
17430 => conv_std_logic_vector(5, 8),
17431 => conv_std_logic_vector(6, 8),
17432 => conv_std_logic_vector(6, 8),
17433 => conv_std_logic_vector(6, 8),
17434 => conv_std_logic_vector(6, 8),
17435 => conv_std_logic_vector(7, 8),
17436 => conv_std_logic_vector(7, 8),
17437 => conv_std_logic_vector(7, 8),
17438 => conv_std_logic_vector(7, 8),
17439 => conv_std_logic_vector(8, 8),
17440 => conv_std_logic_vector(8, 8),
17441 => conv_std_logic_vector(8, 8),
17442 => conv_std_logic_vector(9, 8),
17443 => conv_std_logic_vector(9, 8),
17444 => conv_std_logic_vector(9, 8),
17445 => conv_std_logic_vector(9, 8),
17446 => conv_std_logic_vector(10, 8),
17447 => conv_std_logic_vector(10, 8),
17448 => conv_std_logic_vector(10, 8),
17449 => conv_std_logic_vector(10, 8),
17450 => conv_std_logic_vector(11, 8),
17451 => conv_std_logic_vector(11, 8),
17452 => conv_std_logic_vector(11, 8),
17453 => conv_std_logic_vector(11, 8),
17454 => conv_std_logic_vector(12, 8),
17455 => conv_std_logic_vector(12, 8),
17456 => conv_std_logic_vector(12, 8),
17457 => conv_std_logic_vector(13, 8),
17458 => conv_std_logic_vector(13, 8),
17459 => conv_std_logic_vector(13, 8),
17460 => conv_std_logic_vector(13, 8),
17461 => conv_std_logic_vector(14, 8),
17462 => conv_std_logic_vector(14, 8),
17463 => conv_std_logic_vector(14, 8),
17464 => conv_std_logic_vector(14, 8),
17465 => conv_std_logic_vector(15, 8),
17466 => conv_std_logic_vector(15, 8),
17467 => conv_std_logic_vector(15, 8),
17468 => conv_std_logic_vector(15, 8),
17469 => conv_std_logic_vector(16, 8),
17470 => conv_std_logic_vector(16, 8),
17471 => conv_std_logic_vector(16, 8),
17472 => conv_std_logic_vector(17, 8),
17473 => conv_std_logic_vector(17, 8),
17474 => conv_std_logic_vector(17, 8),
17475 => conv_std_logic_vector(17, 8),
17476 => conv_std_logic_vector(18, 8),
17477 => conv_std_logic_vector(18, 8),
17478 => conv_std_logic_vector(18, 8),
17479 => conv_std_logic_vector(18, 8),
17480 => conv_std_logic_vector(19, 8),
17481 => conv_std_logic_vector(19, 8),
17482 => conv_std_logic_vector(19, 8),
17483 => conv_std_logic_vector(19, 8),
17484 => conv_std_logic_vector(20, 8),
17485 => conv_std_logic_vector(20, 8),
17486 => conv_std_logic_vector(20, 8),
17487 => conv_std_logic_vector(20, 8),
17488 => conv_std_logic_vector(21, 8),
17489 => conv_std_logic_vector(21, 8),
17490 => conv_std_logic_vector(21, 8),
17491 => conv_std_logic_vector(22, 8),
17492 => conv_std_logic_vector(22, 8),
17493 => conv_std_logic_vector(22, 8),
17494 => conv_std_logic_vector(22, 8),
17495 => conv_std_logic_vector(23, 8),
17496 => conv_std_logic_vector(23, 8),
17497 => conv_std_logic_vector(23, 8),
17498 => conv_std_logic_vector(23, 8),
17499 => conv_std_logic_vector(24, 8),
17500 => conv_std_logic_vector(24, 8),
17501 => conv_std_logic_vector(24, 8),
17502 => conv_std_logic_vector(24, 8),
17503 => conv_std_logic_vector(25, 8),
17504 => conv_std_logic_vector(25, 8),
17505 => conv_std_logic_vector(25, 8),
17506 => conv_std_logic_vector(26, 8),
17507 => conv_std_logic_vector(26, 8),
17508 => conv_std_logic_vector(26, 8),
17509 => conv_std_logic_vector(26, 8),
17510 => conv_std_logic_vector(27, 8),
17511 => conv_std_logic_vector(27, 8),
17512 => conv_std_logic_vector(27, 8),
17513 => conv_std_logic_vector(27, 8),
17514 => conv_std_logic_vector(28, 8),
17515 => conv_std_logic_vector(28, 8),
17516 => conv_std_logic_vector(28, 8),
17517 => conv_std_logic_vector(28, 8),
17518 => conv_std_logic_vector(29, 8),
17519 => conv_std_logic_vector(29, 8),
17520 => conv_std_logic_vector(29, 8),
17521 => conv_std_logic_vector(30, 8),
17522 => conv_std_logic_vector(30, 8),
17523 => conv_std_logic_vector(30, 8),
17524 => conv_std_logic_vector(30, 8),
17525 => conv_std_logic_vector(31, 8),
17526 => conv_std_logic_vector(31, 8),
17527 => conv_std_logic_vector(31, 8),
17528 => conv_std_logic_vector(31, 8),
17529 => conv_std_logic_vector(32, 8),
17530 => conv_std_logic_vector(32, 8),
17531 => conv_std_logic_vector(32, 8),
17532 => conv_std_logic_vector(32, 8),
17533 => conv_std_logic_vector(33, 8),
17534 => conv_std_logic_vector(33, 8),
17535 => conv_std_logic_vector(33, 8),
17536 => conv_std_logic_vector(34, 8),
17537 => conv_std_logic_vector(34, 8),
17538 => conv_std_logic_vector(34, 8),
17539 => conv_std_logic_vector(34, 8),
17540 => conv_std_logic_vector(35, 8),
17541 => conv_std_logic_vector(35, 8),
17542 => conv_std_logic_vector(35, 8),
17543 => conv_std_logic_vector(35, 8),
17544 => conv_std_logic_vector(36, 8),
17545 => conv_std_logic_vector(36, 8),
17546 => conv_std_logic_vector(36, 8),
17547 => conv_std_logic_vector(36, 8),
17548 => conv_std_logic_vector(37, 8),
17549 => conv_std_logic_vector(37, 8),
17550 => conv_std_logic_vector(37, 8),
17551 => conv_std_logic_vector(37, 8),
17552 => conv_std_logic_vector(38, 8),
17553 => conv_std_logic_vector(38, 8),
17554 => conv_std_logic_vector(38, 8),
17555 => conv_std_logic_vector(39, 8),
17556 => conv_std_logic_vector(39, 8),
17557 => conv_std_logic_vector(39, 8),
17558 => conv_std_logic_vector(39, 8),
17559 => conv_std_logic_vector(40, 8),
17560 => conv_std_logic_vector(40, 8),
17561 => conv_std_logic_vector(40, 8),
17562 => conv_std_logic_vector(40, 8),
17563 => conv_std_logic_vector(41, 8),
17564 => conv_std_logic_vector(41, 8),
17565 => conv_std_logic_vector(41, 8),
17566 => conv_std_logic_vector(41, 8),
17567 => conv_std_logic_vector(42, 8),
17568 => conv_std_logic_vector(42, 8),
17569 => conv_std_logic_vector(42, 8),
17570 => conv_std_logic_vector(43, 8),
17571 => conv_std_logic_vector(43, 8),
17572 => conv_std_logic_vector(43, 8),
17573 => conv_std_logic_vector(43, 8),
17574 => conv_std_logic_vector(44, 8),
17575 => conv_std_logic_vector(44, 8),
17576 => conv_std_logic_vector(44, 8),
17577 => conv_std_logic_vector(44, 8),
17578 => conv_std_logic_vector(45, 8),
17579 => conv_std_logic_vector(45, 8),
17580 => conv_std_logic_vector(45, 8),
17581 => conv_std_logic_vector(45, 8),
17582 => conv_std_logic_vector(46, 8),
17583 => conv_std_logic_vector(46, 8),
17584 => conv_std_logic_vector(46, 8),
17585 => conv_std_logic_vector(47, 8),
17586 => conv_std_logic_vector(47, 8),
17587 => conv_std_logic_vector(47, 8),
17588 => conv_std_logic_vector(47, 8),
17589 => conv_std_logic_vector(48, 8),
17590 => conv_std_logic_vector(48, 8),
17591 => conv_std_logic_vector(48, 8),
17592 => conv_std_logic_vector(48, 8),
17593 => conv_std_logic_vector(49, 8),
17594 => conv_std_logic_vector(49, 8),
17595 => conv_std_logic_vector(49, 8),
17596 => conv_std_logic_vector(49, 8),
17597 => conv_std_logic_vector(50, 8),
17598 => conv_std_logic_vector(50, 8),
17599 => conv_std_logic_vector(50, 8),
17600 => conv_std_logic_vector(51, 8),
17601 => conv_std_logic_vector(51, 8),
17602 => conv_std_logic_vector(51, 8),
17603 => conv_std_logic_vector(51, 8),
17604 => conv_std_logic_vector(52, 8),
17605 => conv_std_logic_vector(52, 8),
17606 => conv_std_logic_vector(52, 8),
17607 => conv_std_logic_vector(52, 8),
17608 => conv_std_logic_vector(53, 8),
17609 => conv_std_logic_vector(53, 8),
17610 => conv_std_logic_vector(53, 8),
17611 => conv_std_logic_vector(53, 8),
17612 => conv_std_logic_vector(54, 8),
17613 => conv_std_logic_vector(54, 8),
17614 => conv_std_logic_vector(54, 8),
17615 => conv_std_logic_vector(54, 8),
17616 => conv_std_logic_vector(55, 8),
17617 => conv_std_logic_vector(55, 8),
17618 => conv_std_logic_vector(55, 8),
17619 => conv_std_logic_vector(56, 8),
17620 => conv_std_logic_vector(56, 8),
17621 => conv_std_logic_vector(56, 8),
17622 => conv_std_logic_vector(56, 8),
17623 => conv_std_logic_vector(57, 8),
17624 => conv_std_logic_vector(57, 8),
17625 => conv_std_logic_vector(57, 8),
17626 => conv_std_logic_vector(57, 8),
17627 => conv_std_logic_vector(58, 8),
17628 => conv_std_logic_vector(58, 8),
17629 => conv_std_logic_vector(58, 8),
17630 => conv_std_logic_vector(58, 8),
17631 => conv_std_logic_vector(59, 8),
17632 => conv_std_logic_vector(59, 8),
17633 => conv_std_logic_vector(59, 8),
17634 => conv_std_logic_vector(60, 8),
17635 => conv_std_logic_vector(60, 8),
17636 => conv_std_logic_vector(60, 8),
17637 => conv_std_logic_vector(60, 8),
17638 => conv_std_logic_vector(61, 8),
17639 => conv_std_logic_vector(61, 8),
17640 => conv_std_logic_vector(61, 8),
17641 => conv_std_logic_vector(61, 8),
17642 => conv_std_logic_vector(62, 8),
17643 => conv_std_logic_vector(62, 8),
17644 => conv_std_logic_vector(62, 8),
17645 => conv_std_logic_vector(62, 8),
17646 => conv_std_logic_vector(63, 8),
17647 => conv_std_logic_vector(63, 8),
17648 => conv_std_logic_vector(63, 8),
17649 => conv_std_logic_vector(64, 8),
17650 => conv_std_logic_vector(64, 8),
17651 => conv_std_logic_vector(64, 8),
17652 => conv_std_logic_vector(64, 8),
17653 => conv_std_logic_vector(65, 8),
17654 => conv_std_logic_vector(65, 8),
17655 => conv_std_logic_vector(65, 8),
17656 => conv_std_logic_vector(65, 8),
17657 => conv_std_logic_vector(66, 8),
17658 => conv_std_logic_vector(66, 8),
17659 => conv_std_logic_vector(66, 8),
17660 => conv_std_logic_vector(66, 8),
17661 => conv_std_logic_vector(67, 8),
17662 => conv_std_logic_vector(67, 8),
17663 => conv_std_logic_vector(67, 8),
17664 => conv_std_logic_vector(0, 8),
17665 => conv_std_logic_vector(0, 8),
17666 => conv_std_logic_vector(0, 8),
17667 => conv_std_logic_vector(0, 8),
17668 => conv_std_logic_vector(1, 8),
17669 => conv_std_logic_vector(1, 8),
17670 => conv_std_logic_vector(1, 8),
17671 => conv_std_logic_vector(1, 8),
17672 => conv_std_logic_vector(2, 8),
17673 => conv_std_logic_vector(2, 8),
17674 => conv_std_logic_vector(2, 8),
17675 => conv_std_logic_vector(2, 8),
17676 => conv_std_logic_vector(3, 8),
17677 => conv_std_logic_vector(3, 8),
17678 => conv_std_logic_vector(3, 8),
17679 => conv_std_logic_vector(4, 8),
17680 => conv_std_logic_vector(4, 8),
17681 => conv_std_logic_vector(4, 8),
17682 => conv_std_logic_vector(4, 8),
17683 => conv_std_logic_vector(5, 8),
17684 => conv_std_logic_vector(5, 8),
17685 => conv_std_logic_vector(5, 8),
17686 => conv_std_logic_vector(5, 8),
17687 => conv_std_logic_vector(6, 8),
17688 => conv_std_logic_vector(6, 8),
17689 => conv_std_logic_vector(6, 8),
17690 => conv_std_logic_vector(7, 8),
17691 => conv_std_logic_vector(7, 8),
17692 => conv_std_logic_vector(7, 8),
17693 => conv_std_logic_vector(7, 8),
17694 => conv_std_logic_vector(8, 8),
17695 => conv_std_logic_vector(8, 8),
17696 => conv_std_logic_vector(8, 8),
17697 => conv_std_logic_vector(8, 8),
17698 => conv_std_logic_vector(9, 8),
17699 => conv_std_logic_vector(9, 8),
17700 => conv_std_logic_vector(9, 8),
17701 => conv_std_logic_vector(9, 8),
17702 => conv_std_logic_vector(10, 8),
17703 => conv_std_logic_vector(10, 8),
17704 => conv_std_logic_vector(10, 8),
17705 => conv_std_logic_vector(11, 8),
17706 => conv_std_logic_vector(11, 8),
17707 => conv_std_logic_vector(11, 8),
17708 => conv_std_logic_vector(11, 8),
17709 => conv_std_logic_vector(12, 8),
17710 => conv_std_logic_vector(12, 8),
17711 => conv_std_logic_vector(12, 8),
17712 => conv_std_logic_vector(12, 8),
17713 => conv_std_logic_vector(13, 8),
17714 => conv_std_logic_vector(13, 8),
17715 => conv_std_logic_vector(13, 8),
17716 => conv_std_logic_vector(14, 8),
17717 => conv_std_logic_vector(14, 8),
17718 => conv_std_logic_vector(14, 8),
17719 => conv_std_logic_vector(14, 8),
17720 => conv_std_logic_vector(15, 8),
17721 => conv_std_logic_vector(15, 8),
17722 => conv_std_logic_vector(15, 8),
17723 => conv_std_logic_vector(15, 8),
17724 => conv_std_logic_vector(16, 8),
17725 => conv_std_logic_vector(16, 8),
17726 => conv_std_logic_vector(16, 8),
17727 => conv_std_logic_vector(16, 8),
17728 => conv_std_logic_vector(17, 8),
17729 => conv_std_logic_vector(17, 8),
17730 => conv_std_logic_vector(17, 8),
17731 => conv_std_logic_vector(18, 8),
17732 => conv_std_logic_vector(18, 8),
17733 => conv_std_logic_vector(18, 8),
17734 => conv_std_logic_vector(18, 8),
17735 => conv_std_logic_vector(19, 8),
17736 => conv_std_logic_vector(19, 8),
17737 => conv_std_logic_vector(19, 8),
17738 => conv_std_logic_vector(19, 8),
17739 => conv_std_logic_vector(20, 8),
17740 => conv_std_logic_vector(20, 8),
17741 => conv_std_logic_vector(20, 8),
17742 => conv_std_logic_vector(21, 8),
17743 => conv_std_logic_vector(21, 8),
17744 => conv_std_logic_vector(21, 8),
17745 => conv_std_logic_vector(21, 8),
17746 => conv_std_logic_vector(22, 8),
17747 => conv_std_logic_vector(22, 8),
17748 => conv_std_logic_vector(22, 8),
17749 => conv_std_logic_vector(22, 8),
17750 => conv_std_logic_vector(23, 8),
17751 => conv_std_logic_vector(23, 8),
17752 => conv_std_logic_vector(23, 8),
17753 => conv_std_logic_vector(23, 8),
17754 => conv_std_logic_vector(24, 8),
17755 => conv_std_logic_vector(24, 8),
17756 => conv_std_logic_vector(24, 8),
17757 => conv_std_logic_vector(25, 8),
17758 => conv_std_logic_vector(25, 8),
17759 => conv_std_logic_vector(25, 8),
17760 => conv_std_logic_vector(25, 8),
17761 => conv_std_logic_vector(26, 8),
17762 => conv_std_logic_vector(26, 8),
17763 => conv_std_logic_vector(26, 8),
17764 => conv_std_logic_vector(26, 8),
17765 => conv_std_logic_vector(27, 8),
17766 => conv_std_logic_vector(27, 8),
17767 => conv_std_logic_vector(27, 8),
17768 => conv_std_logic_vector(28, 8),
17769 => conv_std_logic_vector(28, 8),
17770 => conv_std_logic_vector(28, 8),
17771 => conv_std_logic_vector(28, 8),
17772 => conv_std_logic_vector(29, 8),
17773 => conv_std_logic_vector(29, 8),
17774 => conv_std_logic_vector(29, 8),
17775 => conv_std_logic_vector(29, 8),
17776 => conv_std_logic_vector(30, 8),
17777 => conv_std_logic_vector(30, 8),
17778 => conv_std_logic_vector(30, 8),
17779 => conv_std_logic_vector(30, 8),
17780 => conv_std_logic_vector(31, 8),
17781 => conv_std_logic_vector(31, 8),
17782 => conv_std_logic_vector(31, 8),
17783 => conv_std_logic_vector(32, 8),
17784 => conv_std_logic_vector(32, 8),
17785 => conv_std_logic_vector(32, 8),
17786 => conv_std_logic_vector(32, 8),
17787 => conv_std_logic_vector(33, 8),
17788 => conv_std_logic_vector(33, 8),
17789 => conv_std_logic_vector(33, 8),
17790 => conv_std_logic_vector(33, 8),
17791 => conv_std_logic_vector(34, 8),
17792 => conv_std_logic_vector(34, 8),
17793 => conv_std_logic_vector(34, 8),
17794 => conv_std_logic_vector(35, 8),
17795 => conv_std_logic_vector(35, 8),
17796 => conv_std_logic_vector(35, 8),
17797 => conv_std_logic_vector(35, 8),
17798 => conv_std_logic_vector(36, 8),
17799 => conv_std_logic_vector(36, 8),
17800 => conv_std_logic_vector(36, 8),
17801 => conv_std_logic_vector(36, 8),
17802 => conv_std_logic_vector(37, 8),
17803 => conv_std_logic_vector(37, 8),
17804 => conv_std_logic_vector(37, 8),
17805 => conv_std_logic_vector(38, 8),
17806 => conv_std_logic_vector(38, 8),
17807 => conv_std_logic_vector(38, 8),
17808 => conv_std_logic_vector(38, 8),
17809 => conv_std_logic_vector(39, 8),
17810 => conv_std_logic_vector(39, 8),
17811 => conv_std_logic_vector(39, 8),
17812 => conv_std_logic_vector(39, 8),
17813 => conv_std_logic_vector(40, 8),
17814 => conv_std_logic_vector(40, 8),
17815 => conv_std_logic_vector(40, 8),
17816 => conv_std_logic_vector(40, 8),
17817 => conv_std_logic_vector(41, 8),
17818 => conv_std_logic_vector(41, 8),
17819 => conv_std_logic_vector(41, 8),
17820 => conv_std_logic_vector(42, 8),
17821 => conv_std_logic_vector(42, 8),
17822 => conv_std_logic_vector(42, 8),
17823 => conv_std_logic_vector(42, 8),
17824 => conv_std_logic_vector(43, 8),
17825 => conv_std_logic_vector(43, 8),
17826 => conv_std_logic_vector(43, 8),
17827 => conv_std_logic_vector(43, 8),
17828 => conv_std_logic_vector(44, 8),
17829 => conv_std_logic_vector(44, 8),
17830 => conv_std_logic_vector(44, 8),
17831 => conv_std_logic_vector(45, 8),
17832 => conv_std_logic_vector(45, 8),
17833 => conv_std_logic_vector(45, 8),
17834 => conv_std_logic_vector(45, 8),
17835 => conv_std_logic_vector(46, 8),
17836 => conv_std_logic_vector(46, 8),
17837 => conv_std_logic_vector(46, 8),
17838 => conv_std_logic_vector(46, 8),
17839 => conv_std_logic_vector(47, 8),
17840 => conv_std_logic_vector(47, 8),
17841 => conv_std_logic_vector(47, 8),
17842 => conv_std_logic_vector(47, 8),
17843 => conv_std_logic_vector(48, 8),
17844 => conv_std_logic_vector(48, 8),
17845 => conv_std_logic_vector(48, 8),
17846 => conv_std_logic_vector(49, 8),
17847 => conv_std_logic_vector(49, 8),
17848 => conv_std_logic_vector(49, 8),
17849 => conv_std_logic_vector(49, 8),
17850 => conv_std_logic_vector(50, 8),
17851 => conv_std_logic_vector(50, 8),
17852 => conv_std_logic_vector(50, 8),
17853 => conv_std_logic_vector(50, 8),
17854 => conv_std_logic_vector(51, 8),
17855 => conv_std_logic_vector(51, 8),
17856 => conv_std_logic_vector(51, 8),
17857 => conv_std_logic_vector(52, 8),
17858 => conv_std_logic_vector(52, 8),
17859 => conv_std_logic_vector(52, 8),
17860 => conv_std_logic_vector(52, 8),
17861 => conv_std_logic_vector(53, 8),
17862 => conv_std_logic_vector(53, 8),
17863 => conv_std_logic_vector(53, 8),
17864 => conv_std_logic_vector(53, 8),
17865 => conv_std_logic_vector(54, 8),
17866 => conv_std_logic_vector(54, 8),
17867 => conv_std_logic_vector(54, 8),
17868 => conv_std_logic_vector(54, 8),
17869 => conv_std_logic_vector(55, 8),
17870 => conv_std_logic_vector(55, 8),
17871 => conv_std_logic_vector(55, 8),
17872 => conv_std_logic_vector(56, 8),
17873 => conv_std_logic_vector(56, 8),
17874 => conv_std_logic_vector(56, 8),
17875 => conv_std_logic_vector(56, 8),
17876 => conv_std_logic_vector(57, 8),
17877 => conv_std_logic_vector(57, 8),
17878 => conv_std_logic_vector(57, 8),
17879 => conv_std_logic_vector(57, 8),
17880 => conv_std_logic_vector(58, 8),
17881 => conv_std_logic_vector(58, 8),
17882 => conv_std_logic_vector(58, 8),
17883 => conv_std_logic_vector(59, 8),
17884 => conv_std_logic_vector(59, 8),
17885 => conv_std_logic_vector(59, 8),
17886 => conv_std_logic_vector(59, 8),
17887 => conv_std_logic_vector(60, 8),
17888 => conv_std_logic_vector(60, 8),
17889 => conv_std_logic_vector(60, 8),
17890 => conv_std_logic_vector(60, 8),
17891 => conv_std_logic_vector(61, 8),
17892 => conv_std_logic_vector(61, 8),
17893 => conv_std_logic_vector(61, 8),
17894 => conv_std_logic_vector(61, 8),
17895 => conv_std_logic_vector(62, 8),
17896 => conv_std_logic_vector(62, 8),
17897 => conv_std_logic_vector(62, 8),
17898 => conv_std_logic_vector(63, 8),
17899 => conv_std_logic_vector(63, 8),
17900 => conv_std_logic_vector(63, 8),
17901 => conv_std_logic_vector(63, 8),
17902 => conv_std_logic_vector(64, 8),
17903 => conv_std_logic_vector(64, 8),
17904 => conv_std_logic_vector(64, 8),
17905 => conv_std_logic_vector(64, 8),
17906 => conv_std_logic_vector(65, 8),
17907 => conv_std_logic_vector(65, 8),
17908 => conv_std_logic_vector(65, 8),
17909 => conv_std_logic_vector(66, 8),
17910 => conv_std_logic_vector(66, 8),
17911 => conv_std_logic_vector(66, 8),
17912 => conv_std_logic_vector(66, 8),
17913 => conv_std_logic_vector(67, 8),
17914 => conv_std_logic_vector(67, 8),
17915 => conv_std_logic_vector(67, 8),
17916 => conv_std_logic_vector(67, 8),
17917 => conv_std_logic_vector(68, 8),
17918 => conv_std_logic_vector(68, 8),
17919 => conv_std_logic_vector(68, 8),
17920 => conv_std_logic_vector(0, 8),
17921 => conv_std_logic_vector(0, 8),
17922 => conv_std_logic_vector(0, 8),
17923 => conv_std_logic_vector(0, 8),
17924 => conv_std_logic_vector(1, 8),
17925 => conv_std_logic_vector(1, 8),
17926 => conv_std_logic_vector(1, 8),
17927 => conv_std_logic_vector(1, 8),
17928 => conv_std_logic_vector(2, 8),
17929 => conv_std_logic_vector(2, 8),
17930 => conv_std_logic_vector(2, 8),
17931 => conv_std_logic_vector(3, 8),
17932 => conv_std_logic_vector(3, 8),
17933 => conv_std_logic_vector(3, 8),
17934 => conv_std_logic_vector(3, 8),
17935 => conv_std_logic_vector(4, 8),
17936 => conv_std_logic_vector(4, 8),
17937 => conv_std_logic_vector(4, 8),
17938 => conv_std_logic_vector(4, 8),
17939 => conv_std_logic_vector(5, 8),
17940 => conv_std_logic_vector(5, 8),
17941 => conv_std_logic_vector(5, 8),
17942 => conv_std_logic_vector(6, 8),
17943 => conv_std_logic_vector(6, 8),
17944 => conv_std_logic_vector(6, 8),
17945 => conv_std_logic_vector(6, 8),
17946 => conv_std_logic_vector(7, 8),
17947 => conv_std_logic_vector(7, 8),
17948 => conv_std_logic_vector(7, 8),
17949 => conv_std_logic_vector(7, 8),
17950 => conv_std_logic_vector(8, 8),
17951 => conv_std_logic_vector(8, 8),
17952 => conv_std_logic_vector(8, 8),
17953 => conv_std_logic_vector(9, 8),
17954 => conv_std_logic_vector(9, 8),
17955 => conv_std_logic_vector(9, 8),
17956 => conv_std_logic_vector(9, 8),
17957 => conv_std_logic_vector(10, 8),
17958 => conv_std_logic_vector(10, 8),
17959 => conv_std_logic_vector(10, 8),
17960 => conv_std_logic_vector(10, 8),
17961 => conv_std_logic_vector(11, 8),
17962 => conv_std_logic_vector(11, 8),
17963 => conv_std_logic_vector(11, 8),
17964 => conv_std_logic_vector(12, 8),
17965 => conv_std_logic_vector(12, 8),
17966 => conv_std_logic_vector(12, 8),
17967 => conv_std_logic_vector(12, 8),
17968 => conv_std_logic_vector(13, 8),
17969 => conv_std_logic_vector(13, 8),
17970 => conv_std_logic_vector(13, 8),
17971 => conv_std_logic_vector(13, 8),
17972 => conv_std_logic_vector(14, 8),
17973 => conv_std_logic_vector(14, 8),
17974 => conv_std_logic_vector(14, 8),
17975 => conv_std_logic_vector(15, 8),
17976 => conv_std_logic_vector(15, 8),
17977 => conv_std_logic_vector(15, 8),
17978 => conv_std_logic_vector(15, 8),
17979 => conv_std_logic_vector(16, 8),
17980 => conv_std_logic_vector(16, 8),
17981 => conv_std_logic_vector(16, 8),
17982 => conv_std_logic_vector(16, 8),
17983 => conv_std_logic_vector(17, 8),
17984 => conv_std_logic_vector(17, 8),
17985 => conv_std_logic_vector(17, 8),
17986 => conv_std_logic_vector(18, 8),
17987 => conv_std_logic_vector(18, 8),
17988 => conv_std_logic_vector(18, 8),
17989 => conv_std_logic_vector(18, 8),
17990 => conv_std_logic_vector(19, 8),
17991 => conv_std_logic_vector(19, 8),
17992 => conv_std_logic_vector(19, 8),
17993 => conv_std_logic_vector(19, 8),
17994 => conv_std_logic_vector(20, 8),
17995 => conv_std_logic_vector(20, 8),
17996 => conv_std_logic_vector(20, 8),
17997 => conv_std_logic_vector(21, 8),
17998 => conv_std_logic_vector(21, 8),
17999 => conv_std_logic_vector(21, 8),
18000 => conv_std_logic_vector(21, 8),
18001 => conv_std_logic_vector(22, 8),
18002 => conv_std_logic_vector(22, 8),
18003 => conv_std_logic_vector(22, 8),
18004 => conv_std_logic_vector(22, 8),
18005 => conv_std_logic_vector(23, 8),
18006 => conv_std_logic_vector(23, 8),
18007 => conv_std_logic_vector(23, 8),
18008 => conv_std_logic_vector(24, 8),
18009 => conv_std_logic_vector(24, 8),
18010 => conv_std_logic_vector(24, 8),
18011 => conv_std_logic_vector(24, 8),
18012 => conv_std_logic_vector(25, 8),
18013 => conv_std_logic_vector(25, 8),
18014 => conv_std_logic_vector(25, 8),
18015 => conv_std_logic_vector(25, 8),
18016 => conv_std_logic_vector(26, 8),
18017 => conv_std_logic_vector(26, 8),
18018 => conv_std_logic_vector(26, 8),
18019 => conv_std_logic_vector(27, 8),
18020 => conv_std_logic_vector(27, 8),
18021 => conv_std_logic_vector(27, 8),
18022 => conv_std_logic_vector(27, 8),
18023 => conv_std_logic_vector(28, 8),
18024 => conv_std_logic_vector(28, 8),
18025 => conv_std_logic_vector(28, 8),
18026 => conv_std_logic_vector(28, 8),
18027 => conv_std_logic_vector(29, 8),
18028 => conv_std_logic_vector(29, 8),
18029 => conv_std_logic_vector(29, 8),
18030 => conv_std_logic_vector(30, 8),
18031 => conv_std_logic_vector(30, 8),
18032 => conv_std_logic_vector(30, 8),
18033 => conv_std_logic_vector(30, 8),
18034 => conv_std_logic_vector(31, 8),
18035 => conv_std_logic_vector(31, 8),
18036 => conv_std_logic_vector(31, 8),
18037 => conv_std_logic_vector(31, 8),
18038 => conv_std_logic_vector(32, 8),
18039 => conv_std_logic_vector(32, 8),
18040 => conv_std_logic_vector(32, 8),
18041 => conv_std_logic_vector(33, 8),
18042 => conv_std_logic_vector(33, 8),
18043 => conv_std_logic_vector(33, 8),
18044 => conv_std_logic_vector(33, 8),
18045 => conv_std_logic_vector(34, 8),
18046 => conv_std_logic_vector(34, 8),
18047 => conv_std_logic_vector(34, 8),
18048 => conv_std_logic_vector(35, 8),
18049 => conv_std_logic_vector(35, 8),
18050 => conv_std_logic_vector(35, 8),
18051 => conv_std_logic_vector(35, 8),
18052 => conv_std_logic_vector(36, 8),
18053 => conv_std_logic_vector(36, 8),
18054 => conv_std_logic_vector(36, 8),
18055 => conv_std_logic_vector(36, 8),
18056 => conv_std_logic_vector(37, 8),
18057 => conv_std_logic_vector(37, 8),
18058 => conv_std_logic_vector(37, 8),
18059 => conv_std_logic_vector(38, 8),
18060 => conv_std_logic_vector(38, 8),
18061 => conv_std_logic_vector(38, 8),
18062 => conv_std_logic_vector(38, 8),
18063 => conv_std_logic_vector(39, 8),
18064 => conv_std_logic_vector(39, 8),
18065 => conv_std_logic_vector(39, 8),
18066 => conv_std_logic_vector(39, 8),
18067 => conv_std_logic_vector(40, 8),
18068 => conv_std_logic_vector(40, 8),
18069 => conv_std_logic_vector(40, 8),
18070 => conv_std_logic_vector(41, 8),
18071 => conv_std_logic_vector(41, 8),
18072 => conv_std_logic_vector(41, 8),
18073 => conv_std_logic_vector(41, 8),
18074 => conv_std_logic_vector(42, 8),
18075 => conv_std_logic_vector(42, 8),
18076 => conv_std_logic_vector(42, 8),
18077 => conv_std_logic_vector(42, 8),
18078 => conv_std_logic_vector(43, 8),
18079 => conv_std_logic_vector(43, 8),
18080 => conv_std_logic_vector(43, 8),
18081 => conv_std_logic_vector(44, 8),
18082 => conv_std_logic_vector(44, 8),
18083 => conv_std_logic_vector(44, 8),
18084 => conv_std_logic_vector(44, 8),
18085 => conv_std_logic_vector(45, 8),
18086 => conv_std_logic_vector(45, 8),
18087 => conv_std_logic_vector(45, 8),
18088 => conv_std_logic_vector(45, 8),
18089 => conv_std_logic_vector(46, 8),
18090 => conv_std_logic_vector(46, 8),
18091 => conv_std_logic_vector(46, 8),
18092 => conv_std_logic_vector(47, 8),
18093 => conv_std_logic_vector(47, 8),
18094 => conv_std_logic_vector(47, 8),
18095 => conv_std_logic_vector(47, 8),
18096 => conv_std_logic_vector(48, 8),
18097 => conv_std_logic_vector(48, 8),
18098 => conv_std_logic_vector(48, 8),
18099 => conv_std_logic_vector(48, 8),
18100 => conv_std_logic_vector(49, 8),
18101 => conv_std_logic_vector(49, 8),
18102 => conv_std_logic_vector(49, 8),
18103 => conv_std_logic_vector(50, 8),
18104 => conv_std_logic_vector(50, 8),
18105 => conv_std_logic_vector(50, 8),
18106 => conv_std_logic_vector(50, 8),
18107 => conv_std_logic_vector(51, 8),
18108 => conv_std_logic_vector(51, 8),
18109 => conv_std_logic_vector(51, 8),
18110 => conv_std_logic_vector(51, 8),
18111 => conv_std_logic_vector(52, 8),
18112 => conv_std_logic_vector(52, 8),
18113 => conv_std_logic_vector(52, 8),
18114 => conv_std_logic_vector(53, 8),
18115 => conv_std_logic_vector(53, 8),
18116 => conv_std_logic_vector(53, 8),
18117 => conv_std_logic_vector(53, 8),
18118 => conv_std_logic_vector(54, 8),
18119 => conv_std_logic_vector(54, 8),
18120 => conv_std_logic_vector(54, 8),
18121 => conv_std_logic_vector(54, 8),
18122 => conv_std_logic_vector(55, 8),
18123 => conv_std_logic_vector(55, 8),
18124 => conv_std_logic_vector(55, 8),
18125 => conv_std_logic_vector(56, 8),
18126 => conv_std_logic_vector(56, 8),
18127 => conv_std_logic_vector(56, 8),
18128 => conv_std_logic_vector(56, 8),
18129 => conv_std_logic_vector(57, 8),
18130 => conv_std_logic_vector(57, 8),
18131 => conv_std_logic_vector(57, 8),
18132 => conv_std_logic_vector(57, 8),
18133 => conv_std_logic_vector(58, 8),
18134 => conv_std_logic_vector(58, 8),
18135 => conv_std_logic_vector(58, 8),
18136 => conv_std_logic_vector(59, 8),
18137 => conv_std_logic_vector(59, 8),
18138 => conv_std_logic_vector(59, 8),
18139 => conv_std_logic_vector(59, 8),
18140 => conv_std_logic_vector(60, 8),
18141 => conv_std_logic_vector(60, 8),
18142 => conv_std_logic_vector(60, 8),
18143 => conv_std_logic_vector(60, 8),
18144 => conv_std_logic_vector(61, 8),
18145 => conv_std_logic_vector(61, 8),
18146 => conv_std_logic_vector(61, 8),
18147 => conv_std_logic_vector(62, 8),
18148 => conv_std_logic_vector(62, 8),
18149 => conv_std_logic_vector(62, 8),
18150 => conv_std_logic_vector(62, 8),
18151 => conv_std_logic_vector(63, 8),
18152 => conv_std_logic_vector(63, 8),
18153 => conv_std_logic_vector(63, 8),
18154 => conv_std_logic_vector(63, 8),
18155 => conv_std_logic_vector(64, 8),
18156 => conv_std_logic_vector(64, 8),
18157 => conv_std_logic_vector(64, 8),
18158 => conv_std_logic_vector(65, 8),
18159 => conv_std_logic_vector(65, 8),
18160 => conv_std_logic_vector(65, 8),
18161 => conv_std_logic_vector(65, 8),
18162 => conv_std_logic_vector(66, 8),
18163 => conv_std_logic_vector(66, 8),
18164 => conv_std_logic_vector(66, 8),
18165 => conv_std_logic_vector(66, 8),
18166 => conv_std_logic_vector(67, 8),
18167 => conv_std_logic_vector(67, 8),
18168 => conv_std_logic_vector(67, 8),
18169 => conv_std_logic_vector(68, 8),
18170 => conv_std_logic_vector(68, 8),
18171 => conv_std_logic_vector(68, 8),
18172 => conv_std_logic_vector(68, 8),
18173 => conv_std_logic_vector(69, 8),
18174 => conv_std_logic_vector(69, 8),
18175 => conv_std_logic_vector(69, 8),
18176 => conv_std_logic_vector(0, 8),
18177 => conv_std_logic_vector(0, 8),
18178 => conv_std_logic_vector(0, 8),
18179 => conv_std_logic_vector(0, 8),
18180 => conv_std_logic_vector(1, 8),
18181 => conv_std_logic_vector(1, 8),
18182 => conv_std_logic_vector(1, 8),
18183 => conv_std_logic_vector(1, 8),
18184 => conv_std_logic_vector(2, 8),
18185 => conv_std_logic_vector(2, 8),
18186 => conv_std_logic_vector(2, 8),
18187 => conv_std_logic_vector(3, 8),
18188 => conv_std_logic_vector(3, 8),
18189 => conv_std_logic_vector(3, 8),
18190 => conv_std_logic_vector(3, 8),
18191 => conv_std_logic_vector(4, 8),
18192 => conv_std_logic_vector(4, 8),
18193 => conv_std_logic_vector(4, 8),
18194 => conv_std_logic_vector(4, 8),
18195 => conv_std_logic_vector(5, 8),
18196 => conv_std_logic_vector(5, 8),
18197 => conv_std_logic_vector(5, 8),
18198 => conv_std_logic_vector(6, 8),
18199 => conv_std_logic_vector(6, 8),
18200 => conv_std_logic_vector(6, 8),
18201 => conv_std_logic_vector(6, 8),
18202 => conv_std_logic_vector(7, 8),
18203 => conv_std_logic_vector(7, 8),
18204 => conv_std_logic_vector(7, 8),
18205 => conv_std_logic_vector(8, 8),
18206 => conv_std_logic_vector(8, 8),
18207 => conv_std_logic_vector(8, 8),
18208 => conv_std_logic_vector(8, 8),
18209 => conv_std_logic_vector(9, 8),
18210 => conv_std_logic_vector(9, 8),
18211 => conv_std_logic_vector(9, 8),
18212 => conv_std_logic_vector(9, 8),
18213 => conv_std_logic_vector(10, 8),
18214 => conv_std_logic_vector(10, 8),
18215 => conv_std_logic_vector(10, 8),
18216 => conv_std_logic_vector(11, 8),
18217 => conv_std_logic_vector(11, 8),
18218 => conv_std_logic_vector(11, 8),
18219 => conv_std_logic_vector(11, 8),
18220 => conv_std_logic_vector(12, 8),
18221 => conv_std_logic_vector(12, 8),
18222 => conv_std_logic_vector(12, 8),
18223 => conv_std_logic_vector(13, 8),
18224 => conv_std_logic_vector(13, 8),
18225 => conv_std_logic_vector(13, 8),
18226 => conv_std_logic_vector(13, 8),
18227 => conv_std_logic_vector(14, 8),
18228 => conv_std_logic_vector(14, 8),
18229 => conv_std_logic_vector(14, 8),
18230 => conv_std_logic_vector(14, 8),
18231 => conv_std_logic_vector(15, 8),
18232 => conv_std_logic_vector(15, 8),
18233 => conv_std_logic_vector(15, 8),
18234 => conv_std_logic_vector(16, 8),
18235 => conv_std_logic_vector(16, 8),
18236 => conv_std_logic_vector(16, 8),
18237 => conv_std_logic_vector(16, 8),
18238 => conv_std_logic_vector(17, 8),
18239 => conv_std_logic_vector(17, 8),
18240 => conv_std_logic_vector(17, 8),
18241 => conv_std_logic_vector(18, 8),
18242 => conv_std_logic_vector(18, 8),
18243 => conv_std_logic_vector(18, 8),
18244 => conv_std_logic_vector(18, 8),
18245 => conv_std_logic_vector(19, 8),
18246 => conv_std_logic_vector(19, 8),
18247 => conv_std_logic_vector(19, 8),
18248 => conv_std_logic_vector(19, 8),
18249 => conv_std_logic_vector(20, 8),
18250 => conv_std_logic_vector(20, 8),
18251 => conv_std_logic_vector(20, 8),
18252 => conv_std_logic_vector(21, 8),
18253 => conv_std_logic_vector(21, 8),
18254 => conv_std_logic_vector(21, 8),
18255 => conv_std_logic_vector(21, 8),
18256 => conv_std_logic_vector(22, 8),
18257 => conv_std_logic_vector(22, 8),
18258 => conv_std_logic_vector(22, 8),
18259 => conv_std_logic_vector(23, 8),
18260 => conv_std_logic_vector(23, 8),
18261 => conv_std_logic_vector(23, 8),
18262 => conv_std_logic_vector(23, 8),
18263 => conv_std_logic_vector(24, 8),
18264 => conv_std_logic_vector(24, 8),
18265 => conv_std_logic_vector(24, 8),
18266 => conv_std_logic_vector(24, 8),
18267 => conv_std_logic_vector(25, 8),
18268 => conv_std_logic_vector(25, 8),
18269 => conv_std_logic_vector(25, 8),
18270 => conv_std_logic_vector(26, 8),
18271 => conv_std_logic_vector(26, 8),
18272 => conv_std_logic_vector(26, 8),
18273 => conv_std_logic_vector(26, 8),
18274 => conv_std_logic_vector(27, 8),
18275 => conv_std_logic_vector(27, 8),
18276 => conv_std_logic_vector(27, 8),
18277 => conv_std_logic_vector(28, 8),
18278 => conv_std_logic_vector(28, 8),
18279 => conv_std_logic_vector(28, 8),
18280 => conv_std_logic_vector(28, 8),
18281 => conv_std_logic_vector(29, 8),
18282 => conv_std_logic_vector(29, 8),
18283 => conv_std_logic_vector(29, 8),
18284 => conv_std_logic_vector(29, 8),
18285 => conv_std_logic_vector(30, 8),
18286 => conv_std_logic_vector(30, 8),
18287 => conv_std_logic_vector(30, 8),
18288 => conv_std_logic_vector(31, 8),
18289 => conv_std_logic_vector(31, 8),
18290 => conv_std_logic_vector(31, 8),
18291 => conv_std_logic_vector(31, 8),
18292 => conv_std_logic_vector(32, 8),
18293 => conv_std_logic_vector(32, 8),
18294 => conv_std_logic_vector(32, 8),
18295 => conv_std_logic_vector(33, 8),
18296 => conv_std_logic_vector(33, 8),
18297 => conv_std_logic_vector(33, 8),
18298 => conv_std_logic_vector(33, 8),
18299 => conv_std_logic_vector(34, 8),
18300 => conv_std_logic_vector(34, 8),
18301 => conv_std_logic_vector(34, 8),
18302 => conv_std_logic_vector(34, 8),
18303 => conv_std_logic_vector(35, 8),
18304 => conv_std_logic_vector(35, 8),
18305 => conv_std_logic_vector(35, 8),
18306 => conv_std_logic_vector(36, 8),
18307 => conv_std_logic_vector(36, 8),
18308 => conv_std_logic_vector(36, 8),
18309 => conv_std_logic_vector(36, 8),
18310 => conv_std_logic_vector(37, 8),
18311 => conv_std_logic_vector(37, 8),
18312 => conv_std_logic_vector(37, 8),
18313 => conv_std_logic_vector(37, 8),
18314 => conv_std_logic_vector(38, 8),
18315 => conv_std_logic_vector(38, 8),
18316 => conv_std_logic_vector(38, 8),
18317 => conv_std_logic_vector(39, 8),
18318 => conv_std_logic_vector(39, 8),
18319 => conv_std_logic_vector(39, 8),
18320 => conv_std_logic_vector(39, 8),
18321 => conv_std_logic_vector(40, 8),
18322 => conv_std_logic_vector(40, 8),
18323 => conv_std_logic_vector(40, 8),
18324 => conv_std_logic_vector(41, 8),
18325 => conv_std_logic_vector(41, 8),
18326 => conv_std_logic_vector(41, 8),
18327 => conv_std_logic_vector(41, 8),
18328 => conv_std_logic_vector(42, 8),
18329 => conv_std_logic_vector(42, 8),
18330 => conv_std_logic_vector(42, 8),
18331 => conv_std_logic_vector(42, 8),
18332 => conv_std_logic_vector(43, 8),
18333 => conv_std_logic_vector(43, 8),
18334 => conv_std_logic_vector(43, 8),
18335 => conv_std_logic_vector(44, 8),
18336 => conv_std_logic_vector(44, 8),
18337 => conv_std_logic_vector(44, 8),
18338 => conv_std_logic_vector(44, 8),
18339 => conv_std_logic_vector(45, 8),
18340 => conv_std_logic_vector(45, 8),
18341 => conv_std_logic_vector(45, 8),
18342 => conv_std_logic_vector(46, 8),
18343 => conv_std_logic_vector(46, 8),
18344 => conv_std_logic_vector(46, 8),
18345 => conv_std_logic_vector(46, 8),
18346 => conv_std_logic_vector(47, 8),
18347 => conv_std_logic_vector(47, 8),
18348 => conv_std_logic_vector(47, 8),
18349 => conv_std_logic_vector(47, 8),
18350 => conv_std_logic_vector(48, 8),
18351 => conv_std_logic_vector(48, 8),
18352 => conv_std_logic_vector(48, 8),
18353 => conv_std_logic_vector(49, 8),
18354 => conv_std_logic_vector(49, 8),
18355 => conv_std_logic_vector(49, 8),
18356 => conv_std_logic_vector(49, 8),
18357 => conv_std_logic_vector(50, 8),
18358 => conv_std_logic_vector(50, 8),
18359 => conv_std_logic_vector(50, 8),
18360 => conv_std_logic_vector(51, 8),
18361 => conv_std_logic_vector(51, 8),
18362 => conv_std_logic_vector(51, 8),
18363 => conv_std_logic_vector(51, 8),
18364 => conv_std_logic_vector(52, 8),
18365 => conv_std_logic_vector(52, 8),
18366 => conv_std_logic_vector(52, 8),
18367 => conv_std_logic_vector(52, 8),
18368 => conv_std_logic_vector(53, 8),
18369 => conv_std_logic_vector(53, 8),
18370 => conv_std_logic_vector(53, 8),
18371 => conv_std_logic_vector(54, 8),
18372 => conv_std_logic_vector(54, 8),
18373 => conv_std_logic_vector(54, 8),
18374 => conv_std_logic_vector(54, 8),
18375 => conv_std_logic_vector(55, 8),
18376 => conv_std_logic_vector(55, 8),
18377 => conv_std_logic_vector(55, 8),
18378 => conv_std_logic_vector(56, 8),
18379 => conv_std_logic_vector(56, 8),
18380 => conv_std_logic_vector(56, 8),
18381 => conv_std_logic_vector(56, 8),
18382 => conv_std_logic_vector(57, 8),
18383 => conv_std_logic_vector(57, 8),
18384 => conv_std_logic_vector(57, 8),
18385 => conv_std_logic_vector(57, 8),
18386 => conv_std_logic_vector(58, 8),
18387 => conv_std_logic_vector(58, 8),
18388 => conv_std_logic_vector(58, 8),
18389 => conv_std_logic_vector(59, 8),
18390 => conv_std_logic_vector(59, 8),
18391 => conv_std_logic_vector(59, 8),
18392 => conv_std_logic_vector(59, 8),
18393 => conv_std_logic_vector(60, 8),
18394 => conv_std_logic_vector(60, 8),
18395 => conv_std_logic_vector(60, 8),
18396 => conv_std_logic_vector(61, 8),
18397 => conv_std_logic_vector(61, 8),
18398 => conv_std_logic_vector(61, 8),
18399 => conv_std_logic_vector(61, 8),
18400 => conv_std_logic_vector(62, 8),
18401 => conv_std_logic_vector(62, 8),
18402 => conv_std_logic_vector(62, 8),
18403 => conv_std_logic_vector(62, 8),
18404 => conv_std_logic_vector(63, 8),
18405 => conv_std_logic_vector(63, 8),
18406 => conv_std_logic_vector(63, 8),
18407 => conv_std_logic_vector(64, 8),
18408 => conv_std_logic_vector(64, 8),
18409 => conv_std_logic_vector(64, 8),
18410 => conv_std_logic_vector(64, 8),
18411 => conv_std_logic_vector(65, 8),
18412 => conv_std_logic_vector(65, 8),
18413 => conv_std_logic_vector(65, 8),
18414 => conv_std_logic_vector(66, 8),
18415 => conv_std_logic_vector(66, 8),
18416 => conv_std_logic_vector(66, 8),
18417 => conv_std_logic_vector(66, 8),
18418 => conv_std_logic_vector(67, 8),
18419 => conv_std_logic_vector(67, 8),
18420 => conv_std_logic_vector(67, 8),
18421 => conv_std_logic_vector(67, 8),
18422 => conv_std_logic_vector(68, 8),
18423 => conv_std_logic_vector(68, 8),
18424 => conv_std_logic_vector(68, 8),
18425 => conv_std_logic_vector(69, 8),
18426 => conv_std_logic_vector(69, 8),
18427 => conv_std_logic_vector(69, 8),
18428 => conv_std_logic_vector(69, 8),
18429 => conv_std_logic_vector(70, 8),
18430 => conv_std_logic_vector(70, 8),
18431 => conv_std_logic_vector(70, 8),
18432 => conv_std_logic_vector(0, 8),
18433 => conv_std_logic_vector(0, 8),
18434 => conv_std_logic_vector(0, 8),
18435 => conv_std_logic_vector(0, 8),
18436 => conv_std_logic_vector(1, 8),
18437 => conv_std_logic_vector(1, 8),
18438 => conv_std_logic_vector(1, 8),
18439 => conv_std_logic_vector(1, 8),
18440 => conv_std_logic_vector(2, 8),
18441 => conv_std_logic_vector(2, 8),
18442 => conv_std_logic_vector(2, 8),
18443 => conv_std_logic_vector(3, 8),
18444 => conv_std_logic_vector(3, 8),
18445 => conv_std_logic_vector(3, 8),
18446 => conv_std_logic_vector(3, 8),
18447 => conv_std_logic_vector(4, 8),
18448 => conv_std_logic_vector(4, 8),
18449 => conv_std_logic_vector(4, 8),
18450 => conv_std_logic_vector(5, 8),
18451 => conv_std_logic_vector(5, 8),
18452 => conv_std_logic_vector(5, 8),
18453 => conv_std_logic_vector(5, 8),
18454 => conv_std_logic_vector(6, 8),
18455 => conv_std_logic_vector(6, 8),
18456 => conv_std_logic_vector(6, 8),
18457 => conv_std_logic_vector(7, 8),
18458 => conv_std_logic_vector(7, 8),
18459 => conv_std_logic_vector(7, 8),
18460 => conv_std_logic_vector(7, 8),
18461 => conv_std_logic_vector(8, 8),
18462 => conv_std_logic_vector(8, 8),
18463 => conv_std_logic_vector(8, 8),
18464 => conv_std_logic_vector(9, 8),
18465 => conv_std_logic_vector(9, 8),
18466 => conv_std_logic_vector(9, 8),
18467 => conv_std_logic_vector(9, 8),
18468 => conv_std_logic_vector(10, 8),
18469 => conv_std_logic_vector(10, 8),
18470 => conv_std_logic_vector(10, 8),
18471 => conv_std_logic_vector(10, 8),
18472 => conv_std_logic_vector(11, 8),
18473 => conv_std_logic_vector(11, 8),
18474 => conv_std_logic_vector(11, 8),
18475 => conv_std_logic_vector(12, 8),
18476 => conv_std_logic_vector(12, 8),
18477 => conv_std_logic_vector(12, 8),
18478 => conv_std_logic_vector(12, 8),
18479 => conv_std_logic_vector(13, 8),
18480 => conv_std_logic_vector(13, 8),
18481 => conv_std_logic_vector(13, 8),
18482 => conv_std_logic_vector(14, 8),
18483 => conv_std_logic_vector(14, 8),
18484 => conv_std_logic_vector(14, 8),
18485 => conv_std_logic_vector(14, 8),
18486 => conv_std_logic_vector(15, 8),
18487 => conv_std_logic_vector(15, 8),
18488 => conv_std_logic_vector(15, 8),
18489 => conv_std_logic_vector(16, 8),
18490 => conv_std_logic_vector(16, 8),
18491 => conv_std_logic_vector(16, 8),
18492 => conv_std_logic_vector(16, 8),
18493 => conv_std_logic_vector(17, 8),
18494 => conv_std_logic_vector(17, 8),
18495 => conv_std_logic_vector(17, 8),
18496 => conv_std_logic_vector(18, 8),
18497 => conv_std_logic_vector(18, 8),
18498 => conv_std_logic_vector(18, 8),
18499 => conv_std_logic_vector(18, 8),
18500 => conv_std_logic_vector(19, 8),
18501 => conv_std_logic_vector(19, 8),
18502 => conv_std_logic_vector(19, 8),
18503 => conv_std_logic_vector(19, 8),
18504 => conv_std_logic_vector(20, 8),
18505 => conv_std_logic_vector(20, 8),
18506 => conv_std_logic_vector(20, 8),
18507 => conv_std_logic_vector(21, 8),
18508 => conv_std_logic_vector(21, 8),
18509 => conv_std_logic_vector(21, 8),
18510 => conv_std_logic_vector(21, 8),
18511 => conv_std_logic_vector(22, 8),
18512 => conv_std_logic_vector(22, 8),
18513 => conv_std_logic_vector(22, 8),
18514 => conv_std_logic_vector(23, 8),
18515 => conv_std_logic_vector(23, 8),
18516 => conv_std_logic_vector(23, 8),
18517 => conv_std_logic_vector(23, 8),
18518 => conv_std_logic_vector(24, 8),
18519 => conv_std_logic_vector(24, 8),
18520 => conv_std_logic_vector(24, 8),
18521 => conv_std_logic_vector(25, 8),
18522 => conv_std_logic_vector(25, 8),
18523 => conv_std_logic_vector(25, 8),
18524 => conv_std_logic_vector(25, 8),
18525 => conv_std_logic_vector(26, 8),
18526 => conv_std_logic_vector(26, 8),
18527 => conv_std_logic_vector(26, 8),
18528 => conv_std_logic_vector(27, 8),
18529 => conv_std_logic_vector(27, 8),
18530 => conv_std_logic_vector(27, 8),
18531 => conv_std_logic_vector(27, 8),
18532 => conv_std_logic_vector(28, 8),
18533 => conv_std_logic_vector(28, 8),
18534 => conv_std_logic_vector(28, 8),
18535 => conv_std_logic_vector(28, 8),
18536 => conv_std_logic_vector(29, 8),
18537 => conv_std_logic_vector(29, 8),
18538 => conv_std_logic_vector(29, 8),
18539 => conv_std_logic_vector(30, 8),
18540 => conv_std_logic_vector(30, 8),
18541 => conv_std_logic_vector(30, 8),
18542 => conv_std_logic_vector(30, 8),
18543 => conv_std_logic_vector(31, 8),
18544 => conv_std_logic_vector(31, 8),
18545 => conv_std_logic_vector(31, 8),
18546 => conv_std_logic_vector(32, 8),
18547 => conv_std_logic_vector(32, 8),
18548 => conv_std_logic_vector(32, 8),
18549 => conv_std_logic_vector(32, 8),
18550 => conv_std_logic_vector(33, 8),
18551 => conv_std_logic_vector(33, 8),
18552 => conv_std_logic_vector(33, 8),
18553 => conv_std_logic_vector(34, 8),
18554 => conv_std_logic_vector(34, 8),
18555 => conv_std_logic_vector(34, 8),
18556 => conv_std_logic_vector(34, 8),
18557 => conv_std_logic_vector(35, 8),
18558 => conv_std_logic_vector(35, 8),
18559 => conv_std_logic_vector(35, 8),
18560 => conv_std_logic_vector(36, 8),
18561 => conv_std_logic_vector(36, 8),
18562 => conv_std_logic_vector(36, 8),
18563 => conv_std_logic_vector(36, 8),
18564 => conv_std_logic_vector(37, 8),
18565 => conv_std_logic_vector(37, 8),
18566 => conv_std_logic_vector(37, 8),
18567 => conv_std_logic_vector(37, 8),
18568 => conv_std_logic_vector(38, 8),
18569 => conv_std_logic_vector(38, 8),
18570 => conv_std_logic_vector(38, 8),
18571 => conv_std_logic_vector(39, 8),
18572 => conv_std_logic_vector(39, 8),
18573 => conv_std_logic_vector(39, 8),
18574 => conv_std_logic_vector(39, 8),
18575 => conv_std_logic_vector(40, 8),
18576 => conv_std_logic_vector(40, 8),
18577 => conv_std_logic_vector(40, 8),
18578 => conv_std_logic_vector(41, 8),
18579 => conv_std_logic_vector(41, 8),
18580 => conv_std_logic_vector(41, 8),
18581 => conv_std_logic_vector(41, 8),
18582 => conv_std_logic_vector(42, 8),
18583 => conv_std_logic_vector(42, 8),
18584 => conv_std_logic_vector(42, 8),
18585 => conv_std_logic_vector(43, 8),
18586 => conv_std_logic_vector(43, 8),
18587 => conv_std_logic_vector(43, 8),
18588 => conv_std_logic_vector(43, 8),
18589 => conv_std_logic_vector(44, 8),
18590 => conv_std_logic_vector(44, 8),
18591 => conv_std_logic_vector(44, 8),
18592 => conv_std_logic_vector(45, 8),
18593 => conv_std_logic_vector(45, 8),
18594 => conv_std_logic_vector(45, 8),
18595 => conv_std_logic_vector(45, 8),
18596 => conv_std_logic_vector(46, 8),
18597 => conv_std_logic_vector(46, 8),
18598 => conv_std_logic_vector(46, 8),
18599 => conv_std_logic_vector(46, 8),
18600 => conv_std_logic_vector(47, 8),
18601 => conv_std_logic_vector(47, 8),
18602 => conv_std_logic_vector(47, 8),
18603 => conv_std_logic_vector(48, 8),
18604 => conv_std_logic_vector(48, 8),
18605 => conv_std_logic_vector(48, 8),
18606 => conv_std_logic_vector(48, 8),
18607 => conv_std_logic_vector(49, 8),
18608 => conv_std_logic_vector(49, 8),
18609 => conv_std_logic_vector(49, 8),
18610 => conv_std_logic_vector(50, 8),
18611 => conv_std_logic_vector(50, 8),
18612 => conv_std_logic_vector(50, 8),
18613 => conv_std_logic_vector(50, 8),
18614 => conv_std_logic_vector(51, 8),
18615 => conv_std_logic_vector(51, 8),
18616 => conv_std_logic_vector(51, 8),
18617 => conv_std_logic_vector(52, 8),
18618 => conv_std_logic_vector(52, 8),
18619 => conv_std_logic_vector(52, 8),
18620 => conv_std_logic_vector(52, 8),
18621 => conv_std_logic_vector(53, 8),
18622 => conv_std_logic_vector(53, 8),
18623 => conv_std_logic_vector(53, 8),
18624 => conv_std_logic_vector(54, 8),
18625 => conv_std_logic_vector(54, 8),
18626 => conv_std_logic_vector(54, 8),
18627 => conv_std_logic_vector(54, 8),
18628 => conv_std_logic_vector(55, 8),
18629 => conv_std_logic_vector(55, 8),
18630 => conv_std_logic_vector(55, 8),
18631 => conv_std_logic_vector(55, 8),
18632 => conv_std_logic_vector(56, 8),
18633 => conv_std_logic_vector(56, 8),
18634 => conv_std_logic_vector(56, 8),
18635 => conv_std_logic_vector(57, 8),
18636 => conv_std_logic_vector(57, 8),
18637 => conv_std_logic_vector(57, 8),
18638 => conv_std_logic_vector(57, 8),
18639 => conv_std_logic_vector(58, 8),
18640 => conv_std_logic_vector(58, 8),
18641 => conv_std_logic_vector(58, 8),
18642 => conv_std_logic_vector(59, 8),
18643 => conv_std_logic_vector(59, 8),
18644 => conv_std_logic_vector(59, 8),
18645 => conv_std_logic_vector(59, 8),
18646 => conv_std_logic_vector(60, 8),
18647 => conv_std_logic_vector(60, 8),
18648 => conv_std_logic_vector(60, 8),
18649 => conv_std_logic_vector(61, 8),
18650 => conv_std_logic_vector(61, 8),
18651 => conv_std_logic_vector(61, 8),
18652 => conv_std_logic_vector(61, 8),
18653 => conv_std_logic_vector(62, 8),
18654 => conv_std_logic_vector(62, 8),
18655 => conv_std_logic_vector(62, 8),
18656 => conv_std_logic_vector(63, 8),
18657 => conv_std_logic_vector(63, 8),
18658 => conv_std_logic_vector(63, 8),
18659 => conv_std_logic_vector(63, 8),
18660 => conv_std_logic_vector(64, 8),
18661 => conv_std_logic_vector(64, 8),
18662 => conv_std_logic_vector(64, 8),
18663 => conv_std_logic_vector(64, 8),
18664 => conv_std_logic_vector(65, 8),
18665 => conv_std_logic_vector(65, 8),
18666 => conv_std_logic_vector(65, 8),
18667 => conv_std_logic_vector(66, 8),
18668 => conv_std_logic_vector(66, 8),
18669 => conv_std_logic_vector(66, 8),
18670 => conv_std_logic_vector(66, 8),
18671 => conv_std_logic_vector(67, 8),
18672 => conv_std_logic_vector(67, 8),
18673 => conv_std_logic_vector(67, 8),
18674 => conv_std_logic_vector(68, 8),
18675 => conv_std_logic_vector(68, 8),
18676 => conv_std_logic_vector(68, 8),
18677 => conv_std_logic_vector(68, 8),
18678 => conv_std_logic_vector(69, 8),
18679 => conv_std_logic_vector(69, 8),
18680 => conv_std_logic_vector(69, 8),
18681 => conv_std_logic_vector(70, 8),
18682 => conv_std_logic_vector(70, 8),
18683 => conv_std_logic_vector(70, 8),
18684 => conv_std_logic_vector(70, 8),
18685 => conv_std_logic_vector(71, 8),
18686 => conv_std_logic_vector(71, 8),
18687 => conv_std_logic_vector(71, 8),
18688 => conv_std_logic_vector(0, 8),
18689 => conv_std_logic_vector(0, 8),
18690 => conv_std_logic_vector(0, 8),
18691 => conv_std_logic_vector(0, 8),
18692 => conv_std_logic_vector(1, 8),
18693 => conv_std_logic_vector(1, 8),
18694 => conv_std_logic_vector(1, 8),
18695 => conv_std_logic_vector(1, 8),
18696 => conv_std_logic_vector(2, 8),
18697 => conv_std_logic_vector(2, 8),
18698 => conv_std_logic_vector(2, 8),
18699 => conv_std_logic_vector(3, 8),
18700 => conv_std_logic_vector(3, 8),
18701 => conv_std_logic_vector(3, 8),
18702 => conv_std_logic_vector(3, 8),
18703 => conv_std_logic_vector(4, 8),
18704 => conv_std_logic_vector(4, 8),
18705 => conv_std_logic_vector(4, 8),
18706 => conv_std_logic_vector(5, 8),
18707 => conv_std_logic_vector(5, 8),
18708 => conv_std_logic_vector(5, 8),
18709 => conv_std_logic_vector(5, 8),
18710 => conv_std_logic_vector(6, 8),
18711 => conv_std_logic_vector(6, 8),
18712 => conv_std_logic_vector(6, 8),
18713 => conv_std_logic_vector(7, 8),
18714 => conv_std_logic_vector(7, 8),
18715 => conv_std_logic_vector(7, 8),
18716 => conv_std_logic_vector(7, 8),
18717 => conv_std_logic_vector(8, 8),
18718 => conv_std_logic_vector(8, 8),
18719 => conv_std_logic_vector(8, 8),
18720 => conv_std_logic_vector(9, 8),
18721 => conv_std_logic_vector(9, 8),
18722 => conv_std_logic_vector(9, 8),
18723 => conv_std_logic_vector(9, 8),
18724 => conv_std_logic_vector(10, 8),
18725 => conv_std_logic_vector(10, 8),
18726 => conv_std_logic_vector(10, 8),
18727 => conv_std_logic_vector(11, 8),
18728 => conv_std_logic_vector(11, 8),
18729 => conv_std_logic_vector(11, 8),
18730 => conv_std_logic_vector(11, 8),
18731 => conv_std_logic_vector(12, 8),
18732 => conv_std_logic_vector(12, 8),
18733 => conv_std_logic_vector(12, 8),
18734 => conv_std_logic_vector(13, 8),
18735 => conv_std_logic_vector(13, 8),
18736 => conv_std_logic_vector(13, 8),
18737 => conv_std_logic_vector(13, 8),
18738 => conv_std_logic_vector(14, 8),
18739 => conv_std_logic_vector(14, 8),
18740 => conv_std_logic_vector(14, 8),
18741 => conv_std_logic_vector(15, 8),
18742 => conv_std_logic_vector(15, 8),
18743 => conv_std_logic_vector(15, 8),
18744 => conv_std_logic_vector(15, 8),
18745 => conv_std_logic_vector(16, 8),
18746 => conv_std_logic_vector(16, 8),
18747 => conv_std_logic_vector(16, 8),
18748 => conv_std_logic_vector(17, 8),
18749 => conv_std_logic_vector(17, 8),
18750 => conv_std_logic_vector(17, 8),
18751 => conv_std_logic_vector(17, 8),
18752 => conv_std_logic_vector(18, 8),
18753 => conv_std_logic_vector(18, 8),
18754 => conv_std_logic_vector(18, 8),
18755 => conv_std_logic_vector(19, 8),
18756 => conv_std_logic_vector(19, 8),
18757 => conv_std_logic_vector(19, 8),
18758 => conv_std_logic_vector(19, 8),
18759 => conv_std_logic_vector(20, 8),
18760 => conv_std_logic_vector(20, 8),
18761 => conv_std_logic_vector(20, 8),
18762 => conv_std_logic_vector(21, 8),
18763 => conv_std_logic_vector(21, 8),
18764 => conv_std_logic_vector(21, 8),
18765 => conv_std_logic_vector(21, 8),
18766 => conv_std_logic_vector(22, 8),
18767 => conv_std_logic_vector(22, 8),
18768 => conv_std_logic_vector(22, 8),
18769 => conv_std_logic_vector(23, 8),
18770 => conv_std_logic_vector(23, 8),
18771 => conv_std_logic_vector(23, 8),
18772 => conv_std_logic_vector(23, 8),
18773 => conv_std_logic_vector(24, 8),
18774 => conv_std_logic_vector(24, 8),
18775 => conv_std_logic_vector(24, 8),
18776 => conv_std_logic_vector(25, 8),
18777 => conv_std_logic_vector(25, 8),
18778 => conv_std_logic_vector(25, 8),
18779 => conv_std_logic_vector(25, 8),
18780 => conv_std_logic_vector(26, 8),
18781 => conv_std_logic_vector(26, 8),
18782 => conv_std_logic_vector(26, 8),
18783 => conv_std_logic_vector(27, 8),
18784 => conv_std_logic_vector(27, 8),
18785 => conv_std_logic_vector(27, 8),
18786 => conv_std_logic_vector(27, 8),
18787 => conv_std_logic_vector(28, 8),
18788 => conv_std_logic_vector(28, 8),
18789 => conv_std_logic_vector(28, 8),
18790 => conv_std_logic_vector(29, 8),
18791 => conv_std_logic_vector(29, 8),
18792 => conv_std_logic_vector(29, 8),
18793 => conv_std_logic_vector(29, 8),
18794 => conv_std_logic_vector(30, 8),
18795 => conv_std_logic_vector(30, 8),
18796 => conv_std_logic_vector(30, 8),
18797 => conv_std_logic_vector(31, 8),
18798 => conv_std_logic_vector(31, 8),
18799 => conv_std_logic_vector(31, 8),
18800 => conv_std_logic_vector(31, 8),
18801 => conv_std_logic_vector(32, 8),
18802 => conv_std_logic_vector(32, 8),
18803 => conv_std_logic_vector(32, 8),
18804 => conv_std_logic_vector(33, 8),
18805 => conv_std_logic_vector(33, 8),
18806 => conv_std_logic_vector(33, 8),
18807 => conv_std_logic_vector(33, 8),
18808 => conv_std_logic_vector(34, 8),
18809 => conv_std_logic_vector(34, 8),
18810 => conv_std_logic_vector(34, 8),
18811 => conv_std_logic_vector(35, 8),
18812 => conv_std_logic_vector(35, 8),
18813 => conv_std_logic_vector(35, 8),
18814 => conv_std_logic_vector(35, 8),
18815 => conv_std_logic_vector(36, 8),
18816 => conv_std_logic_vector(36, 8),
18817 => conv_std_logic_vector(36, 8),
18818 => conv_std_logic_vector(37, 8),
18819 => conv_std_logic_vector(37, 8),
18820 => conv_std_logic_vector(37, 8),
18821 => conv_std_logic_vector(37, 8),
18822 => conv_std_logic_vector(38, 8),
18823 => conv_std_logic_vector(38, 8),
18824 => conv_std_logic_vector(38, 8),
18825 => conv_std_logic_vector(39, 8),
18826 => conv_std_logic_vector(39, 8),
18827 => conv_std_logic_vector(39, 8),
18828 => conv_std_logic_vector(39, 8),
18829 => conv_std_logic_vector(40, 8),
18830 => conv_std_logic_vector(40, 8),
18831 => conv_std_logic_vector(40, 8),
18832 => conv_std_logic_vector(41, 8),
18833 => conv_std_logic_vector(41, 8),
18834 => conv_std_logic_vector(41, 8),
18835 => conv_std_logic_vector(41, 8),
18836 => conv_std_logic_vector(42, 8),
18837 => conv_std_logic_vector(42, 8),
18838 => conv_std_logic_vector(42, 8),
18839 => conv_std_logic_vector(43, 8),
18840 => conv_std_logic_vector(43, 8),
18841 => conv_std_logic_vector(43, 8),
18842 => conv_std_logic_vector(43, 8),
18843 => conv_std_logic_vector(44, 8),
18844 => conv_std_logic_vector(44, 8),
18845 => conv_std_logic_vector(44, 8),
18846 => conv_std_logic_vector(45, 8),
18847 => conv_std_logic_vector(45, 8),
18848 => conv_std_logic_vector(45, 8),
18849 => conv_std_logic_vector(45, 8),
18850 => conv_std_logic_vector(46, 8),
18851 => conv_std_logic_vector(46, 8),
18852 => conv_std_logic_vector(46, 8),
18853 => conv_std_logic_vector(47, 8),
18854 => conv_std_logic_vector(47, 8),
18855 => conv_std_logic_vector(47, 8),
18856 => conv_std_logic_vector(47, 8),
18857 => conv_std_logic_vector(48, 8),
18858 => conv_std_logic_vector(48, 8),
18859 => conv_std_logic_vector(48, 8),
18860 => conv_std_logic_vector(49, 8),
18861 => conv_std_logic_vector(49, 8),
18862 => conv_std_logic_vector(49, 8),
18863 => conv_std_logic_vector(49, 8),
18864 => conv_std_logic_vector(50, 8),
18865 => conv_std_logic_vector(50, 8),
18866 => conv_std_logic_vector(50, 8),
18867 => conv_std_logic_vector(51, 8),
18868 => conv_std_logic_vector(51, 8),
18869 => conv_std_logic_vector(51, 8),
18870 => conv_std_logic_vector(51, 8),
18871 => conv_std_logic_vector(52, 8),
18872 => conv_std_logic_vector(52, 8),
18873 => conv_std_logic_vector(52, 8),
18874 => conv_std_logic_vector(53, 8),
18875 => conv_std_logic_vector(53, 8),
18876 => conv_std_logic_vector(53, 8),
18877 => conv_std_logic_vector(53, 8),
18878 => conv_std_logic_vector(54, 8),
18879 => conv_std_logic_vector(54, 8),
18880 => conv_std_logic_vector(54, 8),
18881 => conv_std_logic_vector(55, 8),
18882 => conv_std_logic_vector(55, 8),
18883 => conv_std_logic_vector(55, 8),
18884 => conv_std_logic_vector(55, 8),
18885 => conv_std_logic_vector(56, 8),
18886 => conv_std_logic_vector(56, 8),
18887 => conv_std_logic_vector(56, 8),
18888 => conv_std_logic_vector(57, 8),
18889 => conv_std_logic_vector(57, 8),
18890 => conv_std_logic_vector(57, 8),
18891 => conv_std_logic_vector(57, 8),
18892 => conv_std_logic_vector(58, 8),
18893 => conv_std_logic_vector(58, 8),
18894 => conv_std_logic_vector(58, 8),
18895 => conv_std_logic_vector(59, 8),
18896 => conv_std_logic_vector(59, 8),
18897 => conv_std_logic_vector(59, 8),
18898 => conv_std_logic_vector(59, 8),
18899 => conv_std_logic_vector(60, 8),
18900 => conv_std_logic_vector(60, 8),
18901 => conv_std_logic_vector(60, 8),
18902 => conv_std_logic_vector(61, 8),
18903 => conv_std_logic_vector(61, 8),
18904 => conv_std_logic_vector(61, 8),
18905 => conv_std_logic_vector(61, 8),
18906 => conv_std_logic_vector(62, 8),
18907 => conv_std_logic_vector(62, 8),
18908 => conv_std_logic_vector(62, 8),
18909 => conv_std_logic_vector(63, 8),
18910 => conv_std_logic_vector(63, 8),
18911 => conv_std_logic_vector(63, 8),
18912 => conv_std_logic_vector(63, 8),
18913 => conv_std_logic_vector(64, 8),
18914 => conv_std_logic_vector(64, 8),
18915 => conv_std_logic_vector(64, 8),
18916 => conv_std_logic_vector(65, 8),
18917 => conv_std_logic_vector(65, 8),
18918 => conv_std_logic_vector(65, 8),
18919 => conv_std_logic_vector(65, 8),
18920 => conv_std_logic_vector(66, 8),
18921 => conv_std_logic_vector(66, 8),
18922 => conv_std_logic_vector(66, 8),
18923 => conv_std_logic_vector(67, 8),
18924 => conv_std_logic_vector(67, 8),
18925 => conv_std_logic_vector(67, 8),
18926 => conv_std_logic_vector(67, 8),
18927 => conv_std_logic_vector(68, 8),
18928 => conv_std_logic_vector(68, 8),
18929 => conv_std_logic_vector(68, 8),
18930 => conv_std_logic_vector(69, 8),
18931 => conv_std_logic_vector(69, 8),
18932 => conv_std_logic_vector(69, 8),
18933 => conv_std_logic_vector(69, 8),
18934 => conv_std_logic_vector(70, 8),
18935 => conv_std_logic_vector(70, 8),
18936 => conv_std_logic_vector(70, 8),
18937 => conv_std_logic_vector(71, 8),
18938 => conv_std_logic_vector(71, 8),
18939 => conv_std_logic_vector(71, 8),
18940 => conv_std_logic_vector(71, 8),
18941 => conv_std_logic_vector(72, 8),
18942 => conv_std_logic_vector(72, 8),
18943 => conv_std_logic_vector(72, 8),
18944 => conv_std_logic_vector(0, 8),
18945 => conv_std_logic_vector(0, 8),
18946 => conv_std_logic_vector(0, 8),
18947 => conv_std_logic_vector(0, 8),
18948 => conv_std_logic_vector(1, 8),
18949 => conv_std_logic_vector(1, 8),
18950 => conv_std_logic_vector(1, 8),
18951 => conv_std_logic_vector(2, 8),
18952 => conv_std_logic_vector(2, 8),
18953 => conv_std_logic_vector(2, 8),
18954 => conv_std_logic_vector(2, 8),
18955 => conv_std_logic_vector(3, 8),
18956 => conv_std_logic_vector(3, 8),
18957 => conv_std_logic_vector(3, 8),
18958 => conv_std_logic_vector(4, 8),
18959 => conv_std_logic_vector(4, 8),
18960 => conv_std_logic_vector(4, 8),
18961 => conv_std_logic_vector(4, 8),
18962 => conv_std_logic_vector(5, 8),
18963 => conv_std_logic_vector(5, 8),
18964 => conv_std_logic_vector(5, 8),
18965 => conv_std_logic_vector(6, 8),
18966 => conv_std_logic_vector(6, 8),
18967 => conv_std_logic_vector(6, 8),
18968 => conv_std_logic_vector(6, 8),
18969 => conv_std_logic_vector(7, 8),
18970 => conv_std_logic_vector(7, 8),
18971 => conv_std_logic_vector(7, 8),
18972 => conv_std_logic_vector(8, 8),
18973 => conv_std_logic_vector(8, 8),
18974 => conv_std_logic_vector(8, 8),
18975 => conv_std_logic_vector(8, 8),
18976 => conv_std_logic_vector(9, 8),
18977 => conv_std_logic_vector(9, 8),
18978 => conv_std_logic_vector(9, 8),
18979 => conv_std_logic_vector(10, 8),
18980 => conv_std_logic_vector(10, 8),
18981 => conv_std_logic_vector(10, 8),
18982 => conv_std_logic_vector(10, 8),
18983 => conv_std_logic_vector(11, 8),
18984 => conv_std_logic_vector(11, 8),
18985 => conv_std_logic_vector(11, 8),
18986 => conv_std_logic_vector(12, 8),
18987 => conv_std_logic_vector(12, 8),
18988 => conv_std_logic_vector(12, 8),
18989 => conv_std_logic_vector(13, 8),
18990 => conv_std_logic_vector(13, 8),
18991 => conv_std_logic_vector(13, 8),
18992 => conv_std_logic_vector(13, 8),
18993 => conv_std_logic_vector(14, 8),
18994 => conv_std_logic_vector(14, 8),
18995 => conv_std_logic_vector(14, 8),
18996 => conv_std_logic_vector(15, 8),
18997 => conv_std_logic_vector(15, 8),
18998 => conv_std_logic_vector(15, 8),
18999 => conv_std_logic_vector(15, 8),
19000 => conv_std_logic_vector(16, 8),
19001 => conv_std_logic_vector(16, 8),
19002 => conv_std_logic_vector(16, 8),
19003 => conv_std_logic_vector(17, 8),
19004 => conv_std_logic_vector(17, 8),
19005 => conv_std_logic_vector(17, 8),
19006 => conv_std_logic_vector(17, 8),
19007 => conv_std_logic_vector(18, 8),
19008 => conv_std_logic_vector(18, 8),
19009 => conv_std_logic_vector(18, 8),
19010 => conv_std_logic_vector(19, 8),
19011 => conv_std_logic_vector(19, 8),
19012 => conv_std_logic_vector(19, 8),
19013 => conv_std_logic_vector(19, 8),
19014 => conv_std_logic_vector(20, 8),
19015 => conv_std_logic_vector(20, 8),
19016 => conv_std_logic_vector(20, 8),
19017 => conv_std_logic_vector(21, 8),
19018 => conv_std_logic_vector(21, 8),
19019 => conv_std_logic_vector(21, 8),
19020 => conv_std_logic_vector(21, 8),
19021 => conv_std_logic_vector(22, 8),
19022 => conv_std_logic_vector(22, 8),
19023 => conv_std_logic_vector(22, 8),
19024 => conv_std_logic_vector(23, 8),
19025 => conv_std_logic_vector(23, 8),
19026 => conv_std_logic_vector(23, 8),
19027 => conv_std_logic_vector(23, 8),
19028 => conv_std_logic_vector(24, 8),
19029 => conv_std_logic_vector(24, 8),
19030 => conv_std_logic_vector(24, 8),
19031 => conv_std_logic_vector(25, 8),
19032 => conv_std_logic_vector(25, 8),
19033 => conv_std_logic_vector(25, 8),
19034 => conv_std_logic_vector(26, 8),
19035 => conv_std_logic_vector(26, 8),
19036 => conv_std_logic_vector(26, 8),
19037 => conv_std_logic_vector(26, 8),
19038 => conv_std_logic_vector(27, 8),
19039 => conv_std_logic_vector(27, 8),
19040 => conv_std_logic_vector(27, 8),
19041 => conv_std_logic_vector(28, 8),
19042 => conv_std_logic_vector(28, 8),
19043 => conv_std_logic_vector(28, 8),
19044 => conv_std_logic_vector(28, 8),
19045 => conv_std_logic_vector(29, 8),
19046 => conv_std_logic_vector(29, 8),
19047 => conv_std_logic_vector(29, 8),
19048 => conv_std_logic_vector(30, 8),
19049 => conv_std_logic_vector(30, 8),
19050 => conv_std_logic_vector(30, 8),
19051 => conv_std_logic_vector(30, 8),
19052 => conv_std_logic_vector(31, 8),
19053 => conv_std_logic_vector(31, 8),
19054 => conv_std_logic_vector(31, 8),
19055 => conv_std_logic_vector(32, 8),
19056 => conv_std_logic_vector(32, 8),
19057 => conv_std_logic_vector(32, 8),
19058 => conv_std_logic_vector(32, 8),
19059 => conv_std_logic_vector(33, 8),
19060 => conv_std_logic_vector(33, 8),
19061 => conv_std_logic_vector(33, 8),
19062 => conv_std_logic_vector(34, 8),
19063 => conv_std_logic_vector(34, 8),
19064 => conv_std_logic_vector(34, 8),
19065 => conv_std_logic_vector(34, 8),
19066 => conv_std_logic_vector(35, 8),
19067 => conv_std_logic_vector(35, 8),
19068 => conv_std_logic_vector(35, 8),
19069 => conv_std_logic_vector(36, 8),
19070 => conv_std_logic_vector(36, 8),
19071 => conv_std_logic_vector(36, 8),
19072 => conv_std_logic_vector(37, 8),
19073 => conv_std_logic_vector(37, 8),
19074 => conv_std_logic_vector(37, 8),
19075 => conv_std_logic_vector(37, 8),
19076 => conv_std_logic_vector(38, 8),
19077 => conv_std_logic_vector(38, 8),
19078 => conv_std_logic_vector(38, 8),
19079 => conv_std_logic_vector(39, 8),
19080 => conv_std_logic_vector(39, 8),
19081 => conv_std_logic_vector(39, 8),
19082 => conv_std_logic_vector(39, 8),
19083 => conv_std_logic_vector(40, 8),
19084 => conv_std_logic_vector(40, 8),
19085 => conv_std_logic_vector(40, 8),
19086 => conv_std_logic_vector(41, 8),
19087 => conv_std_logic_vector(41, 8),
19088 => conv_std_logic_vector(41, 8),
19089 => conv_std_logic_vector(41, 8),
19090 => conv_std_logic_vector(42, 8),
19091 => conv_std_logic_vector(42, 8),
19092 => conv_std_logic_vector(42, 8),
19093 => conv_std_logic_vector(43, 8),
19094 => conv_std_logic_vector(43, 8),
19095 => conv_std_logic_vector(43, 8),
19096 => conv_std_logic_vector(43, 8),
19097 => conv_std_logic_vector(44, 8),
19098 => conv_std_logic_vector(44, 8),
19099 => conv_std_logic_vector(44, 8),
19100 => conv_std_logic_vector(45, 8),
19101 => conv_std_logic_vector(45, 8),
19102 => conv_std_logic_vector(45, 8),
19103 => conv_std_logic_vector(45, 8),
19104 => conv_std_logic_vector(46, 8),
19105 => conv_std_logic_vector(46, 8),
19106 => conv_std_logic_vector(46, 8),
19107 => conv_std_logic_vector(47, 8),
19108 => conv_std_logic_vector(47, 8),
19109 => conv_std_logic_vector(47, 8),
19110 => conv_std_logic_vector(47, 8),
19111 => conv_std_logic_vector(48, 8),
19112 => conv_std_logic_vector(48, 8),
19113 => conv_std_logic_vector(48, 8),
19114 => conv_std_logic_vector(49, 8),
19115 => conv_std_logic_vector(49, 8),
19116 => conv_std_logic_vector(49, 8),
19117 => conv_std_logic_vector(50, 8),
19118 => conv_std_logic_vector(50, 8),
19119 => conv_std_logic_vector(50, 8),
19120 => conv_std_logic_vector(50, 8),
19121 => conv_std_logic_vector(51, 8),
19122 => conv_std_logic_vector(51, 8),
19123 => conv_std_logic_vector(51, 8),
19124 => conv_std_logic_vector(52, 8),
19125 => conv_std_logic_vector(52, 8),
19126 => conv_std_logic_vector(52, 8),
19127 => conv_std_logic_vector(52, 8),
19128 => conv_std_logic_vector(53, 8),
19129 => conv_std_logic_vector(53, 8),
19130 => conv_std_logic_vector(53, 8),
19131 => conv_std_logic_vector(54, 8),
19132 => conv_std_logic_vector(54, 8),
19133 => conv_std_logic_vector(54, 8),
19134 => conv_std_logic_vector(54, 8),
19135 => conv_std_logic_vector(55, 8),
19136 => conv_std_logic_vector(55, 8),
19137 => conv_std_logic_vector(55, 8),
19138 => conv_std_logic_vector(56, 8),
19139 => conv_std_logic_vector(56, 8),
19140 => conv_std_logic_vector(56, 8),
19141 => conv_std_logic_vector(56, 8),
19142 => conv_std_logic_vector(57, 8),
19143 => conv_std_logic_vector(57, 8),
19144 => conv_std_logic_vector(57, 8),
19145 => conv_std_logic_vector(58, 8),
19146 => conv_std_logic_vector(58, 8),
19147 => conv_std_logic_vector(58, 8),
19148 => conv_std_logic_vector(58, 8),
19149 => conv_std_logic_vector(59, 8),
19150 => conv_std_logic_vector(59, 8),
19151 => conv_std_logic_vector(59, 8),
19152 => conv_std_logic_vector(60, 8),
19153 => conv_std_logic_vector(60, 8),
19154 => conv_std_logic_vector(60, 8),
19155 => conv_std_logic_vector(60, 8),
19156 => conv_std_logic_vector(61, 8),
19157 => conv_std_logic_vector(61, 8),
19158 => conv_std_logic_vector(61, 8),
19159 => conv_std_logic_vector(62, 8),
19160 => conv_std_logic_vector(62, 8),
19161 => conv_std_logic_vector(62, 8),
19162 => conv_std_logic_vector(63, 8),
19163 => conv_std_logic_vector(63, 8),
19164 => conv_std_logic_vector(63, 8),
19165 => conv_std_logic_vector(63, 8),
19166 => conv_std_logic_vector(64, 8),
19167 => conv_std_logic_vector(64, 8),
19168 => conv_std_logic_vector(64, 8),
19169 => conv_std_logic_vector(65, 8),
19170 => conv_std_logic_vector(65, 8),
19171 => conv_std_logic_vector(65, 8),
19172 => conv_std_logic_vector(65, 8),
19173 => conv_std_logic_vector(66, 8),
19174 => conv_std_logic_vector(66, 8),
19175 => conv_std_logic_vector(66, 8),
19176 => conv_std_logic_vector(67, 8),
19177 => conv_std_logic_vector(67, 8),
19178 => conv_std_logic_vector(67, 8),
19179 => conv_std_logic_vector(67, 8),
19180 => conv_std_logic_vector(68, 8),
19181 => conv_std_logic_vector(68, 8),
19182 => conv_std_logic_vector(68, 8),
19183 => conv_std_logic_vector(69, 8),
19184 => conv_std_logic_vector(69, 8),
19185 => conv_std_logic_vector(69, 8),
19186 => conv_std_logic_vector(69, 8),
19187 => conv_std_logic_vector(70, 8),
19188 => conv_std_logic_vector(70, 8),
19189 => conv_std_logic_vector(70, 8),
19190 => conv_std_logic_vector(71, 8),
19191 => conv_std_logic_vector(71, 8),
19192 => conv_std_logic_vector(71, 8),
19193 => conv_std_logic_vector(71, 8),
19194 => conv_std_logic_vector(72, 8),
19195 => conv_std_logic_vector(72, 8),
19196 => conv_std_logic_vector(72, 8),
19197 => conv_std_logic_vector(73, 8),
19198 => conv_std_logic_vector(73, 8),
19199 => conv_std_logic_vector(73, 8),
19200 => conv_std_logic_vector(0, 8),
19201 => conv_std_logic_vector(0, 8),
19202 => conv_std_logic_vector(0, 8),
19203 => conv_std_logic_vector(0, 8),
19204 => conv_std_logic_vector(1, 8),
19205 => conv_std_logic_vector(1, 8),
19206 => conv_std_logic_vector(1, 8),
19207 => conv_std_logic_vector(2, 8),
19208 => conv_std_logic_vector(2, 8),
19209 => conv_std_logic_vector(2, 8),
19210 => conv_std_logic_vector(2, 8),
19211 => conv_std_logic_vector(3, 8),
19212 => conv_std_logic_vector(3, 8),
19213 => conv_std_logic_vector(3, 8),
19214 => conv_std_logic_vector(4, 8),
19215 => conv_std_logic_vector(4, 8),
19216 => conv_std_logic_vector(4, 8),
19217 => conv_std_logic_vector(4, 8),
19218 => conv_std_logic_vector(5, 8),
19219 => conv_std_logic_vector(5, 8),
19220 => conv_std_logic_vector(5, 8),
19221 => conv_std_logic_vector(6, 8),
19222 => conv_std_logic_vector(6, 8),
19223 => conv_std_logic_vector(6, 8),
19224 => conv_std_logic_vector(7, 8),
19225 => conv_std_logic_vector(7, 8),
19226 => conv_std_logic_vector(7, 8),
19227 => conv_std_logic_vector(7, 8),
19228 => conv_std_logic_vector(8, 8),
19229 => conv_std_logic_vector(8, 8),
19230 => conv_std_logic_vector(8, 8),
19231 => conv_std_logic_vector(9, 8),
19232 => conv_std_logic_vector(9, 8),
19233 => conv_std_logic_vector(9, 8),
19234 => conv_std_logic_vector(9, 8),
19235 => conv_std_logic_vector(10, 8),
19236 => conv_std_logic_vector(10, 8),
19237 => conv_std_logic_vector(10, 8),
19238 => conv_std_logic_vector(11, 8),
19239 => conv_std_logic_vector(11, 8),
19240 => conv_std_logic_vector(11, 8),
19241 => conv_std_logic_vector(12, 8),
19242 => conv_std_logic_vector(12, 8),
19243 => conv_std_logic_vector(12, 8),
19244 => conv_std_logic_vector(12, 8),
19245 => conv_std_logic_vector(13, 8),
19246 => conv_std_logic_vector(13, 8),
19247 => conv_std_logic_vector(13, 8),
19248 => conv_std_logic_vector(14, 8),
19249 => conv_std_logic_vector(14, 8),
19250 => conv_std_logic_vector(14, 8),
19251 => conv_std_logic_vector(14, 8),
19252 => conv_std_logic_vector(15, 8),
19253 => conv_std_logic_vector(15, 8),
19254 => conv_std_logic_vector(15, 8),
19255 => conv_std_logic_vector(16, 8),
19256 => conv_std_logic_vector(16, 8),
19257 => conv_std_logic_vector(16, 8),
19258 => conv_std_logic_vector(16, 8),
19259 => conv_std_logic_vector(17, 8),
19260 => conv_std_logic_vector(17, 8),
19261 => conv_std_logic_vector(17, 8),
19262 => conv_std_logic_vector(18, 8),
19263 => conv_std_logic_vector(18, 8),
19264 => conv_std_logic_vector(18, 8),
19265 => conv_std_logic_vector(19, 8),
19266 => conv_std_logic_vector(19, 8),
19267 => conv_std_logic_vector(19, 8),
19268 => conv_std_logic_vector(19, 8),
19269 => conv_std_logic_vector(20, 8),
19270 => conv_std_logic_vector(20, 8),
19271 => conv_std_logic_vector(20, 8),
19272 => conv_std_logic_vector(21, 8),
19273 => conv_std_logic_vector(21, 8),
19274 => conv_std_logic_vector(21, 8),
19275 => conv_std_logic_vector(21, 8),
19276 => conv_std_logic_vector(22, 8),
19277 => conv_std_logic_vector(22, 8),
19278 => conv_std_logic_vector(22, 8),
19279 => conv_std_logic_vector(23, 8),
19280 => conv_std_logic_vector(23, 8),
19281 => conv_std_logic_vector(23, 8),
19282 => conv_std_logic_vector(24, 8),
19283 => conv_std_logic_vector(24, 8),
19284 => conv_std_logic_vector(24, 8),
19285 => conv_std_logic_vector(24, 8),
19286 => conv_std_logic_vector(25, 8),
19287 => conv_std_logic_vector(25, 8),
19288 => conv_std_logic_vector(25, 8),
19289 => conv_std_logic_vector(26, 8),
19290 => conv_std_logic_vector(26, 8),
19291 => conv_std_logic_vector(26, 8),
19292 => conv_std_logic_vector(26, 8),
19293 => conv_std_logic_vector(27, 8),
19294 => conv_std_logic_vector(27, 8),
19295 => conv_std_logic_vector(27, 8),
19296 => conv_std_logic_vector(28, 8),
19297 => conv_std_logic_vector(28, 8),
19298 => conv_std_logic_vector(28, 8),
19299 => conv_std_logic_vector(29, 8),
19300 => conv_std_logic_vector(29, 8),
19301 => conv_std_logic_vector(29, 8),
19302 => conv_std_logic_vector(29, 8),
19303 => conv_std_logic_vector(30, 8),
19304 => conv_std_logic_vector(30, 8),
19305 => conv_std_logic_vector(30, 8),
19306 => conv_std_logic_vector(31, 8),
19307 => conv_std_logic_vector(31, 8),
19308 => conv_std_logic_vector(31, 8),
19309 => conv_std_logic_vector(31, 8),
19310 => conv_std_logic_vector(32, 8),
19311 => conv_std_logic_vector(32, 8),
19312 => conv_std_logic_vector(32, 8),
19313 => conv_std_logic_vector(33, 8),
19314 => conv_std_logic_vector(33, 8),
19315 => conv_std_logic_vector(33, 8),
19316 => conv_std_logic_vector(33, 8),
19317 => conv_std_logic_vector(34, 8),
19318 => conv_std_logic_vector(34, 8),
19319 => conv_std_logic_vector(34, 8),
19320 => conv_std_logic_vector(35, 8),
19321 => conv_std_logic_vector(35, 8),
19322 => conv_std_logic_vector(35, 8),
19323 => conv_std_logic_vector(36, 8),
19324 => conv_std_logic_vector(36, 8),
19325 => conv_std_logic_vector(36, 8),
19326 => conv_std_logic_vector(36, 8),
19327 => conv_std_logic_vector(37, 8),
19328 => conv_std_logic_vector(37, 8),
19329 => conv_std_logic_vector(37, 8),
19330 => conv_std_logic_vector(38, 8),
19331 => conv_std_logic_vector(38, 8),
19332 => conv_std_logic_vector(38, 8),
19333 => conv_std_logic_vector(38, 8),
19334 => conv_std_logic_vector(39, 8),
19335 => conv_std_logic_vector(39, 8),
19336 => conv_std_logic_vector(39, 8),
19337 => conv_std_logic_vector(40, 8),
19338 => conv_std_logic_vector(40, 8),
19339 => conv_std_logic_vector(40, 8),
19340 => conv_std_logic_vector(41, 8),
19341 => conv_std_logic_vector(41, 8),
19342 => conv_std_logic_vector(41, 8),
19343 => conv_std_logic_vector(41, 8),
19344 => conv_std_logic_vector(42, 8),
19345 => conv_std_logic_vector(42, 8),
19346 => conv_std_logic_vector(42, 8),
19347 => conv_std_logic_vector(43, 8),
19348 => conv_std_logic_vector(43, 8),
19349 => conv_std_logic_vector(43, 8),
19350 => conv_std_logic_vector(43, 8),
19351 => conv_std_logic_vector(44, 8),
19352 => conv_std_logic_vector(44, 8),
19353 => conv_std_logic_vector(44, 8),
19354 => conv_std_logic_vector(45, 8),
19355 => conv_std_logic_vector(45, 8),
19356 => conv_std_logic_vector(45, 8),
19357 => conv_std_logic_vector(45, 8),
19358 => conv_std_logic_vector(46, 8),
19359 => conv_std_logic_vector(46, 8),
19360 => conv_std_logic_vector(46, 8),
19361 => conv_std_logic_vector(47, 8),
19362 => conv_std_logic_vector(47, 8),
19363 => conv_std_logic_vector(47, 8),
19364 => conv_std_logic_vector(48, 8),
19365 => conv_std_logic_vector(48, 8),
19366 => conv_std_logic_vector(48, 8),
19367 => conv_std_logic_vector(48, 8),
19368 => conv_std_logic_vector(49, 8),
19369 => conv_std_logic_vector(49, 8),
19370 => conv_std_logic_vector(49, 8),
19371 => conv_std_logic_vector(50, 8),
19372 => conv_std_logic_vector(50, 8),
19373 => conv_std_logic_vector(50, 8),
19374 => conv_std_logic_vector(50, 8),
19375 => conv_std_logic_vector(51, 8),
19376 => conv_std_logic_vector(51, 8),
19377 => conv_std_logic_vector(51, 8),
19378 => conv_std_logic_vector(52, 8),
19379 => conv_std_logic_vector(52, 8),
19380 => conv_std_logic_vector(52, 8),
19381 => conv_std_logic_vector(53, 8),
19382 => conv_std_logic_vector(53, 8),
19383 => conv_std_logic_vector(53, 8),
19384 => conv_std_logic_vector(53, 8),
19385 => conv_std_logic_vector(54, 8),
19386 => conv_std_logic_vector(54, 8),
19387 => conv_std_logic_vector(54, 8),
19388 => conv_std_logic_vector(55, 8),
19389 => conv_std_logic_vector(55, 8),
19390 => conv_std_logic_vector(55, 8),
19391 => conv_std_logic_vector(55, 8),
19392 => conv_std_logic_vector(56, 8),
19393 => conv_std_logic_vector(56, 8),
19394 => conv_std_logic_vector(56, 8),
19395 => conv_std_logic_vector(57, 8),
19396 => conv_std_logic_vector(57, 8),
19397 => conv_std_logic_vector(57, 8),
19398 => conv_std_logic_vector(58, 8),
19399 => conv_std_logic_vector(58, 8),
19400 => conv_std_logic_vector(58, 8),
19401 => conv_std_logic_vector(58, 8),
19402 => conv_std_logic_vector(59, 8),
19403 => conv_std_logic_vector(59, 8),
19404 => conv_std_logic_vector(59, 8),
19405 => conv_std_logic_vector(60, 8),
19406 => conv_std_logic_vector(60, 8),
19407 => conv_std_logic_vector(60, 8),
19408 => conv_std_logic_vector(60, 8),
19409 => conv_std_logic_vector(61, 8),
19410 => conv_std_logic_vector(61, 8),
19411 => conv_std_logic_vector(61, 8),
19412 => conv_std_logic_vector(62, 8),
19413 => conv_std_logic_vector(62, 8),
19414 => conv_std_logic_vector(62, 8),
19415 => conv_std_logic_vector(62, 8),
19416 => conv_std_logic_vector(63, 8),
19417 => conv_std_logic_vector(63, 8),
19418 => conv_std_logic_vector(63, 8),
19419 => conv_std_logic_vector(64, 8),
19420 => conv_std_logic_vector(64, 8),
19421 => conv_std_logic_vector(64, 8),
19422 => conv_std_logic_vector(65, 8),
19423 => conv_std_logic_vector(65, 8),
19424 => conv_std_logic_vector(65, 8),
19425 => conv_std_logic_vector(65, 8),
19426 => conv_std_logic_vector(66, 8),
19427 => conv_std_logic_vector(66, 8),
19428 => conv_std_logic_vector(66, 8),
19429 => conv_std_logic_vector(67, 8),
19430 => conv_std_logic_vector(67, 8),
19431 => conv_std_logic_vector(67, 8),
19432 => conv_std_logic_vector(67, 8),
19433 => conv_std_logic_vector(68, 8),
19434 => conv_std_logic_vector(68, 8),
19435 => conv_std_logic_vector(68, 8),
19436 => conv_std_logic_vector(69, 8),
19437 => conv_std_logic_vector(69, 8),
19438 => conv_std_logic_vector(69, 8),
19439 => conv_std_logic_vector(70, 8),
19440 => conv_std_logic_vector(70, 8),
19441 => conv_std_logic_vector(70, 8),
19442 => conv_std_logic_vector(70, 8),
19443 => conv_std_logic_vector(71, 8),
19444 => conv_std_logic_vector(71, 8),
19445 => conv_std_logic_vector(71, 8),
19446 => conv_std_logic_vector(72, 8),
19447 => conv_std_logic_vector(72, 8),
19448 => conv_std_logic_vector(72, 8),
19449 => conv_std_logic_vector(72, 8),
19450 => conv_std_logic_vector(73, 8),
19451 => conv_std_logic_vector(73, 8),
19452 => conv_std_logic_vector(73, 8),
19453 => conv_std_logic_vector(74, 8),
19454 => conv_std_logic_vector(74, 8),
19455 => conv_std_logic_vector(74, 8),
19456 => conv_std_logic_vector(0, 8),
19457 => conv_std_logic_vector(0, 8),
19458 => conv_std_logic_vector(0, 8),
19459 => conv_std_logic_vector(0, 8),
19460 => conv_std_logic_vector(1, 8),
19461 => conv_std_logic_vector(1, 8),
19462 => conv_std_logic_vector(1, 8),
19463 => conv_std_logic_vector(2, 8),
19464 => conv_std_logic_vector(2, 8),
19465 => conv_std_logic_vector(2, 8),
19466 => conv_std_logic_vector(2, 8),
19467 => conv_std_logic_vector(3, 8),
19468 => conv_std_logic_vector(3, 8),
19469 => conv_std_logic_vector(3, 8),
19470 => conv_std_logic_vector(4, 8),
19471 => conv_std_logic_vector(4, 8),
19472 => conv_std_logic_vector(4, 8),
19473 => conv_std_logic_vector(5, 8),
19474 => conv_std_logic_vector(5, 8),
19475 => conv_std_logic_vector(5, 8),
19476 => conv_std_logic_vector(5, 8),
19477 => conv_std_logic_vector(6, 8),
19478 => conv_std_logic_vector(6, 8),
19479 => conv_std_logic_vector(6, 8),
19480 => conv_std_logic_vector(7, 8),
19481 => conv_std_logic_vector(7, 8),
19482 => conv_std_logic_vector(7, 8),
19483 => conv_std_logic_vector(8, 8),
19484 => conv_std_logic_vector(8, 8),
19485 => conv_std_logic_vector(8, 8),
19486 => conv_std_logic_vector(8, 8),
19487 => conv_std_logic_vector(9, 8),
19488 => conv_std_logic_vector(9, 8),
19489 => conv_std_logic_vector(9, 8),
19490 => conv_std_logic_vector(10, 8),
19491 => conv_std_logic_vector(10, 8),
19492 => conv_std_logic_vector(10, 8),
19493 => conv_std_logic_vector(10, 8),
19494 => conv_std_logic_vector(11, 8),
19495 => conv_std_logic_vector(11, 8),
19496 => conv_std_logic_vector(11, 8),
19497 => conv_std_logic_vector(12, 8),
19498 => conv_std_logic_vector(12, 8),
19499 => conv_std_logic_vector(12, 8),
19500 => conv_std_logic_vector(13, 8),
19501 => conv_std_logic_vector(13, 8),
19502 => conv_std_logic_vector(13, 8),
19503 => conv_std_logic_vector(13, 8),
19504 => conv_std_logic_vector(14, 8),
19505 => conv_std_logic_vector(14, 8),
19506 => conv_std_logic_vector(14, 8),
19507 => conv_std_logic_vector(15, 8),
19508 => conv_std_logic_vector(15, 8),
19509 => conv_std_logic_vector(15, 8),
19510 => conv_std_logic_vector(16, 8),
19511 => conv_std_logic_vector(16, 8),
19512 => conv_std_logic_vector(16, 8),
19513 => conv_std_logic_vector(16, 8),
19514 => conv_std_logic_vector(17, 8),
19515 => conv_std_logic_vector(17, 8),
19516 => conv_std_logic_vector(17, 8),
19517 => conv_std_logic_vector(18, 8),
19518 => conv_std_logic_vector(18, 8),
19519 => conv_std_logic_vector(18, 8),
19520 => conv_std_logic_vector(19, 8),
19521 => conv_std_logic_vector(19, 8),
19522 => conv_std_logic_vector(19, 8),
19523 => conv_std_logic_vector(19, 8),
19524 => conv_std_logic_vector(20, 8),
19525 => conv_std_logic_vector(20, 8),
19526 => conv_std_logic_vector(20, 8),
19527 => conv_std_logic_vector(21, 8),
19528 => conv_std_logic_vector(21, 8),
19529 => conv_std_logic_vector(21, 8),
19530 => conv_std_logic_vector(21, 8),
19531 => conv_std_logic_vector(22, 8),
19532 => conv_std_logic_vector(22, 8),
19533 => conv_std_logic_vector(22, 8),
19534 => conv_std_logic_vector(23, 8),
19535 => conv_std_logic_vector(23, 8),
19536 => conv_std_logic_vector(23, 8),
19537 => conv_std_logic_vector(24, 8),
19538 => conv_std_logic_vector(24, 8),
19539 => conv_std_logic_vector(24, 8),
19540 => conv_std_logic_vector(24, 8),
19541 => conv_std_logic_vector(25, 8),
19542 => conv_std_logic_vector(25, 8),
19543 => conv_std_logic_vector(25, 8),
19544 => conv_std_logic_vector(26, 8),
19545 => conv_std_logic_vector(26, 8),
19546 => conv_std_logic_vector(26, 8),
19547 => conv_std_logic_vector(27, 8),
19548 => conv_std_logic_vector(27, 8),
19549 => conv_std_logic_vector(27, 8),
19550 => conv_std_logic_vector(27, 8),
19551 => conv_std_logic_vector(28, 8),
19552 => conv_std_logic_vector(28, 8),
19553 => conv_std_logic_vector(28, 8),
19554 => conv_std_logic_vector(29, 8),
19555 => conv_std_logic_vector(29, 8),
19556 => conv_std_logic_vector(29, 8),
19557 => conv_std_logic_vector(29, 8),
19558 => conv_std_logic_vector(30, 8),
19559 => conv_std_logic_vector(30, 8),
19560 => conv_std_logic_vector(30, 8),
19561 => conv_std_logic_vector(31, 8),
19562 => conv_std_logic_vector(31, 8),
19563 => conv_std_logic_vector(31, 8),
19564 => conv_std_logic_vector(32, 8),
19565 => conv_std_logic_vector(32, 8),
19566 => conv_std_logic_vector(32, 8),
19567 => conv_std_logic_vector(32, 8),
19568 => conv_std_logic_vector(33, 8),
19569 => conv_std_logic_vector(33, 8),
19570 => conv_std_logic_vector(33, 8),
19571 => conv_std_logic_vector(34, 8),
19572 => conv_std_logic_vector(34, 8),
19573 => conv_std_logic_vector(34, 8),
19574 => conv_std_logic_vector(35, 8),
19575 => conv_std_logic_vector(35, 8),
19576 => conv_std_logic_vector(35, 8),
19577 => conv_std_logic_vector(35, 8),
19578 => conv_std_logic_vector(36, 8),
19579 => conv_std_logic_vector(36, 8),
19580 => conv_std_logic_vector(36, 8),
19581 => conv_std_logic_vector(37, 8),
19582 => conv_std_logic_vector(37, 8),
19583 => conv_std_logic_vector(37, 8),
19584 => conv_std_logic_vector(38, 8),
19585 => conv_std_logic_vector(38, 8),
19586 => conv_std_logic_vector(38, 8),
19587 => conv_std_logic_vector(38, 8),
19588 => conv_std_logic_vector(39, 8),
19589 => conv_std_logic_vector(39, 8),
19590 => conv_std_logic_vector(39, 8),
19591 => conv_std_logic_vector(40, 8),
19592 => conv_std_logic_vector(40, 8),
19593 => conv_std_logic_vector(40, 8),
19594 => conv_std_logic_vector(40, 8),
19595 => conv_std_logic_vector(41, 8),
19596 => conv_std_logic_vector(41, 8),
19597 => conv_std_logic_vector(41, 8),
19598 => conv_std_logic_vector(42, 8),
19599 => conv_std_logic_vector(42, 8),
19600 => conv_std_logic_vector(42, 8),
19601 => conv_std_logic_vector(43, 8),
19602 => conv_std_logic_vector(43, 8),
19603 => conv_std_logic_vector(43, 8),
19604 => conv_std_logic_vector(43, 8),
19605 => conv_std_logic_vector(44, 8),
19606 => conv_std_logic_vector(44, 8),
19607 => conv_std_logic_vector(44, 8),
19608 => conv_std_logic_vector(45, 8),
19609 => conv_std_logic_vector(45, 8),
19610 => conv_std_logic_vector(45, 8),
19611 => conv_std_logic_vector(46, 8),
19612 => conv_std_logic_vector(46, 8),
19613 => conv_std_logic_vector(46, 8),
19614 => conv_std_logic_vector(46, 8),
19615 => conv_std_logic_vector(47, 8),
19616 => conv_std_logic_vector(47, 8),
19617 => conv_std_logic_vector(47, 8),
19618 => conv_std_logic_vector(48, 8),
19619 => conv_std_logic_vector(48, 8),
19620 => conv_std_logic_vector(48, 8),
19621 => conv_std_logic_vector(48, 8),
19622 => conv_std_logic_vector(49, 8),
19623 => conv_std_logic_vector(49, 8),
19624 => conv_std_logic_vector(49, 8),
19625 => conv_std_logic_vector(50, 8),
19626 => conv_std_logic_vector(50, 8),
19627 => conv_std_logic_vector(50, 8),
19628 => conv_std_logic_vector(51, 8),
19629 => conv_std_logic_vector(51, 8),
19630 => conv_std_logic_vector(51, 8),
19631 => conv_std_logic_vector(51, 8),
19632 => conv_std_logic_vector(52, 8),
19633 => conv_std_logic_vector(52, 8),
19634 => conv_std_logic_vector(52, 8),
19635 => conv_std_logic_vector(53, 8),
19636 => conv_std_logic_vector(53, 8),
19637 => conv_std_logic_vector(53, 8),
19638 => conv_std_logic_vector(54, 8),
19639 => conv_std_logic_vector(54, 8),
19640 => conv_std_logic_vector(54, 8),
19641 => conv_std_logic_vector(54, 8),
19642 => conv_std_logic_vector(55, 8),
19643 => conv_std_logic_vector(55, 8),
19644 => conv_std_logic_vector(55, 8),
19645 => conv_std_logic_vector(56, 8),
19646 => conv_std_logic_vector(56, 8),
19647 => conv_std_logic_vector(56, 8),
19648 => conv_std_logic_vector(57, 8),
19649 => conv_std_logic_vector(57, 8),
19650 => conv_std_logic_vector(57, 8),
19651 => conv_std_logic_vector(57, 8),
19652 => conv_std_logic_vector(58, 8),
19653 => conv_std_logic_vector(58, 8),
19654 => conv_std_logic_vector(58, 8),
19655 => conv_std_logic_vector(59, 8),
19656 => conv_std_logic_vector(59, 8),
19657 => conv_std_logic_vector(59, 8),
19658 => conv_std_logic_vector(59, 8),
19659 => conv_std_logic_vector(60, 8),
19660 => conv_std_logic_vector(60, 8),
19661 => conv_std_logic_vector(60, 8),
19662 => conv_std_logic_vector(61, 8),
19663 => conv_std_logic_vector(61, 8),
19664 => conv_std_logic_vector(61, 8),
19665 => conv_std_logic_vector(62, 8),
19666 => conv_std_logic_vector(62, 8),
19667 => conv_std_logic_vector(62, 8),
19668 => conv_std_logic_vector(62, 8),
19669 => conv_std_logic_vector(63, 8),
19670 => conv_std_logic_vector(63, 8),
19671 => conv_std_logic_vector(63, 8),
19672 => conv_std_logic_vector(64, 8),
19673 => conv_std_logic_vector(64, 8),
19674 => conv_std_logic_vector(64, 8),
19675 => conv_std_logic_vector(65, 8),
19676 => conv_std_logic_vector(65, 8),
19677 => conv_std_logic_vector(65, 8),
19678 => conv_std_logic_vector(65, 8),
19679 => conv_std_logic_vector(66, 8),
19680 => conv_std_logic_vector(66, 8),
19681 => conv_std_logic_vector(66, 8),
19682 => conv_std_logic_vector(67, 8),
19683 => conv_std_logic_vector(67, 8),
19684 => conv_std_logic_vector(67, 8),
19685 => conv_std_logic_vector(67, 8),
19686 => conv_std_logic_vector(68, 8),
19687 => conv_std_logic_vector(68, 8),
19688 => conv_std_logic_vector(68, 8),
19689 => conv_std_logic_vector(69, 8),
19690 => conv_std_logic_vector(69, 8),
19691 => conv_std_logic_vector(69, 8),
19692 => conv_std_logic_vector(70, 8),
19693 => conv_std_logic_vector(70, 8),
19694 => conv_std_logic_vector(70, 8),
19695 => conv_std_logic_vector(70, 8),
19696 => conv_std_logic_vector(71, 8),
19697 => conv_std_logic_vector(71, 8),
19698 => conv_std_logic_vector(71, 8),
19699 => conv_std_logic_vector(72, 8),
19700 => conv_std_logic_vector(72, 8),
19701 => conv_std_logic_vector(72, 8),
19702 => conv_std_logic_vector(73, 8),
19703 => conv_std_logic_vector(73, 8),
19704 => conv_std_logic_vector(73, 8),
19705 => conv_std_logic_vector(73, 8),
19706 => conv_std_logic_vector(74, 8),
19707 => conv_std_logic_vector(74, 8),
19708 => conv_std_logic_vector(74, 8),
19709 => conv_std_logic_vector(75, 8),
19710 => conv_std_logic_vector(75, 8),
19711 => conv_std_logic_vector(75, 8),
19712 => conv_std_logic_vector(0, 8),
19713 => conv_std_logic_vector(0, 8),
19714 => conv_std_logic_vector(0, 8),
19715 => conv_std_logic_vector(0, 8),
19716 => conv_std_logic_vector(1, 8),
19717 => conv_std_logic_vector(1, 8),
19718 => conv_std_logic_vector(1, 8),
19719 => conv_std_logic_vector(2, 8),
19720 => conv_std_logic_vector(2, 8),
19721 => conv_std_logic_vector(2, 8),
19722 => conv_std_logic_vector(3, 8),
19723 => conv_std_logic_vector(3, 8),
19724 => conv_std_logic_vector(3, 8),
19725 => conv_std_logic_vector(3, 8),
19726 => conv_std_logic_vector(4, 8),
19727 => conv_std_logic_vector(4, 8),
19728 => conv_std_logic_vector(4, 8),
19729 => conv_std_logic_vector(5, 8),
19730 => conv_std_logic_vector(5, 8),
19731 => conv_std_logic_vector(5, 8),
19732 => conv_std_logic_vector(6, 8),
19733 => conv_std_logic_vector(6, 8),
19734 => conv_std_logic_vector(6, 8),
19735 => conv_std_logic_vector(6, 8),
19736 => conv_std_logic_vector(7, 8),
19737 => conv_std_logic_vector(7, 8),
19738 => conv_std_logic_vector(7, 8),
19739 => conv_std_logic_vector(8, 8),
19740 => conv_std_logic_vector(8, 8),
19741 => conv_std_logic_vector(8, 8),
19742 => conv_std_logic_vector(9, 8),
19743 => conv_std_logic_vector(9, 8),
19744 => conv_std_logic_vector(9, 8),
19745 => conv_std_logic_vector(9, 8),
19746 => conv_std_logic_vector(10, 8),
19747 => conv_std_logic_vector(10, 8),
19748 => conv_std_logic_vector(10, 8),
19749 => conv_std_logic_vector(11, 8),
19750 => conv_std_logic_vector(11, 8),
19751 => conv_std_logic_vector(11, 8),
19752 => conv_std_logic_vector(12, 8),
19753 => conv_std_logic_vector(12, 8),
19754 => conv_std_logic_vector(12, 8),
19755 => conv_std_logic_vector(12, 8),
19756 => conv_std_logic_vector(13, 8),
19757 => conv_std_logic_vector(13, 8),
19758 => conv_std_logic_vector(13, 8),
19759 => conv_std_logic_vector(14, 8),
19760 => conv_std_logic_vector(14, 8),
19761 => conv_std_logic_vector(14, 8),
19762 => conv_std_logic_vector(15, 8),
19763 => conv_std_logic_vector(15, 8),
19764 => conv_std_logic_vector(15, 8),
19765 => conv_std_logic_vector(15, 8),
19766 => conv_std_logic_vector(16, 8),
19767 => conv_std_logic_vector(16, 8),
19768 => conv_std_logic_vector(16, 8),
19769 => conv_std_logic_vector(17, 8),
19770 => conv_std_logic_vector(17, 8),
19771 => conv_std_logic_vector(17, 8),
19772 => conv_std_logic_vector(18, 8),
19773 => conv_std_logic_vector(18, 8),
19774 => conv_std_logic_vector(18, 8),
19775 => conv_std_logic_vector(18, 8),
19776 => conv_std_logic_vector(19, 8),
19777 => conv_std_logic_vector(19, 8),
19778 => conv_std_logic_vector(19, 8),
19779 => conv_std_logic_vector(20, 8),
19780 => conv_std_logic_vector(20, 8),
19781 => conv_std_logic_vector(20, 8),
19782 => conv_std_logic_vector(21, 8),
19783 => conv_std_logic_vector(21, 8),
19784 => conv_std_logic_vector(21, 8),
19785 => conv_std_logic_vector(21, 8),
19786 => conv_std_logic_vector(22, 8),
19787 => conv_std_logic_vector(22, 8),
19788 => conv_std_logic_vector(22, 8),
19789 => conv_std_logic_vector(23, 8),
19790 => conv_std_logic_vector(23, 8),
19791 => conv_std_logic_vector(23, 8),
19792 => conv_std_logic_vector(24, 8),
19793 => conv_std_logic_vector(24, 8),
19794 => conv_std_logic_vector(24, 8),
19795 => conv_std_logic_vector(24, 8),
19796 => conv_std_logic_vector(25, 8),
19797 => conv_std_logic_vector(25, 8),
19798 => conv_std_logic_vector(25, 8),
19799 => conv_std_logic_vector(26, 8),
19800 => conv_std_logic_vector(26, 8),
19801 => conv_std_logic_vector(26, 8),
19802 => conv_std_logic_vector(27, 8),
19803 => conv_std_logic_vector(27, 8),
19804 => conv_std_logic_vector(27, 8),
19805 => conv_std_logic_vector(27, 8),
19806 => conv_std_logic_vector(28, 8),
19807 => conv_std_logic_vector(28, 8),
19808 => conv_std_logic_vector(28, 8),
19809 => conv_std_logic_vector(29, 8),
19810 => conv_std_logic_vector(29, 8),
19811 => conv_std_logic_vector(29, 8),
19812 => conv_std_logic_vector(30, 8),
19813 => conv_std_logic_vector(30, 8),
19814 => conv_std_logic_vector(30, 8),
19815 => conv_std_logic_vector(30, 8),
19816 => conv_std_logic_vector(31, 8),
19817 => conv_std_logic_vector(31, 8),
19818 => conv_std_logic_vector(31, 8),
19819 => conv_std_logic_vector(32, 8),
19820 => conv_std_logic_vector(32, 8),
19821 => conv_std_logic_vector(32, 8),
19822 => conv_std_logic_vector(33, 8),
19823 => conv_std_logic_vector(33, 8),
19824 => conv_std_logic_vector(33, 8),
19825 => conv_std_logic_vector(33, 8),
19826 => conv_std_logic_vector(34, 8),
19827 => conv_std_logic_vector(34, 8),
19828 => conv_std_logic_vector(34, 8),
19829 => conv_std_logic_vector(35, 8),
19830 => conv_std_logic_vector(35, 8),
19831 => conv_std_logic_vector(35, 8),
19832 => conv_std_logic_vector(36, 8),
19833 => conv_std_logic_vector(36, 8),
19834 => conv_std_logic_vector(36, 8),
19835 => conv_std_logic_vector(36, 8),
19836 => conv_std_logic_vector(37, 8),
19837 => conv_std_logic_vector(37, 8),
19838 => conv_std_logic_vector(37, 8),
19839 => conv_std_logic_vector(38, 8),
19840 => conv_std_logic_vector(38, 8),
19841 => conv_std_logic_vector(38, 8),
19842 => conv_std_logic_vector(39, 8),
19843 => conv_std_logic_vector(39, 8),
19844 => conv_std_logic_vector(39, 8),
19845 => conv_std_logic_vector(40, 8),
19846 => conv_std_logic_vector(40, 8),
19847 => conv_std_logic_vector(40, 8),
19848 => conv_std_logic_vector(40, 8),
19849 => conv_std_logic_vector(41, 8),
19850 => conv_std_logic_vector(41, 8),
19851 => conv_std_logic_vector(41, 8),
19852 => conv_std_logic_vector(42, 8),
19853 => conv_std_logic_vector(42, 8),
19854 => conv_std_logic_vector(42, 8),
19855 => conv_std_logic_vector(43, 8),
19856 => conv_std_logic_vector(43, 8),
19857 => conv_std_logic_vector(43, 8),
19858 => conv_std_logic_vector(43, 8),
19859 => conv_std_logic_vector(44, 8),
19860 => conv_std_logic_vector(44, 8),
19861 => conv_std_logic_vector(44, 8),
19862 => conv_std_logic_vector(45, 8),
19863 => conv_std_logic_vector(45, 8),
19864 => conv_std_logic_vector(45, 8),
19865 => conv_std_logic_vector(46, 8),
19866 => conv_std_logic_vector(46, 8),
19867 => conv_std_logic_vector(46, 8),
19868 => conv_std_logic_vector(46, 8),
19869 => conv_std_logic_vector(47, 8),
19870 => conv_std_logic_vector(47, 8),
19871 => conv_std_logic_vector(47, 8),
19872 => conv_std_logic_vector(48, 8),
19873 => conv_std_logic_vector(48, 8),
19874 => conv_std_logic_vector(48, 8),
19875 => conv_std_logic_vector(49, 8),
19876 => conv_std_logic_vector(49, 8),
19877 => conv_std_logic_vector(49, 8),
19878 => conv_std_logic_vector(49, 8),
19879 => conv_std_logic_vector(50, 8),
19880 => conv_std_logic_vector(50, 8),
19881 => conv_std_logic_vector(50, 8),
19882 => conv_std_logic_vector(51, 8),
19883 => conv_std_logic_vector(51, 8),
19884 => conv_std_logic_vector(51, 8),
19885 => conv_std_logic_vector(52, 8),
19886 => conv_std_logic_vector(52, 8),
19887 => conv_std_logic_vector(52, 8),
19888 => conv_std_logic_vector(52, 8),
19889 => conv_std_logic_vector(53, 8),
19890 => conv_std_logic_vector(53, 8),
19891 => conv_std_logic_vector(53, 8),
19892 => conv_std_logic_vector(54, 8),
19893 => conv_std_logic_vector(54, 8),
19894 => conv_std_logic_vector(54, 8),
19895 => conv_std_logic_vector(55, 8),
19896 => conv_std_logic_vector(55, 8),
19897 => conv_std_logic_vector(55, 8),
19898 => conv_std_logic_vector(55, 8),
19899 => conv_std_logic_vector(56, 8),
19900 => conv_std_logic_vector(56, 8),
19901 => conv_std_logic_vector(56, 8),
19902 => conv_std_logic_vector(57, 8),
19903 => conv_std_logic_vector(57, 8),
19904 => conv_std_logic_vector(57, 8),
19905 => conv_std_logic_vector(58, 8),
19906 => conv_std_logic_vector(58, 8),
19907 => conv_std_logic_vector(58, 8),
19908 => conv_std_logic_vector(58, 8),
19909 => conv_std_logic_vector(59, 8),
19910 => conv_std_logic_vector(59, 8),
19911 => conv_std_logic_vector(59, 8),
19912 => conv_std_logic_vector(60, 8),
19913 => conv_std_logic_vector(60, 8),
19914 => conv_std_logic_vector(60, 8),
19915 => conv_std_logic_vector(61, 8),
19916 => conv_std_logic_vector(61, 8),
19917 => conv_std_logic_vector(61, 8),
19918 => conv_std_logic_vector(61, 8),
19919 => conv_std_logic_vector(62, 8),
19920 => conv_std_logic_vector(62, 8),
19921 => conv_std_logic_vector(62, 8),
19922 => conv_std_logic_vector(63, 8),
19923 => conv_std_logic_vector(63, 8),
19924 => conv_std_logic_vector(63, 8),
19925 => conv_std_logic_vector(64, 8),
19926 => conv_std_logic_vector(64, 8),
19927 => conv_std_logic_vector(64, 8),
19928 => conv_std_logic_vector(64, 8),
19929 => conv_std_logic_vector(65, 8),
19930 => conv_std_logic_vector(65, 8),
19931 => conv_std_logic_vector(65, 8),
19932 => conv_std_logic_vector(66, 8),
19933 => conv_std_logic_vector(66, 8),
19934 => conv_std_logic_vector(66, 8),
19935 => conv_std_logic_vector(67, 8),
19936 => conv_std_logic_vector(67, 8),
19937 => conv_std_logic_vector(67, 8),
19938 => conv_std_logic_vector(67, 8),
19939 => conv_std_logic_vector(68, 8),
19940 => conv_std_logic_vector(68, 8),
19941 => conv_std_logic_vector(68, 8),
19942 => conv_std_logic_vector(69, 8),
19943 => conv_std_logic_vector(69, 8),
19944 => conv_std_logic_vector(69, 8),
19945 => conv_std_logic_vector(70, 8),
19946 => conv_std_logic_vector(70, 8),
19947 => conv_std_logic_vector(70, 8),
19948 => conv_std_logic_vector(70, 8),
19949 => conv_std_logic_vector(71, 8),
19950 => conv_std_logic_vector(71, 8),
19951 => conv_std_logic_vector(71, 8),
19952 => conv_std_logic_vector(72, 8),
19953 => conv_std_logic_vector(72, 8),
19954 => conv_std_logic_vector(72, 8),
19955 => conv_std_logic_vector(73, 8),
19956 => conv_std_logic_vector(73, 8),
19957 => conv_std_logic_vector(73, 8),
19958 => conv_std_logic_vector(73, 8),
19959 => conv_std_logic_vector(74, 8),
19960 => conv_std_logic_vector(74, 8),
19961 => conv_std_logic_vector(74, 8),
19962 => conv_std_logic_vector(75, 8),
19963 => conv_std_logic_vector(75, 8),
19964 => conv_std_logic_vector(75, 8),
19965 => conv_std_logic_vector(76, 8),
19966 => conv_std_logic_vector(76, 8),
19967 => conv_std_logic_vector(76, 8),
19968 => conv_std_logic_vector(0, 8),
19969 => conv_std_logic_vector(0, 8),
19970 => conv_std_logic_vector(0, 8),
19971 => conv_std_logic_vector(0, 8),
19972 => conv_std_logic_vector(1, 8),
19973 => conv_std_logic_vector(1, 8),
19974 => conv_std_logic_vector(1, 8),
19975 => conv_std_logic_vector(2, 8),
19976 => conv_std_logic_vector(2, 8),
19977 => conv_std_logic_vector(2, 8),
19978 => conv_std_logic_vector(3, 8),
19979 => conv_std_logic_vector(3, 8),
19980 => conv_std_logic_vector(3, 8),
19981 => conv_std_logic_vector(3, 8),
19982 => conv_std_logic_vector(4, 8),
19983 => conv_std_logic_vector(4, 8),
19984 => conv_std_logic_vector(4, 8),
19985 => conv_std_logic_vector(5, 8),
19986 => conv_std_logic_vector(5, 8),
19987 => conv_std_logic_vector(5, 8),
19988 => conv_std_logic_vector(6, 8),
19989 => conv_std_logic_vector(6, 8),
19990 => conv_std_logic_vector(6, 8),
19991 => conv_std_logic_vector(7, 8),
19992 => conv_std_logic_vector(7, 8),
19993 => conv_std_logic_vector(7, 8),
19994 => conv_std_logic_vector(7, 8),
19995 => conv_std_logic_vector(8, 8),
19996 => conv_std_logic_vector(8, 8),
19997 => conv_std_logic_vector(8, 8),
19998 => conv_std_logic_vector(9, 8),
19999 => conv_std_logic_vector(9, 8),
20000 => conv_std_logic_vector(9, 8),
20001 => conv_std_logic_vector(10, 8),
20002 => conv_std_logic_vector(10, 8),
20003 => conv_std_logic_vector(10, 8),
20004 => conv_std_logic_vector(10, 8),
20005 => conv_std_logic_vector(11, 8),
20006 => conv_std_logic_vector(11, 8),
20007 => conv_std_logic_vector(11, 8),
20008 => conv_std_logic_vector(12, 8),
20009 => conv_std_logic_vector(12, 8),
20010 => conv_std_logic_vector(12, 8),
20011 => conv_std_logic_vector(13, 8),
20012 => conv_std_logic_vector(13, 8),
20013 => conv_std_logic_vector(13, 8),
20014 => conv_std_logic_vector(14, 8),
20015 => conv_std_logic_vector(14, 8),
20016 => conv_std_logic_vector(14, 8),
20017 => conv_std_logic_vector(14, 8),
20018 => conv_std_logic_vector(15, 8),
20019 => conv_std_logic_vector(15, 8),
20020 => conv_std_logic_vector(15, 8),
20021 => conv_std_logic_vector(16, 8),
20022 => conv_std_logic_vector(16, 8),
20023 => conv_std_logic_vector(16, 8),
20024 => conv_std_logic_vector(17, 8),
20025 => conv_std_logic_vector(17, 8),
20026 => conv_std_logic_vector(17, 8),
20027 => conv_std_logic_vector(17, 8),
20028 => conv_std_logic_vector(18, 8),
20029 => conv_std_logic_vector(18, 8),
20030 => conv_std_logic_vector(18, 8),
20031 => conv_std_logic_vector(19, 8),
20032 => conv_std_logic_vector(19, 8),
20033 => conv_std_logic_vector(19, 8),
20034 => conv_std_logic_vector(20, 8),
20035 => conv_std_logic_vector(20, 8),
20036 => conv_std_logic_vector(20, 8),
20037 => conv_std_logic_vector(21, 8),
20038 => conv_std_logic_vector(21, 8),
20039 => conv_std_logic_vector(21, 8),
20040 => conv_std_logic_vector(21, 8),
20041 => conv_std_logic_vector(22, 8),
20042 => conv_std_logic_vector(22, 8),
20043 => conv_std_logic_vector(22, 8),
20044 => conv_std_logic_vector(23, 8),
20045 => conv_std_logic_vector(23, 8),
20046 => conv_std_logic_vector(23, 8),
20047 => conv_std_logic_vector(24, 8),
20048 => conv_std_logic_vector(24, 8),
20049 => conv_std_logic_vector(24, 8),
20050 => conv_std_logic_vector(24, 8),
20051 => conv_std_logic_vector(25, 8),
20052 => conv_std_logic_vector(25, 8),
20053 => conv_std_logic_vector(25, 8),
20054 => conv_std_logic_vector(26, 8),
20055 => conv_std_logic_vector(26, 8),
20056 => conv_std_logic_vector(26, 8),
20057 => conv_std_logic_vector(27, 8),
20058 => conv_std_logic_vector(27, 8),
20059 => conv_std_logic_vector(27, 8),
20060 => conv_std_logic_vector(28, 8),
20061 => conv_std_logic_vector(28, 8),
20062 => conv_std_logic_vector(28, 8),
20063 => conv_std_logic_vector(28, 8),
20064 => conv_std_logic_vector(29, 8),
20065 => conv_std_logic_vector(29, 8),
20066 => conv_std_logic_vector(29, 8),
20067 => conv_std_logic_vector(30, 8),
20068 => conv_std_logic_vector(30, 8),
20069 => conv_std_logic_vector(30, 8),
20070 => conv_std_logic_vector(31, 8),
20071 => conv_std_logic_vector(31, 8),
20072 => conv_std_logic_vector(31, 8),
20073 => conv_std_logic_vector(31, 8),
20074 => conv_std_logic_vector(32, 8),
20075 => conv_std_logic_vector(32, 8),
20076 => conv_std_logic_vector(32, 8),
20077 => conv_std_logic_vector(33, 8),
20078 => conv_std_logic_vector(33, 8),
20079 => conv_std_logic_vector(33, 8),
20080 => conv_std_logic_vector(34, 8),
20081 => conv_std_logic_vector(34, 8),
20082 => conv_std_logic_vector(34, 8),
20083 => conv_std_logic_vector(35, 8),
20084 => conv_std_logic_vector(35, 8),
20085 => conv_std_logic_vector(35, 8),
20086 => conv_std_logic_vector(35, 8),
20087 => conv_std_logic_vector(36, 8),
20088 => conv_std_logic_vector(36, 8),
20089 => conv_std_logic_vector(36, 8),
20090 => conv_std_logic_vector(37, 8),
20091 => conv_std_logic_vector(37, 8),
20092 => conv_std_logic_vector(37, 8),
20093 => conv_std_logic_vector(38, 8),
20094 => conv_std_logic_vector(38, 8),
20095 => conv_std_logic_vector(38, 8),
20096 => conv_std_logic_vector(39, 8),
20097 => conv_std_logic_vector(39, 8),
20098 => conv_std_logic_vector(39, 8),
20099 => conv_std_logic_vector(39, 8),
20100 => conv_std_logic_vector(40, 8),
20101 => conv_std_logic_vector(40, 8),
20102 => conv_std_logic_vector(40, 8),
20103 => conv_std_logic_vector(41, 8),
20104 => conv_std_logic_vector(41, 8),
20105 => conv_std_logic_vector(41, 8),
20106 => conv_std_logic_vector(42, 8),
20107 => conv_std_logic_vector(42, 8),
20108 => conv_std_logic_vector(42, 8),
20109 => conv_std_logic_vector(42, 8),
20110 => conv_std_logic_vector(43, 8),
20111 => conv_std_logic_vector(43, 8),
20112 => conv_std_logic_vector(43, 8),
20113 => conv_std_logic_vector(44, 8),
20114 => conv_std_logic_vector(44, 8),
20115 => conv_std_logic_vector(44, 8),
20116 => conv_std_logic_vector(45, 8),
20117 => conv_std_logic_vector(45, 8),
20118 => conv_std_logic_vector(45, 8),
20119 => conv_std_logic_vector(46, 8),
20120 => conv_std_logic_vector(46, 8),
20121 => conv_std_logic_vector(46, 8),
20122 => conv_std_logic_vector(46, 8),
20123 => conv_std_logic_vector(47, 8),
20124 => conv_std_logic_vector(47, 8),
20125 => conv_std_logic_vector(47, 8),
20126 => conv_std_logic_vector(48, 8),
20127 => conv_std_logic_vector(48, 8),
20128 => conv_std_logic_vector(48, 8),
20129 => conv_std_logic_vector(49, 8),
20130 => conv_std_logic_vector(49, 8),
20131 => conv_std_logic_vector(49, 8),
20132 => conv_std_logic_vector(49, 8),
20133 => conv_std_logic_vector(50, 8),
20134 => conv_std_logic_vector(50, 8),
20135 => conv_std_logic_vector(50, 8),
20136 => conv_std_logic_vector(51, 8),
20137 => conv_std_logic_vector(51, 8),
20138 => conv_std_logic_vector(51, 8),
20139 => conv_std_logic_vector(52, 8),
20140 => conv_std_logic_vector(52, 8),
20141 => conv_std_logic_vector(52, 8),
20142 => conv_std_logic_vector(53, 8),
20143 => conv_std_logic_vector(53, 8),
20144 => conv_std_logic_vector(53, 8),
20145 => conv_std_logic_vector(53, 8),
20146 => conv_std_logic_vector(54, 8),
20147 => conv_std_logic_vector(54, 8),
20148 => conv_std_logic_vector(54, 8),
20149 => conv_std_logic_vector(55, 8),
20150 => conv_std_logic_vector(55, 8),
20151 => conv_std_logic_vector(55, 8),
20152 => conv_std_logic_vector(56, 8),
20153 => conv_std_logic_vector(56, 8),
20154 => conv_std_logic_vector(56, 8),
20155 => conv_std_logic_vector(56, 8),
20156 => conv_std_logic_vector(57, 8),
20157 => conv_std_logic_vector(57, 8),
20158 => conv_std_logic_vector(57, 8),
20159 => conv_std_logic_vector(58, 8),
20160 => conv_std_logic_vector(58, 8),
20161 => conv_std_logic_vector(58, 8),
20162 => conv_std_logic_vector(59, 8),
20163 => conv_std_logic_vector(59, 8),
20164 => conv_std_logic_vector(59, 8),
20165 => conv_std_logic_vector(60, 8),
20166 => conv_std_logic_vector(60, 8),
20167 => conv_std_logic_vector(60, 8),
20168 => conv_std_logic_vector(60, 8),
20169 => conv_std_logic_vector(61, 8),
20170 => conv_std_logic_vector(61, 8),
20171 => conv_std_logic_vector(61, 8),
20172 => conv_std_logic_vector(62, 8),
20173 => conv_std_logic_vector(62, 8),
20174 => conv_std_logic_vector(62, 8),
20175 => conv_std_logic_vector(63, 8),
20176 => conv_std_logic_vector(63, 8),
20177 => conv_std_logic_vector(63, 8),
20178 => conv_std_logic_vector(63, 8),
20179 => conv_std_logic_vector(64, 8),
20180 => conv_std_logic_vector(64, 8),
20181 => conv_std_logic_vector(64, 8),
20182 => conv_std_logic_vector(65, 8),
20183 => conv_std_logic_vector(65, 8),
20184 => conv_std_logic_vector(65, 8),
20185 => conv_std_logic_vector(66, 8),
20186 => conv_std_logic_vector(66, 8),
20187 => conv_std_logic_vector(66, 8),
20188 => conv_std_logic_vector(67, 8),
20189 => conv_std_logic_vector(67, 8),
20190 => conv_std_logic_vector(67, 8),
20191 => conv_std_logic_vector(67, 8),
20192 => conv_std_logic_vector(68, 8),
20193 => conv_std_logic_vector(68, 8),
20194 => conv_std_logic_vector(68, 8),
20195 => conv_std_logic_vector(69, 8),
20196 => conv_std_logic_vector(69, 8),
20197 => conv_std_logic_vector(69, 8),
20198 => conv_std_logic_vector(70, 8),
20199 => conv_std_logic_vector(70, 8),
20200 => conv_std_logic_vector(70, 8),
20201 => conv_std_logic_vector(70, 8),
20202 => conv_std_logic_vector(71, 8),
20203 => conv_std_logic_vector(71, 8),
20204 => conv_std_logic_vector(71, 8),
20205 => conv_std_logic_vector(72, 8),
20206 => conv_std_logic_vector(72, 8),
20207 => conv_std_logic_vector(72, 8),
20208 => conv_std_logic_vector(73, 8),
20209 => conv_std_logic_vector(73, 8),
20210 => conv_std_logic_vector(73, 8),
20211 => conv_std_logic_vector(74, 8),
20212 => conv_std_logic_vector(74, 8),
20213 => conv_std_logic_vector(74, 8),
20214 => conv_std_logic_vector(74, 8),
20215 => conv_std_logic_vector(75, 8),
20216 => conv_std_logic_vector(75, 8),
20217 => conv_std_logic_vector(75, 8),
20218 => conv_std_logic_vector(76, 8),
20219 => conv_std_logic_vector(76, 8),
20220 => conv_std_logic_vector(76, 8),
20221 => conv_std_logic_vector(77, 8),
20222 => conv_std_logic_vector(77, 8),
20223 => conv_std_logic_vector(77, 8),
20224 => conv_std_logic_vector(0, 8),
20225 => conv_std_logic_vector(0, 8),
20226 => conv_std_logic_vector(0, 8),
20227 => conv_std_logic_vector(0, 8),
20228 => conv_std_logic_vector(1, 8),
20229 => conv_std_logic_vector(1, 8),
20230 => conv_std_logic_vector(1, 8),
20231 => conv_std_logic_vector(2, 8),
20232 => conv_std_logic_vector(2, 8),
20233 => conv_std_logic_vector(2, 8),
20234 => conv_std_logic_vector(3, 8),
20235 => conv_std_logic_vector(3, 8),
20236 => conv_std_logic_vector(3, 8),
20237 => conv_std_logic_vector(4, 8),
20238 => conv_std_logic_vector(4, 8),
20239 => conv_std_logic_vector(4, 8),
20240 => conv_std_logic_vector(4, 8),
20241 => conv_std_logic_vector(5, 8),
20242 => conv_std_logic_vector(5, 8),
20243 => conv_std_logic_vector(5, 8),
20244 => conv_std_logic_vector(6, 8),
20245 => conv_std_logic_vector(6, 8),
20246 => conv_std_logic_vector(6, 8),
20247 => conv_std_logic_vector(7, 8),
20248 => conv_std_logic_vector(7, 8),
20249 => conv_std_logic_vector(7, 8),
20250 => conv_std_logic_vector(8, 8),
20251 => conv_std_logic_vector(8, 8),
20252 => conv_std_logic_vector(8, 8),
20253 => conv_std_logic_vector(8, 8),
20254 => conv_std_logic_vector(9, 8),
20255 => conv_std_logic_vector(9, 8),
20256 => conv_std_logic_vector(9, 8),
20257 => conv_std_logic_vector(10, 8),
20258 => conv_std_logic_vector(10, 8),
20259 => conv_std_logic_vector(10, 8),
20260 => conv_std_logic_vector(11, 8),
20261 => conv_std_logic_vector(11, 8),
20262 => conv_std_logic_vector(11, 8),
20263 => conv_std_logic_vector(12, 8),
20264 => conv_std_logic_vector(12, 8),
20265 => conv_std_logic_vector(12, 8),
20266 => conv_std_logic_vector(12, 8),
20267 => conv_std_logic_vector(13, 8),
20268 => conv_std_logic_vector(13, 8),
20269 => conv_std_logic_vector(13, 8),
20270 => conv_std_logic_vector(14, 8),
20271 => conv_std_logic_vector(14, 8),
20272 => conv_std_logic_vector(14, 8),
20273 => conv_std_logic_vector(15, 8),
20274 => conv_std_logic_vector(15, 8),
20275 => conv_std_logic_vector(15, 8),
20276 => conv_std_logic_vector(16, 8),
20277 => conv_std_logic_vector(16, 8),
20278 => conv_std_logic_vector(16, 8),
20279 => conv_std_logic_vector(16, 8),
20280 => conv_std_logic_vector(17, 8),
20281 => conv_std_logic_vector(17, 8),
20282 => conv_std_logic_vector(17, 8),
20283 => conv_std_logic_vector(18, 8),
20284 => conv_std_logic_vector(18, 8),
20285 => conv_std_logic_vector(18, 8),
20286 => conv_std_logic_vector(19, 8),
20287 => conv_std_logic_vector(19, 8),
20288 => conv_std_logic_vector(19, 8),
20289 => conv_std_logic_vector(20, 8),
20290 => conv_std_logic_vector(20, 8),
20291 => conv_std_logic_vector(20, 8),
20292 => conv_std_logic_vector(20, 8),
20293 => conv_std_logic_vector(21, 8),
20294 => conv_std_logic_vector(21, 8),
20295 => conv_std_logic_vector(21, 8),
20296 => conv_std_logic_vector(22, 8),
20297 => conv_std_logic_vector(22, 8),
20298 => conv_std_logic_vector(22, 8),
20299 => conv_std_logic_vector(23, 8),
20300 => conv_std_logic_vector(23, 8),
20301 => conv_std_logic_vector(23, 8),
20302 => conv_std_logic_vector(24, 8),
20303 => conv_std_logic_vector(24, 8),
20304 => conv_std_logic_vector(24, 8),
20305 => conv_std_logic_vector(24, 8),
20306 => conv_std_logic_vector(25, 8),
20307 => conv_std_logic_vector(25, 8),
20308 => conv_std_logic_vector(25, 8),
20309 => conv_std_logic_vector(26, 8),
20310 => conv_std_logic_vector(26, 8),
20311 => conv_std_logic_vector(26, 8),
20312 => conv_std_logic_vector(27, 8),
20313 => conv_std_logic_vector(27, 8),
20314 => conv_std_logic_vector(27, 8),
20315 => conv_std_logic_vector(28, 8),
20316 => conv_std_logic_vector(28, 8),
20317 => conv_std_logic_vector(28, 8),
20318 => conv_std_logic_vector(29, 8),
20319 => conv_std_logic_vector(29, 8),
20320 => conv_std_logic_vector(29, 8),
20321 => conv_std_logic_vector(29, 8),
20322 => conv_std_logic_vector(30, 8),
20323 => conv_std_logic_vector(30, 8),
20324 => conv_std_logic_vector(30, 8),
20325 => conv_std_logic_vector(31, 8),
20326 => conv_std_logic_vector(31, 8),
20327 => conv_std_logic_vector(31, 8),
20328 => conv_std_logic_vector(32, 8),
20329 => conv_std_logic_vector(32, 8),
20330 => conv_std_logic_vector(32, 8),
20331 => conv_std_logic_vector(33, 8),
20332 => conv_std_logic_vector(33, 8),
20333 => conv_std_logic_vector(33, 8),
20334 => conv_std_logic_vector(33, 8),
20335 => conv_std_logic_vector(34, 8),
20336 => conv_std_logic_vector(34, 8),
20337 => conv_std_logic_vector(34, 8),
20338 => conv_std_logic_vector(35, 8),
20339 => conv_std_logic_vector(35, 8),
20340 => conv_std_logic_vector(35, 8),
20341 => conv_std_logic_vector(36, 8),
20342 => conv_std_logic_vector(36, 8),
20343 => conv_std_logic_vector(36, 8),
20344 => conv_std_logic_vector(37, 8),
20345 => conv_std_logic_vector(37, 8),
20346 => conv_std_logic_vector(37, 8),
20347 => conv_std_logic_vector(37, 8),
20348 => conv_std_logic_vector(38, 8),
20349 => conv_std_logic_vector(38, 8),
20350 => conv_std_logic_vector(38, 8),
20351 => conv_std_logic_vector(39, 8),
20352 => conv_std_logic_vector(39, 8),
20353 => conv_std_logic_vector(39, 8),
20354 => conv_std_logic_vector(40, 8),
20355 => conv_std_logic_vector(40, 8),
20356 => conv_std_logic_vector(40, 8),
20357 => conv_std_logic_vector(41, 8),
20358 => conv_std_logic_vector(41, 8),
20359 => conv_std_logic_vector(41, 8),
20360 => conv_std_logic_vector(41, 8),
20361 => conv_std_logic_vector(42, 8),
20362 => conv_std_logic_vector(42, 8),
20363 => conv_std_logic_vector(42, 8),
20364 => conv_std_logic_vector(43, 8),
20365 => conv_std_logic_vector(43, 8),
20366 => conv_std_logic_vector(43, 8),
20367 => conv_std_logic_vector(44, 8),
20368 => conv_std_logic_vector(44, 8),
20369 => conv_std_logic_vector(44, 8),
20370 => conv_std_logic_vector(45, 8),
20371 => conv_std_logic_vector(45, 8),
20372 => conv_std_logic_vector(45, 8),
20373 => conv_std_logic_vector(45, 8),
20374 => conv_std_logic_vector(46, 8),
20375 => conv_std_logic_vector(46, 8),
20376 => conv_std_logic_vector(46, 8),
20377 => conv_std_logic_vector(47, 8),
20378 => conv_std_logic_vector(47, 8),
20379 => conv_std_logic_vector(47, 8),
20380 => conv_std_logic_vector(48, 8),
20381 => conv_std_logic_vector(48, 8),
20382 => conv_std_logic_vector(48, 8),
20383 => conv_std_logic_vector(49, 8),
20384 => conv_std_logic_vector(49, 8),
20385 => conv_std_logic_vector(49, 8),
20386 => conv_std_logic_vector(49, 8),
20387 => conv_std_logic_vector(50, 8),
20388 => conv_std_logic_vector(50, 8),
20389 => conv_std_logic_vector(50, 8),
20390 => conv_std_logic_vector(51, 8),
20391 => conv_std_logic_vector(51, 8),
20392 => conv_std_logic_vector(51, 8),
20393 => conv_std_logic_vector(52, 8),
20394 => conv_std_logic_vector(52, 8),
20395 => conv_std_logic_vector(52, 8),
20396 => conv_std_logic_vector(53, 8),
20397 => conv_std_logic_vector(53, 8),
20398 => conv_std_logic_vector(53, 8),
20399 => conv_std_logic_vector(54, 8),
20400 => conv_std_logic_vector(54, 8),
20401 => conv_std_logic_vector(54, 8),
20402 => conv_std_logic_vector(54, 8),
20403 => conv_std_logic_vector(55, 8),
20404 => conv_std_logic_vector(55, 8),
20405 => conv_std_logic_vector(55, 8),
20406 => conv_std_logic_vector(56, 8),
20407 => conv_std_logic_vector(56, 8),
20408 => conv_std_logic_vector(56, 8),
20409 => conv_std_logic_vector(57, 8),
20410 => conv_std_logic_vector(57, 8),
20411 => conv_std_logic_vector(57, 8),
20412 => conv_std_logic_vector(58, 8),
20413 => conv_std_logic_vector(58, 8),
20414 => conv_std_logic_vector(58, 8),
20415 => conv_std_logic_vector(58, 8),
20416 => conv_std_logic_vector(59, 8),
20417 => conv_std_logic_vector(59, 8),
20418 => conv_std_logic_vector(59, 8),
20419 => conv_std_logic_vector(60, 8),
20420 => conv_std_logic_vector(60, 8),
20421 => conv_std_logic_vector(60, 8),
20422 => conv_std_logic_vector(61, 8),
20423 => conv_std_logic_vector(61, 8),
20424 => conv_std_logic_vector(61, 8),
20425 => conv_std_logic_vector(62, 8),
20426 => conv_std_logic_vector(62, 8),
20427 => conv_std_logic_vector(62, 8),
20428 => conv_std_logic_vector(62, 8),
20429 => conv_std_logic_vector(63, 8),
20430 => conv_std_logic_vector(63, 8),
20431 => conv_std_logic_vector(63, 8),
20432 => conv_std_logic_vector(64, 8),
20433 => conv_std_logic_vector(64, 8),
20434 => conv_std_logic_vector(64, 8),
20435 => conv_std_logic_vector(65, 8),
20436 => conv_std_logic_vector(65, 8),
20437 => conv_std_logic_vector(65, 8),
20438 => conv_std_logic_vector(66, 8),
20439 => conv_std_logic_vector(66, 8),
20440 => conv_std_logic_vector(66, 8),
20441 => conv_std_logic_vector(66, 8),
20442 => conv_std_logic_vector(67, 8),
20443 => conv_std_logic_vector(67, 8),
20444 => conv_std_logic_vector(67, 8),
20445 => conv_std_logic_vector(68, 8),
20446 => conv_std_logic_vector(68, 8),
20447 => conv_std_logic_vector(68, 8),
20448 => conv_std_logic_vector(69, 8),
20449 => conv_std_logic_vector(69, 8),
20450 => conv_std_logic_vector(69, 8),
20451 => conv_std_logic_vector(70, 8),
20452 => conv_std_logic_vector(70, 8),
20453 => conv_std_logic_vector(70, 8),
20454 => conv_std_logic_vector(70, 8),
20455 => conv_std_logic_vector(71, 8),
20456 => conv_std_logic_vector(71, 8),
20457 => conv_std_logic_vector(71, 8),
20458 => conv_std_logic_vector(72, 8),
20459 => conv_std_logic_vector(72, 8),
20460 => conv_std_logic_vector(72, 8),
20461 => conv_std_logic_vector(73, 8),
20462 => conv_std_logic_vector(73, 8),
20463 => conv_std_logic_vector(73, 8),
20464 => conv_std_logic_vector(74, 8),
20465 => conv_std_logic_vector(74, 8),
20466 => conv_std_logic_vector(74, 8),
20467 => conv_std_logic_vector(74, 8),
20468 => conv_std_logic_vector(75, 8),
20469 => conv_std_logic_vector(75, 8),
20470 => conv_std_logic_vector(75, 8),
20471 => conv_std_logic_vector(76, 8),
20472 => conv_std_logic_vector(76, 8),
20473 => conv_std_logic_vector(76, 8),
20474 => conv_std_logic_vector(77, 8),
20475 => conv_std_logic_vector(77, 8),
20476 => conv_std_logic_vector(77, 8),
20477 => conv_std_logic_vector(78, 8),
20478 => conv_std_logic_vector(78, 8),
20479 => conv_std_logic_vector(78, 8),
20480 => conv_std_logic_vector(0, 8),
20481 => conv_std_logic_vector(0, 8),
20482 => conv_std_logic_vector(0, 8),
20483 => conv_std_logic_vector(0, 8),
20484 => conv_std_logic_vector(1, 8),
20485 => conv_std_logic_vector(1, 8),
20486 => conv_std_logic_vector(1, 8),
20487 => conv_std_logic_vector(2, 8),
20488 => conv_std_logic_vector(2, 8),
20489 => conv_std_logic_vector(2, 8),
20490 => conv_std_logic_vector(3, 8),
20491 => conv_std_logic_vector(3, 8),
20492 => conv_std_logic_vector(3, 8),
20493 => conv_std_logic_vector(4, 8),
20494 => conv_std_logic_vector(4, 8),
20495 => conv_std_logic_vector(4, 8),
20496 => conv_std_logic_vector(5, 8),
20497 => conv_std_logic_vector(5, 8),
20498 => conv_std_logic_vector(5, 8),
20499 => conv_std_logic_vector(5, 8),
20500 => conv_std_logic_vector(6, 8),
20501 => conv_std_logic_vector(6, 8),
20502 => conv_std_logic_vector(6, 8),
20503 => conv_std_logic_vector(7, 8),
20504 => conv_std_logic_vector(7, 8),
20505 => conv_std_logic_vector(7, 8),
20506 => conv_std_logic_vector(8, 8),
20507 => conv_std_logic_vector(8, 8),
20508 => conv_std_logic_vector(8, 8),
20509 => conv_std_logic_vector(9, 8),
20510 => conv_std_logic_vector(9, 8),
20511 => conv_std_logic_vector(9, 8),
20512 => conv_std_logic_vector(10, 8),
20513 => conv_std_logic_vector(10, 8),
20514 => conv_std_logic_vector(10, 8),
20515 => conv_std_logic_vector(10, 8),
20516 => conv_std_logic_vector(11, 8),
20517 => conv_std_logic_vector(11, 8),
20518 => conv_std_logic_vector(11, 8),
20519 => conv_std_logic_vector(12, 8),
20520 => conv_std_logic_vector(12, 8),
20521 => conv_std_logic_vector(12, 8),
20522 => conv_std_logic_vector(13, 8),
20523 => conv_std_logic_vector(13, 8),
20524 => conv_std_logic_vector(13, 8),
20525 => conv_std_logic_vector(14, 8),
20526 => conv_std_logic_vector(14, 8),
20527 => conv_std_logic_vector(14, 8),
20528 => conv_std_logic_vector(15, 8),
20529 => conv_std_logic_vector(15, 8),
20530 => conv_std_logic_vector(15, 8),
20531 => conv_std_logic_vector(15, 8),
20532 => conv_std_logic_vector(16, 8),
20533 => conv_std_logic_vector(16, 8),
20534 => conv_std_logic_vector(16, 8),
20535 => conv_std_logic_vector(17, 8),
20536 => conv_std_logic_vector(17, 8),
20537 => conv_std_logic_vector(17, 8),
20538 => conv_std_logic_vector(18, 8),
20539 => conv_std_logic_vector(18, 8),
20540 => conv_std_logic_vector(18, 8),
20541 => conv_std_logic_vector(19, 8),
20542 => conv_std_logic_vector(19, 8),
20543 => conv_std_logic_vector(19, 8),
20544 => conv_std_logic_vector(20, 8),
20545 => conv_std_logic_vector(20, 8),
20546 => conv_std_logic_vector(20, 8),
20547 => conv_std_logic_vector(20, 8),
20548 => conv_std_logic_vector(21, 8),
20549 => conv_std_logic_vector(21, 8),
20550 => conv_std_logic_vector(21, 8),
20551 => conv_std_logic_vector(22, 8),
20552 => conv_std_logic_vector(22, 8),
20553 => conv_std_logic_vector(22, 8),
20554 => conv_std_logic_vector(23, 8),
20555 => conv_std_logic_vector(23, 8),
20556 => conv_std_logic_vector(23, 8),
20557 => conv_std_logic_vector(24, 8),
20558 => conv_std_logic_vector(24, 8),
20559 => conv_std_logic_vector(24, 8),
20560 => conv_std_logic_vector(25, 8),
20561 => conv_std_logic_vector(25, 8),
20562 => conv_std_logic_vector(25, 8),
20563 => conv_std_logic_vector(25, 8),
20564 => conv_std_logic_vector(26, 8),
20565 => conv_std_logic_vector(26, 8),
20566 => conv_std_logic_vector(26, 8),
20567 => conv_std_logic_vector(27, 8),
20568 => conv_std_logic_vector(27, 8),
20569 => conv_std_logic_vector(27, 8),
20570 => conv_std_logic_vector(28, 8),
20571 => conv_std_logic_vector(28, 8),
20572 => conv_std_logic_vector(28, 8),
20573 => conv_std_logic_vector(29, 8),
20574 => conv_std_logic_vector(29, 8),
20575 => conv_std_logic_vector(29, 8),
20576 => conv_std_logic_vector(30, 8),
20577 => conv_std_logic_vector(30, 8),
20578 => conv_std_logic_vector(30, 8),
20579 => conv_std_logic_vector(30, 8),
20580 => conv_std_logic_vector(31, 8),
20581 => conv_std_logic_vector(31, 8),
20582 => conv_std_logic_vector(31, 8),
20583 => conv_std_logic_vector(32, 8),
20584 => conv_std_logic_vector(32, 8),
20585 => conv_std_logic_vector(32, 8),
20586 => conv_std_logic_vector(33, 8),
20587 => conv_std_logic_vector(33, 8),
20588 => conv_std_logic_vector(33, 8),
20589 => conv_std_logic_vector(34, 8),
20590 => conv_std_logic_vector(34, 8),
20591 => conv_std_logic_vector(34, 8),
20592 => conv_std_logic_vector(35, 8),
20593 => conv_std_logic_vector(35, 8),
20594 => conv_std_logic_vector(35, 8),
20595 => conv_std_logic_vector(35, 8),
20596 => conv_std_logic_vector(36, 8),
20597 => conv_std_logic_vector(36, 8),
20598 => conv_std_logic_vector(36, 8),
20599 => conv_std_logic_vector(37, 8),
20600 => conv_std_logic_vector(37, 8),
20601 => conv_std_logic_vector(37, 8),
20602 => conv_std_logic_vector(38, 8),
20603 => conv_std_logic_vector(38, 8),
20604 => conv_std_logic_vector(38, 8),
20605 => conv_std_logic_vector(39, 8),
20606 => conv_std_logic_vector(39, 8),
20607 => conv_std_logic_vector(39, 8),
20608 => conv_std_logic_vector(40, 8),
20609 => conv_std_logic_vector(40, 8),
20610 => conv_std_logic_vector(40, 8),
20611 => conv_std_logic_vector(40, 8),
20612 => conv_std_logic_vector(41, 8),
20613 => conv_std_logic_vector(41, 8),
20614 => conv_std_logic_vector(41, 8),
20615 => conv_std_logic_vector(42, 8),
20616 => conv_std_logic_vector(42, 8),
20617 => conv_std_logic_vector(42, 8),
20618 => conv_std_logic_vector(43, 8),
20619 => conv_std_logic_vector(43, 8),
20620 => conv_std_logic_vector(43, 8),
20621 => conv_std_logic_vector(44, 8),
20622 => conv_std_logic_vector(44, 8),
20623 => conv_std_logic_vector(44, 8),
20624 => conv_std_logic_vector(45, 8),
20625 => conv_std_logic_vector(45, 8),
20626 => conv_std_logic_vector(45, 8),
20627 => conv_std_logic_vector(45, 8),
20628 => conv_std_logic_vector(46, 8),
20629 => conv_std_logic_vector(46, 8),
20630 => conv_std_logic_vector(46, 8),
20631 => conv_std_logic_vector(47, 8),
20632 => conv_std_logic_vector(47, 8),
20633 => conv_std_logic_vector(47, 8),
20634 => conv_std_logic_vector(48, 8),
20635 => conv_std_logic_vector(48, 8),
20636 => conv_std_logic_vector(48, 8),
20637 => conv_std_logic_vector(49, 8),
20638 => conv_std_logic_vector(49, 8),
20639 => conv_std_logic_vector(49, 8),
20640 => conv_std_logic_vector(50, 8),
20641 => conv_std_logic_vector(50, 8),
20642 => conv_std_logic_vector(50, 8),
20643 => conv_std_logic_vector(50, 8),
20644 => conv_std_logic_vector(51, 8),
20645 => conv_std_logic_vector(51, 8),
20646 => conv_std_logic_vector(51, 8),
20647 => conv_std_logic_vector(52, 8),
20648 => conv_std_logic_vector(52, 8),
20649 => conv_std_logic_vector(52, 8),
20650 => conv_std_logic_vector(53, 8),
20651 => conv_std_logic_vector(53, 8),
20652 => conv_std_logic_vector(53, 8),
20653 => conv_std_logic_vector(54, 8),
20654 => conv_std_logic_vector(54, 8),
20655 => conv_std_logic_vector(54, 8),
20656 => conv_std_logic_vector(55, 8),
20657 => conv_std_logic_vector(55, 8),
20658 => conv_std_logic_vector(55, 8),
20659 => conv_std_logic_vector(55, 8),
20660 => conv_std_logic_vector(56, 8),
20661 => conv_std_logic_vector(56, 8),
20662 => conv_std_logic_vector(56, 8),
20663 => conv_std_logic_vector(57, 8),
20664 => conv_std_logic_vector(57, 8),
20665 => conv_std_logic_vector(57, 8),
20666 => conv_std_logic_vector(58, 8),
20667 => conv_std_logic_vector(58, 8),
20668 => conv_std_logic_vector(58, 8),
20669 => conv_std_logic_vector(59, 8),
20670 => conv_std_logic_vector(59, 8),
20671 => conv_std_logic_vector(59, 8),
20672 => conv_std_logic_vector(60, 8),
20673 => conv_std_logic_vector(60, 8),
20674 => conv_std_logic_vector(60, 8),
20675 => conv_std_logic_vector(60, 8),
20676 => conv_std_logic_vector(61, 8),
20677 => conv_std_logic_vector(61, 8),
20678 => conv_std_logic_vector(61, 8),
20679 => conv_std_logic_vector(62, 8),
20680 => conv_std_logic_vector(62, 8),
20681 => conv_std_logic_vector(62, 8),
20682 => conv_std_logic_vector(63, 8),
20683 => conv_std_logic_vector(63, 8),
20684 => conv_std_logic_vector(63, 8),
20685 => conv_std_logic_vector(64, 8),
20686 => conv_std_logic_vector(64, 8),
20687 => conv_std_logic_vector(64, 8),
20688 => conv_std_logic_vector(65, 8),
20689 => conv_std_logic_vector(65, 8),
20690 => conv_std_logic_vector(65, 8),
20691 => conv_std_logic_vector(65, 8),
20692 => conv_std_logic_vector(66, 8),
20693 => conv_std_logic_vector(66, 8),
20694 => conv_std_logic_vector(66, 8),
20695 => conv_std_logic_vector(67, 8),
20696 => conv_std_logic_vector(67, 8),
20697 => conv_std_logic_vector(67, 8),
20698 => conv_std_logic_vector(68, 8),
20699 => conv_std_logic_vector(68, 8),
20700 => conv_std_logic_vector(68, 8),
20701 => conv_std_logic_vector(69, 8),
20702 => conv_std_logic_vector(69, 8),
20703 => conv_std_logic_vector(69, 8),
20704 => conv_std_logic_vector(70, 8),
20705 => conv_std_logic_vector(70, 8),
20706 => conv_std_logic_vector(70, 8),
20707 => conv_std_logic_vector(70, 8),
20708 => conv_std_logic_vector(71, 8),
20709 => conv_std_logic_vector(71, 8),
20710 => conv_std_logic_vector(71, 8),
20711 => conv_std_logic_vector(72, 8),
20712 => conv_std_logic_vector(72, 8),
20713 => conv_std_logic_vector(72, 8),
20714 => conv_std_logic_vector(73, 8),
20715 => conv_std_logic_vector(73, 8),
20716 => conv_std_logic_vector(73, 8),
20717 => conv_std_logic_vector(74, 8),
20718 => conv_std_logic_vector(74, 8),
20719 => conv_std_logic_vector(74, 8),
20720 => conv_std_logic_vector(75, 8),
20721 => conv_std_logic_vector(75, 8),
20722 => conv_std_logic_vector(75, 8),
20723 => conv_std_logic_vector(75, 8),
20724 => conv_std_logic_vector(76, 8),
20725 => conv_std_logic_vector(76, 8),
20726 => conv_std_logic_vector(76, 8),
20727 => conv_std_logic_vector(77, 8),
20728 => conv_std_logic_vector(77, 8),
20729 => conv_std_logic_vector(77, 8),
20730 => conv_std_logic_vector(78, 8),
20731 => conv_std_logic_vector(78, 8),
20732 => conv_std_logic_vector(78, 8),
20733 => conv_std_logic_vector(79, 8),
20734 => conv_std_logic_vector(79, 8),
20735 => conv_std_logic_vector(79, 8),
20736 => conv_std_logic_vector(0, 8),
20737 => conv_std_logic_vector(0, 8),
20738 => conv_std_logic_vector(0, 8),
20739 => conv_std_logic_vector(0, 8),
20740 => conv_std_logic_vector(1, 8),
20741 => conv_std_logic_vector(1, 8),
20742 => conv_std_logic_vector(1, 8),
20743 => conv_std_logic_vector(2, 8),
20744 => conv_std_logic_vector(2, 8),
20745 => conv_std_logic_vector(2, 8),
20746 => conv_std_logic_vector(3, 8),
20747 => conv_std_logic_vector(3, 8),
20748 => conv_std_logic_vector(3, 8),
20749 => conv_std_logic_vector(4, 8),
20750 => conv_std_logic_vector(4, 8),
20751 => conv_std_logic_vector(4, 8),
20752 => conv_std_logic_vector(5, 8),
20753 => conv_std_logic_vector(5, 8),
20754 => conv_std_logic_vector(5, 8),
20755 => conv_std_logic_vector(6, 8),
20756 => conv_std_logic_vector(6, 8),
20757 => conv_std_logic_vector(6, 8),
20758 => conv_std_logic_vector(6, 8),
20759 => conv_std_logic_vector(7, 8),
20760 => conv_std_logic_vector(7, 8),
20761 => conv_std_logic_vector(7, 8),
20762 => conv_std_logic_vector(8, 8),
20763 => conv_std_logic_vector(8, 8),
20764 => conv_std_logic_vector(8, 8),
20765 => conv_std_logic_vector(9, 8),
20766 => conv_std_logic_vector(9, 8),
20767 => conv_std_logic_vector(9, 8),
20768 => conv_std_logic_vector(10, 8),
20769 => conv_std_logic_vector(10, 8),
20770 => conv_std_logic_vector(10, 8),
20771 => conv_std_logic_vector(11, 8),
20772 => conv_std_logic_vector(11, 8),
20773 => conv_std_logic_vector(11, 8),
20774 => conv_std_logic_vector(12, 8),
20775 => conv_std_logic_vector(12, 8),
20776 => conv_std_logic_vector(12, 8),
20777 => conv_std_logic_vector(12, 8),
20778 => conv_std_logic_vector(13, 8),
20779 => conv_std_logic_vector(13, 8),
20780 => conv_std_logic_vector(13, 8),
20781 => conv_std_logic_vector(14, 8),
20782 => conv_std_logic_vector(14, 8),
20783 => conv_std_logic_vector(14, 8),
20784 => conv_std_logic_vector(15, 8),
20785 => conv_std_logic_vector(15, 8),
20786 => conv_std_logic_vector(15, 8),
20787 => conv_std_logic_vector(16, 8),
20788 => conv_std_logic_vector(16, 8),
20789 => conv_std_logic_vector(16, 8),
20790 => conv_std_logic_vector(17, 8),
20791 => conv_std_logic_vector(17, 8),
20792 => conv_std_logic_vector(17, 8),
20793 => conv_std_logic_vector(18, 8),
20794 => conv_std_logic_vector(18, 8),
20795 => conv_std_logic_vector(18, 8),
20796 => conv_std_logic_vector(18, 8),
20797 => conv_std_logic_vector(19, 8),
20798 => conv_std_logic_vector(19, 8),
20799 => conv_std_logic_vector(19, 8),
20800 => conv_std_logic_vector(20, 8),
20801 => conv_std_logic_vector(20, 8),
20802 => conv_std_logic_vector(20, 8),
20803 => conv_std_logic_vector(21, 8),
20804 => conv_std_logic_vector(21, 8),
20805 => conv_std_logic_vector(21, 8),
20806 => conv_std_logic_vector(22, 8),
20807 => conv_std_logic_vector(22, 8),
20808 => conv_std_logic_vector(22, 8),
20809 => conv_std_logic_vector(23, 8),
20810 => conv_std_logic_vector(23, 8),
20811 => conv_std_logic_vector(23, 8),
20812 => conv_std_logic_vector(24, 8),
20813 => conv_std_logic_vector(24, 8),
20814 => conv_std_logic_vector(24, 8),
20815 => conv_std_logic_vector(24, 8),
20816 => conv_std_logic_vector(25, 8),
20817 => conv_std_logic_vector(25, 8),
20818 => conv_std_logic_vector(25, 8),
20819 => conv_std_logic_vector(26, 8),
20820 => conv_std_logic_vector(26, 8),
20821 => conv_std_logic_vector(26, 8),
20822 => conv_std_logic_vector(27, 8),
20823 => conv_std_logic_vector(27, 8),
20824 => conv_std_logic_vector(27, 8),
20825 => conv_std_logic_vector(28, 8),
20826 => conv_std_logic_vector(28, 8),
20827 => conv_std_logic_vector(28, 8),
20828 => conv_std_logic_vector(29, 8),
20829 => conv_std_logic_vector(29, 8),
20830 => conv_std_logic_vector(29, 8),
20831 => conv_std_logic_vector(30, 8),
20832 => conv_std_logic_vector(30, 8),
20833 => conv_std_logic_vector(30, 8),
20834 => conv_std_logic_vector(31, 8),
20835 => conv_std_logic_vector(31, 8),
20836 => conv_std_logic_vector(31, 8),
20837 => conv_std_logic_vector(31, 8),
20838 => conv_std_logic_vector(32, 8),
20839 => conv_std_logic_vector(32, 8),
20840 => conv_std_logic_vector(32, 8),
20841 => conv_std_logic_vector(33, 8),
20842 => conv_std_logic_vector(33, 8),
20843 => conv_std_logic_vector(33, 8),
20844 => conv_std_logic_vector(34, 8),
20845 => conv_std_logic_vector(34, 8),
20846 => conv_std_logic_vector(34, 8),
20847 => conv_std_logic_vector(35, 8),
20848 => conv_std_logic_vector(35, 8),
20849 => conv_std_logic_vector(35, 8),
20850 => conv_std_logic_vector(36, 8),
20851 => conv_std_logic_vector(36, 8),
20852 => conv_std_logic_vector(36, 8),
20853 => conv_std_logic_vector(37, 8),
20854 => conv_std_logic_vector(37, 8),
20855 => conv_std_logic_vector(37, 8),
20856 => conv_std_logic_vector(37, 8),
20857 => conv_std_logic_vector(38, 8),
20858 => conv_std_logic_vector(38, 8),
20859 => conv_std_logic_vector(38, 8),
20860 => conv_std_logic_vector(39, 8),
20861 => conv_std_logic_vector(39, 8),
20862 => conv_std_logic_vector(39, 8),
20863 => conv_std_logic_vector(40, 8),
20864 => conv_std_logic_vector(40, 8),
20865 => conv_std_logic_vector(40, 8),
20866 => conv_std_logic_vector(41, 8),
20867 => conv_std_logic_vector(41, 8),
20868 => conv_std_logic_vector(41, 8),
20869 => conv_std_logic_vector(42, 8),
20870 => conv_std_logic_vector(42, 8),
20871 => conv_std_logic_vector(42, 8),
20872 => conv_std_logic_vector(43, 8),
20873 => conv_std_logic_vector(43, 8),
20874 => conv_std_logic_vector(43, 8),
20875 => conv_std_logic_vector(43, 8),
20876 => conv_std_logic_vector(44, 8),
20877 => conv_std_logic_vector(44, 8),
20878 => conv_std_logic_vector(44, 8),
20879 => conv_std_logic_vector(45, 8),
20880 => conv_std_logic_vector(45, 8),
20881 => conv_std_logic_vector(45, 8),
20882 => conv_std_logic_vector(46, 8),
20883 => conv_std_logic_vector(46, 8),
20884 => conv_std_logic_vector(46, 8),
20885 => conv_std_logic_vector(47, 8),
20886 => conv_std_logic_vector(47, 8),
20887 => conv_std_logic_vector(47, 8),
20888 => conv_std_logic_vector(48, 8),
20889 => conv_std_logic_vector(48, 8),
20890 => conv_std_logic_vector(48, 8),
20891 => conv_std_logic_vector(49, 8),
20892 => conv_std_logic_vector(49, 8),
20893 => conv_std_logic_vector(49, 8),
20894 => conv_std_logic_vector(49, 8),
20895 => conv_std_logic_vector(50, 8),
20896 => conv_std_logic_vector(50, 8),
20897 => conv_std_logic_vector(50, 8),
20898 => conv_std_logic_vector(51, 8),
20899 => conv_std_logic_vector(51, 8),
20900 => conv_std_logic_vector(51, 8),
20901 => conv_std_logic_vector(52, 8),
20902 => conv_std_logic_vector(52, 8),
20903 => conv_std_logic_vector(52, 8),
20904 => conv_std_logic_vector(53, 8),
20905 => conv_std_logic_vector(53, 8),
20906 => conv_std_logic_vector(53, 8),
20907 => conv_std_logic_vector(54, 8),
20908 => conv_std_logic_vector(54, 8),
20909 => conv_std_logic_vector(54, 8),
20910 => conv_std_logic_vector(55, 8),
20911 => conv_std_logic_vector(55, 8),
20912 => conv_std_logic_vector(55, 8),
20913 => conv_std_logic_vector(56, 8),
20914 => conv_std_logic_vector(56, 8),
20915 => conv_std_logic_vector(56, 8),
20916 => conv_std_logic_vector(56, 8),
20917 => conv_std_logic_vector(57, 8),
20918 => conv_std_logic_vector(57, 8),
20919 => conv_std_logic_vector(57, 8),
20920 => conv_std_logic_vector(58, 8),
20921 => conv_std_logic_vector(58, 8),
20922 => conv_std_logic_vector(58, 8),
20923 => conv_std_logic_vector(59, 8),
20924 => conv_std_logic_vector(59, 8),
20925 => conv_std_logic_vector(59, 8),
20926 => conv_std_logic_vector(60, 8),
20927 => conv_std_logic_vector(60, 8),
20928 => conv_std_logic_vector(60, 8),
20929 => conv_std_logic_vector(61, 8),
20930 => conv_std_logic_vector(61, 8),
20931 => conv_std_logic_vector(61, 8),
20932 => conv_std_logic_vector(62, 8),
20933 => conv_std_logic_vector(62, 8),
20934 => conv_std_logic_vector(62, 8),
20935 => conv_std_logic_vector(62, 8),
20936 => conv_std_logic_vector(63, 8),
20937 => conv_std_logic_vector(63, 8),
20938 => conv_std_logic_vector(63, 8),
20939 => conv_std_logic_vector(64, 8),
20940 => conv_std_logic_vector(64, 8),
20941 => conv_std_logic_vector(64, 8),
20942 => conv_std_logic_vector(65, 8),
20943 => conv_std_logic_vector(65, 8),
20944 => conv_std_logic_vector(65, 8),
20945 => conv_std_logic_vector(66, 8),
20946 => conv_std_logic_vector(66, 8),
20947 => conv_std_logic_vector(66, 8),
20948 => conv_std_logic_vector(67, 8),
20949 => conv_std_logic_vector(67, 8),
20950 => conv_std_logic_vector(67, 8),
20951 => conv_std_logic_vector(68, 8),
20952 => conv_std_logic_vector(68, 8),
20953 => conv_std_logic_vector(68, 8),
20954 => conv_std_logic_vector(68, 8),
20955 => conv_std_logic_vector(69, 8),
20956 => conv_std_logic_vector(69, 8),
20957 => conv_std_logic_vector(69, 8),
20958 => conv_std_logic_vector(70, 8),
20959 => conv_std_logic_vector(70, 8),
20960 => conv_std_logic_vector(70, 8),
20961 => conv_std_logic_vector(71, 8),
20962 => conv_std_logic_vector(71, 8),
20963 => conv_std_logic_vector(71, 8),
20964 => conv_std_logic_vector(72, 8),
20965 => conv_std_logic_vector(72, 8),
20966 => conv_std_logic_vector(72, 8),
20967 => conv_std_logic_vector(73, 8),
20968 => conv_std_logic_vector(73, 8),
20969 => conv_std_logic_vector(73, 8),
20970 => conv_std_logic_vector(74, 8),
20971 => conv_std_logic_vector(74, 8),
20972 => conv_std_logic_vector(74, 8),
20973 => conv_std_logic_vector(74, 8),
20974 => conv_std_logic_vector(75, 8),
20975 => conv_std_logic_vector(75, 8),
20976 => conv_std_logic_vector(75, 8),
20977 => conv_std_logic_vector(76, 8),
20978 => conv_std_logic_vector(76, 8),
20979 => conv_std_logic_vector(76, 8),
20980 => conv_std_logic_vector(77, 8),
20981 => conv_std_logic_vector(77, 8),
20982 => conv_std_logic_vector(77, 8),
20983 => conv_std_logic_vector(78, 8),
20984 => conv_std_logic_vector(78, 8),
20985 => conv_std_logic_vector(78, 8),
20986 => conv_std_logic_vector(79, 8),
20987 => conv_std_logic_vector(79, 8),
20988 => conv_std_logic_vector(79, 8),
20989 => conv_std_logic_vector(80, 8),
20990 => conv_std_logic_vector(80, 8),
20991 => conv_std_logic_vector(80, 8),
20992 => conv_std_logic_vector(0, 8),
20993 => conv_std_logic_vector(0, 8),
20994 => conv_std_logic_vector(0, 8),
20995 => conv_std_logic_vector(0, 8),
20996 => conv_std_logic_vector(1, 8),
20997 => conv_std_logic_vector(1, 8),
20998 => conv_std_logic_vector(1, 8),
20999 => conv_std_logic_vector(2, 8),
21000 => conv_std_logic_vector(2, 8),
21001 => conv_std_logic_vector(2, 8),
21002 => conv_std_logic_vector(3, 8),
21003 => conv_std_logic_vector(3, 8),
21004 => conv_std_logic_vector(3, 8),
21005 => conv_std_logic_vector(4, 8),
21006 => conv_std_logic_vector(4, 8),
21007 => conv_std_logic_vector(4, 8),
21008 => conv_std_logic_vector(5, 8),
21009 => conv_std_logic_vector(5, 8),
21010 => conv_std_logic_vector(5, 8),
21011 => conv_std_logic_vector(6, 8),
21012 => conv_std_logic_vector(6, 8),
21013 => conv_std_logic_vector(6, 8),
21014 => conv_std_logic_vector(7, 8),
21015 => conv_std_logic_vector(7, 8),
21016 => conv_std_logic_vector(7, 8),
21017 => conv_std_logic_vector(8, 8),
21018 => conv_std_logic_vector(8, 8),
21019 => conv_std_logic_vector(8, 8),
21020 => conv_std_logic_vector(8, 8),
21021 => conv_std_logic_vector(9, 8),
21022 => conv_std_logic_vector(9, 8),
21023 => conv_std_logic_vector(9, 8),
21024 => conv_std_logic_vector(10, 8),
21025 => conv_std_logic_vector(10, 8),
21026 => conv_std_logic_vector(10, 8),
21027 => conv_std_logic_vector(11, 8),
21028 => conv_std_logic_vector(11, 8),
21029 => conv_std_logic_vector(11, 8),
21030 => conv_std_logic_vector(12, 8),
21031 => conv_std_logic_vector(12, 8),
21032 => conv_std_logic_vector(12, 8),
21033 => conv_std_logic_vector(13, 8),
21034 => conv_std_logic_vector(13, 8),
21035 => conv_std_logic_vector(13, 8),
21036 => conv_std_logic_vector(14, 8),
21037 => conv_std_logic_vector(14, 8),
21038 => conv_std_logic_vector(14, 8),
21039 => conv_std_logic_vector(15, 8),
21040 => conv_std_logic_vector(15, 8),
21041 => conv_std_logic_vector(15, 8),
21042 => conv_std_logic_vector(16, 8),
21043 => conv_std_logic_vector(16, 8),
21044 => conv_std_logic_vector(16, 8),
21045 => conv_std_logic_vector(16, 8),
21046 => conv_std_logic_vector(17, 8),
21047 => conv_std_logic_vector(17, 8),
21048 => conv_std_logic_vector(17, 8),
21049 => conv_std_logic_vector(18, 8),
21050 => conv_std_logic_vector(18, 8),
21051 => conv_std_logic_vector(18, 8),
21052 => conv_std_logic_vector(19, 8),
21053 => conv_std_logic_vector(19, 8),
21054 => conv_std_logic_vector(19, 8),
21055 => conv_std_logic_vector(20, 8),
21056 => conv_std_logic_vector(20, 8),
21057 => conv_std_logic_vector(20, 8),
21058 => conv_std_logic_vector(21, 8),
21059 => conv_std_logic_vector(21, 8),
21060 => conv_std_logic_vector(21, 8),
21061 => conv_std_logic_vector(22, 8),
21062 => conv_std_logic_vector(22, 8),
21063 => conv_std_logic_vector(22, 8),
21064 => conv_std_logic_vector(23, 8),
21065 => conv_std_logic_vector(23, 8),
21066 => conv_std_logic_vector(23, 8),
21067 => conv_std_logic_vector(24, 8),
21068 => conv_std_logic_vector(24, 8),
21069 => conv_std_logic_vector(24, 8),
21070 => conv_std_logic_vector(24, 8),
21071 => conv_std_logic_vector(25, 8),
21072 => conv_std_logic_vector(25, 8),
21073 => conv_std_logic_vector(25, 8),
21074 => conv_std_logic_vector(26, 8),
21075 => conv_std_logic_vector(26, 8),
21076 => conv_std_logic_vector(26, 8),
21077 => conv_std_logic_vector(27, 8),
21078 => conv_std_logic_vector(27, 8),
21079 => conv_std_logic_vector(27, 8),
21080 => conv_std_logic_vector(28, 8),
21081 => conv_std_logic_vector(28, 8),
21082 => conv_std_logic_vector(28, 8),
21083 => conv_std_logic_vector(29, 8),
21084 => conv_std_logic_vector(29, 8),
21085 => conv_std_logic_vector(29, 8),
21086 => conv_std_logic_vector(30, 8),
21087 => conv_std_logic_vector(30, 8),
21088 => conv_std_logic_vector(30, 8),
21089 => conv_std_logic_vector(31, 8),
21090 => conv_std_logic_vector(31, 8),
21091 => conv_std_logic_vector(31, 8),
21092 => conv_std_logic_vector(32, 8),
21093 => conv_std_logic_vector(32, 8),
21094 => conv_std_logic_vector(32, 8),
21095 => conv_std_logic_vector(32, 8),
21096 => conv_std_logic_vector(33, 8),
21097 => conv_std_logic_vector(33, 8),
21098 => conv_std_logic_vector(33, 8),
21099 => conv_std_logic_vector(34, 8),
21100 => conv_std_logic_vector(34, 8),
21101 => conv_std_logic_vector(34, 8),
21102 => conv_std_logic_vector(35, 8),
21103 => conv_std_logic_vector(35, 8),
21104 => conv_std_logic_vector(35, 8),
21105 => conv_std_logic_vector(36, 8),
21106 => conv_std_logic_vector(36, 8),
21107 => conv_std_logic_vector(36, 8),
21108 => conv_std_logic_vector(37, 8),
21109 => conv_std_logic_vector(37, 8),
21110 => conv_std_logic_vector(37, 8),
21111 => conv_std_logic_vector(38, 8),
21112 => conv_std_logic_vector(38, 8),
21113 => conv_std_logic_vector(38, 8),
21114 => conv_std_logic_vector(39, 8),
21115 => conv_std_logic_vector(39, 8),
21116 => conv_std_logic_vector(39, 8),
21117 => conv_std_logic_vector(40, 8),
21118 => conv_std_logic_vector(40, 8),
21119 => conv_std_logic_vector(40, 8),
21120 => conv_std_logic_vector(41, 8),
21121 => conv_std_logic_vector(41, 8),
21122 => conv_std_logic_vector(41, 8),
21123 => conv_std_logic_vector(41, 8),
21124 => conv_std_logic_vector(42, 8),
21125 => conv_std_logic_vector(42, 8),
21126 => conv_std_logic_vector(42, 8),
21127 => conv_std_logic_vector(43, 8),
21128 => conv_std_logic_vector(43, 8),
21129 => conv_std_logic_vector(43, 8),
21130 => conv_std_logic_vector(44, 8),
21131 => conv_std_logic_vector(44, 8),
21132 => conv_std_logic_vector(44, 8),
21133 => conv_std_logic_vector(45, 8),
21134 => conv_std_logic_vector(45, 8),
21135 => conv_std_logic_vector(45, 8),
21136 => conv_std_logic_vector(46, 8),
21137 => conv_std_logic_vector(46, 8),
21138 => conv_std_logic_vector(46, 8),
21139 => conv_std_logic_vector(47, 8),
21140 => conv_std_logic_vector(47, 8),
21141 => conv_std_logic_vector(47, 8),
21142 => conv_std_logic_vector(48, 8),
21143 => conv_std_logic_vector(48, 8),
21144 => conv_std_logic_vector(48, 8),
21145 => conv_std_logic_vector(49, 8),
21146 => conv_std_logic_vector(49, 8),
21147 => conv_std_logic_vector(49, 8),
21148 => conv_std_logic_vector(49, 8),
21149 => conv_std_logic_vector(50, 8),
21150 => conv_std_logic_vector(50, 8),
21151 => conv_std_logic_vector(50, 8),
21152 => conv_std_logic_vector(51, 8),
21153 => conv_std_logic_vector(51, 8),
21154 => conv_std_logic_vector(51, 8),
21155 => conv_std_logic_vector(52, 8),
21156 => conv_std_logic_vector(52, 8),
21157 => conv_std_logic_vector(52, 8),
21158 => conv_std_logic_vector(53, 8),
21159 => conv_std_logic_vector(53, 8),
21160 => conv_std_logic_vector(53, 8),
21161 => conv_std_logic_vector(54, 8),
21162 => conv_std_logic_vector(54, 8),
21163 => conv_std_logic_vector(54, 8),
21164 => conv_std_logic_vector(55, 8),
21165 => conv_std_logic_vector(55, 8),
21166 => conv_std_logic_vector(55, 8),
21167 => conv_std_logic_vector(56, 8),
21168 => conv_std_logic_vector(56, 8),
21169 => conv_std_logic_vector(56, 8),
21170 => conv_std_logic_vector(57, 8),
21171 => conv_std_logic_vector(57, 8),
21172 => conv_std_logic_vector(57, 8),
21173 => conv_std_logic_vector(57, 8),
21174 => conv_std_logic_vector(58, 8),
21175 => conv_std_logic_vector(58, 8),
21176 => conv_std_logic_vector(58, 8),
21177 => conv_std_logic_vector(59, 8),
21178 => conv_std_logic_vector(59, 8),
21179 => conv_std_logic_vector(59, 8),
21180 => conv_std_logic_vector(60, 8),
21181 => conv_std_logic_vector(60, 8),
21182 => conv_std_logic_vector(60, 8),
21183 => conv_std_logic_vector(61, 8),
21184 => conv_std_logic_vector(61, 8),
21185 => conv_std_logic_vector(61, 8),
21186 => conv_std_logic_vector(62, 8),
21187 => conv_std_logic_vector(62, 8),
21188 => conv_std_logic_vector(62, 8),
21189 => conv_std_logic_vector(63, 8),
21190 => conv_std_logic_vector(63, 8),
21191 => conv_std_logic_vector(63, 8),
21192 => conv_std_logic_vector(64, 8),
21193 => conv_std_logic_vector(64, 8),
21194 => conv_std_logic_vector(64, 8),
21195 => conv_std_logic_vector(65, 8),
21196 => conv_std_logic_vector(65, 8),
21197 => conv_std_logic_vector(65, 8),
21198 => conv_std_logic_vector(65, 8),
21199 => conv_std_logic_vector(66, 8),
21200 => conv_std_logic_vector(66, 8),
21201 => conv_std_logic_vector(66, 8),
21202 => conv_std_logic_vector(67, 8),
21203 => conv_std_logic_vector(67, 8),
21204 => conv_std_logic_vector(67, 8),
21205 => conv_std_logic_vector(68, 8),
21206 => conv_std_logic_vector(68, 8),
21207 => conv_std_logic_vector(68, 8),
21208 => conv_std_logic_vector(69, 8),
21209 => conv_std_logic_vector(69, 8),
21210 => conv_std_logic_vector(69, 8),
21211 => conv_std_logic_vector(70, 8),
21212 => conv_std_logic_vector(70, 8),
21213 => conv_std_logic_vector(70, 8),
21214 => conv_std_logic_vector(71, 8),
21215 => conv_std_logic_vector(71, 8),
21216 => conv_std_logic_vector(71, 8),
21217 => conv_std_logic_vector(72, 8),
21218 => conv_std_logic_vector(72, 8),
21219 => conv_std_logic_vector(72, 8),
21220 => conv_std_logic_vector(73, 8),
21221 => conv_std_logic_vector(73, 8),
21222 => conv_std_logic_vector(73, 8),
21223 => conv_std_logic_vector(73, 8),
21224 => conv_std_logic_vector(74, 8),
21225 => conv_std_logic_vector(74, 8),
21226 => conv_std_logic_vector(74, 8),
21227 => conv_std_logic_vector(75, 8),
21228 => conv_std_logic_vector(75, 8),
21229 => conv_std_logic_vector(75, 8),
21230 => conv_std_logic_vector(76, 8),
21231 => conv_std_logic_vector(76, 8),
21232 => conv_std_logic_vector(76, 8),
21233 => conv_std_logic_vector(77, 8),
21234 => conv_std_logic_vector(77, 8),
21235 => conv_std_logic_vector(77, 8),
21236 => conv_std_logic_vector(78, 8),
21237 => conv_std_logic_vector(78, 8),
21238 => conv_std_logic_vector(78, 8),
21239 => conv_std_logic_vector(79, 8),
21240 => conv_std_logic_vector(79, 8),
21241 => conv_std_logic_vector(79, 8),
21242 => conv_std_logic_vector(80, 8),
21243 => conv_std_logic_vector(80, 8),
21244 => conv_std_logic_vector(80, 8),
21245 => conv_std_logic_vector(81, 8),
21246 => conv_std_logic_vector(81, 8),
21247 => conv_std_logic_vector(81, 8),
21248 => conv_std_logic_vector(0, 8),
21249 => conv_std_logic_vector(0, 8),
21250 => conv_std_logic_vector(0, 8),
21251 => conv_std_logic_vector(0, 8),
21252 => conv_std_logic_vector(1, 8),
21253 => conv_std_logic_vector(1, 8),
21254 => conv_std_logic_vector(1, 8),
21255 => conv_std_logic_vector(2, 8),
21256 => conv_std_logic_vector(2, 8),
21257 => conv_std_logic_vector(2, 8),
21258 => conv_std_logic_vector(3, 8),
21259 => conv_std_logic_vector(3, 8),
21260 => conv_std_logic_vector(3, 8),
21261 => conv_std_logic_vector(4, 8),
21262 => conv_std_logic_vector(4, 8),
21263 => conv_std_logic_vector(4, 8),
21264 => conv_std_logic_vector(5, 8),
21265 => conv_std_logic_vector(5, 8),
21266 => conv_std_logic_vector(5, 8),
21267 => conv_std_logic_vector(6, 8),
21268 => conv_std_logic_vector(6, 8),
21269 => conv_std_logic_vector(6, 8),
21270 => conv_std_logic_vector(7, 8),
21271 => conv_std_logic_vector(7, 8),
21272 => conv_std_logic_vector(7, 8),
21273 => conv_std_logic_vector(8, 8),
21274 => conv_std_logic_vector(8, 8),
21275 => conv_std_logic_vector(8, 8),
21276 => conv_std_logic_vector(9, 8),
21277 => conv_std_logic_vector(9, 8),
21278 => conv_std_logic_vector(9, 8),
21279 => conv_std_logic_vector(10, 8),
21280 => conv_std_logic_vector(10, 8),
21281 => conv_std_logic_vector(10, 8),
21282 => conv_std_logic_vector(11, 8),
21283 => conv_std_logic_vector(11, 8),
21284 => conv_std_logic_vector(11, 8),
21285 => conv_std_logic_vector(11, 8),
21286 => conv_std_logic_vector(12, 8),
21287 => conv_std_logic_vector(12, 8),
21288 => conv_std_logic_vector(12, 8),
21289 => conv_std_logic_vector(13, 8),
21290 => conv_std_logic_vector(13, 8),
21291 => conv_std_logic_vector(13, 8),
21292 => conv_std_logic_vector(14, 8),
21293 => conv_std_logic_vector(14, 8),
21294 => conv_std_logic_vector(14, 8),
21295 => conv_std_logic_vector(15, 8),
21296 => conv_std_logic_vector(15, 8),
21297 => conv_std_logic_vector(15, 8),
21298 => conv_std_logic_vector(16, 8),
21299 => conv_std_logic_vector(16, 8),
21300 => conv_std_logic_vector(16, 8),
21301 => conv_std_logic_vector(17, 8),
21302 => conv_std_logic_vector(17, 8),
21303 => conv_std_logic_vector(17, 8),
21304 => conv_std_logic_vector(18, 8),
21305 => conv_std_logic_vector(18, 8),
21306 => conv_std_logic_vector(18, 8),
21307 => conv_std_logic_vector(19, 8),
21308 => conv_std_logic_vector(19, 8),
21309 => conv_std_logic_vector(19, 8),
21310 => conv_std_logic_vector(20, 8),
21311 => conv_std_logic_vector(20, 8),
21312 => conv_std_logic_vector(20, 8),
21313 => conv_std_logic_vector(21, 8),
21314 => conv_std_logic_vector(21, 8),
21315 => conv_std_logic_vector(21, 8),
21316 => conv_std_logic_vector(22, 8),
21317 => conv_std_logic_vector(22, 8),
21318 => conv_std_logic_vector(22, 8),
21319 => conv_std_logic_vector(23, 8),
21320 => conv_std_logic_vector(23, 8),
21321 => conv_std_logic_vector(23, 8),
21322 => conv_std_logic_vector(23, 8),
21323 => conv_std_logic_vector(24, 8),
21324 => conv_std_logic_vector(24, 8),
21325 => conv_std_logic_vector(24, 8),
21326 => conv_std_logic_vector(25, 8),
21327 => conv_std_logic_vector(25, 8),
21328 => conv_std_logic_vector(25, 8),
21329 => conv_std_logic_vector(26, 8),
21330 => conv_std_logic_vector(26, 8),
21331 => conv_std_logic_vector(26, 8),
21332 => conv_std_logic_vector(27, 8),
21333 => conv_std_logic_vector(27, 8),
21334 => conv_std_logic_vector(27, 8),
21335 => conv_std_logic_vector(28, 8),
21336 => conv_std_logic_vector(28, 8),
21337 => conv_std_logic_vector(28, 8),
21338 => conv_std_logic_vector(29, 8),
21339 => conv_std_logic_vector(29, 8),
21340 => conv_std_logic_vector(29, 8),
21341 => conv_std_logic_vector(30, 8),
21342 => conv_std_logic_vector(30, 8),
21343 => conv_std_logic_vector(30, 8),
21344 => conv_std_logic_vector(31, 8),
21345 => conv_std_logic_vector(31, 8),
21346 => conv_std_logic_vector(31, 8),
21347 => conv_std_logic_vector(32, 8),
21348 => conv_std_logic_vector(32, 8),
21349 => conv_std_logic_vector(32, 8),
21350 => conv_std_logic_vector(33, 8),
21351 => conv_std_logic_vector(33, 8),
21352 => conv_std_logic_vector(33, 8),
21353 => conv_std_logic_vector(34, 8),
21354 => conv_std_logic_vector(34, 8),
21355 => conv_std_logic_vector(34, 8),
21356 => conv_std_logic_vector(35, 8),
21357 => conv_std_logic_vector(35, 8),
21358 => conv_std_logic_vector(35, 8),
21359 => conv_std_logic_vector(35, 8),
21360 => conv_std_logic_vector(36, 8),
21361 => conv_std_logic_vector(36, 8),
21362 => conv_std_logic_vector(36, 8),
21363 => conv_std_logic_vector(37, 8),
21364 => conv_std_logic_vector(37, 8),
21365 => conv_std_logic_vector(37, 8),
21366 => conv_std_logic_vector(38, 8),
21367 => conv_std_logic_vector(38, 8),
21368 => conv_std_logic_vector(38, 8),
21369 => conv_std_logic_vector(39, 8),
21370 => conv_std_logic_vector(39, 8),
21371 => conv_std_logic_vector(39, 8),
21372 => conv_std_logic_vector(40, 8),
21373 => conv_std_logic_vector(40, 8),
21374 => conv_std_logic_vector(40, 8),
21375 => conv_std_logic_vector(41, 8),
21376 => conv_std_logic_vector(41, 8),
21377 => conv_std_logic_vector(41, 8),
21378 => conv_std_logic_vector(42, 8),
21379 => conv_std_logic_vector(42, 8),
21380 => conv_std_logic_vector(42, 8),
21381 => conv_std_logic_vector(43, 8),
21382 => conv_std_logic_vector(43, 8),
21383 => conv_std_logic_vector(43, 8),
21384 => conv_std_logic_vector(44, 8),
21385 => conv_std_logic_vector(44, 8),
21386 => conv_std_logic_vector(44, 8),
21387 => conv_std_logic_vector(45, 8),
21388 => conv_std_logic_vector(45, 8),
21389 => conv_std_logic_vector(45, 8),
21390 => conv_std_logic_vector(46, 8),
21391 => conv_std_logic_vector(46, 8),
21392 => conv_std_logic_vector(46, 8),
21393 => conv_std_logic_vector(47, 8),
21394 => conv_std_logic_vector(47, 8),
21395 => conv_std_logic_vector(47, 8),
21396 => conv_std_logic_vector(47, 8),
21397 => conv_std_logic_vector(48, 8),
21398 => conv_std_logic_vector(48, 8),
21399 => conv_std_logic_vector(48, 8),
21400 => conv_std_logic_vector(49, 8),
21401 => conv_std_logic_vector(49, 8),
21402 => conv_std_logic_vector(49, 8),
21403 => conv_std_logic_vector(50, 8),
21404 => conv_std_logic_vector(50, 8),
21405 => conv_std_logic_vector(50, 8),
21406 => conv_std_logic_vector(51, 8),
21407 => conv_std_logic_vector(51, 8),
21408 => conv_std_logic_vector(51, 8),
21409 => conv_std_logic_vector(52, 8),
21410 => conv_std_logic_vector(52, 8),
21411 => conv_std_logic_vector(52, 8),
21412 => conv_std_logic_vector(53, 8),
21413 => conv_std_logic_vector(53, 8),
21414 => conv_std_logic_vector(53, 8),
21415 => conv_std_logic_vector(54, 8),
21416 => conv_std_logic_vector(54, 8),
21417 => conv_std_logic_vector(54, 8),
21418 => conv_std_logic_vector(55, 8),
21419 => conv_std_logic_vector(55, 8),
21420 => conv_std_logic_vector(55, 8),
21421 => conv_std_logic_vector(56, 8),
21422 => conv_std_logic_vector(56, 8),
21423 => conv_std_logic_vector(56, 8),
21424 => conv_std_logic_vector(57, 8),
21425 => conv_std_logic_vector(57, 8),
21426 => conv_std_logic_vector(57, 8),
21427 => conv_std_logic_vector(58, 8),
21428 => conv_std_logic_vector(58, 8),
21429 => conv_std_logic_vector(58, 8),
21430 => conv_std_logic_vector(59, 8),
21431 => conv_std_logic_vector(59, 8),
21432 => conv_std_logic_vector(59, 8),
21433 => conv_std_logic_vector(59, 8),
21434 => conv_std_logic_vector(60, 8),
21435 => conv_std_logic_vector(60, 8),
21436 => conv_std_logic_vector(60, 8),
21437 => conv_std_logic_vector(61, 8),
21438 => conv_std_logic_vector(61, 8),
21439 => conv_std_logic_vector(61, 8),
21440 => conv_std_logic_vector(62, 8),
21441 => conv_std_logic_vector(62, 8),
21442 => conv_std_logic_vector(62, 8),
21443 => conv_std_logic_vector(63, 8),
21444 => conv_std_logic_vector(63, 8),
21445 => conv_std_logic_vector(63, 8),
21446 => conv_std_logic_vector(64, 8),
21447 => conv_std_logic_vector(64, 8),
21448 => conv_std_logic_vector(64, 8),
21449 => conv_std_logic_vector(65, 8),
21450 => conv_std_logic_vector(65, 8),
21451 => conv_std_logic_vector(65, 8),
21452 => conv_std_logic_vector(66, 8),
21453 => conv_std_logic_vector(66, 8),
21454 => conv_std_logic_vector(66, 8),
21455 => conv_std_logic_vector(67, 8),
21456 => conv_std_logic_vector(67, 8),
21457 => conv_std_logic_vector(67, 8),
21458 => conv_std_logic_vector(68, 8),
21459 => conv_std_logic_vector(68, 8),
21460 => conv_std_logic_vector(68, 8),
21461 => conv_std_logic_vector(69, 8),
21462 => conv_std_logic_vector(69, 8),
21463 => conv_std_logic_vector(69, 8),
21464 => conv_std_logic_vector(70, 8),
21465 => conv_std_logic_vector(70, 8),
21466 => conv_std_logic_vector(70, 8),
21467 => conv_std_logic_vector(71, 8),
21468 => conv_std_logic_vector(71, 8),
21469 => conv_std_logic_vector(71, 8),
21470 => conv_std_logic_vector(71, 8),
21471 => conv_std_logic_vector(72, 8),
21472 => conv_std_logic_vector(72, 8),
21473 => conv_std_logic_vector(72, 8),
21474 => conv_std_logic_vector(73, 8),
21475 => conv_std_logic_vector(73, 8),
21476 => conv_std_logic_vector(73, 8),
21477 => conv_std_logic_vector(74, 8),
21478 => conv_std_logic_vector(74, 8),
21479 => conv_std_logic_vector(74, 8),
21480 => conv_std_logic_vector(75, 8),
21481 => conv_std_logic_vector(75, 8),
21482 => conv_std_logic_vector(75, 8),
21483 => conv_std_logic_vector(76, 8),
21484 => conv_std_logic_vector(76, 8),
21485 => conv_std_logic_vector(76, 8),
21486 => conv_std_logic_vector(77, 8),
21487 => conv_std_logic_vector(77, 8),
21488 => conv_std_logic_vector(77, 8),
21489 => conv_std_logic_vector(78, 8),
21490 => conv_std_logic_vector(78, 8),
21491 => conv_std_logic_vector(78, 8),
21492 => conv_std_logic_vector(79, 8),
21493 => conv_std_logic_vector(79, 8),
21494 => conv_std_logic_vector(79, 8),
21495 => conv_std_logic_vector(80, 8),
21496 => conv_std_logic_vector(80, 8),
21497 => conv_std_logic_vector(80, 8),
21498 => conv_std_logic_vector(81, 8),
21499 => conv_std_logic_vector(81, 8),
21500 => conv_std_logic_vector(81, 8),
21501 => conv_std_logic_vector(82, 8),
21502 => conv_std_logic_vector(82, 8),
21503 => conv_std_logic_vector(82, 8),
21504 => conv_std_logic_vector(0, 8),
21505 => conv_std_logic_vector(0, 8),
21506 => conv_std_logic_vector(0, 8),
21507 => conv_std_logic_vector(0, 8),
21508 => conv_std_logic_vector(1, 8),
21509 => conv_std_logic_vector(1, 8),
21510 => conv_std_logic_vector(1, 8),
21511 => conv_std_logic_vector(2, 8),
21512 => conv_std_logic_vector(2, 8),
21513 => conv_std_logic_vector(2, 8),
21514 => conv_std_logic_vector(3, 8),
21515 => conv_std_logic_vector(3, 8),
21516 => conv_std_logic_vector(3, 8),
21517 => conv_std_logic_vector(4, 8),
21518 => conv_std_logic_vector(4, 8),
21519 => conv_std_logic_vector(4, 8),
21520 => conv_std_logic_vector(5, 8),
21521 => conv_std_logic_vector(5, 8),
21522 => conv_std_logic_vector(5, 8),
21523 => conv_std_logic_vector(6, 8),
21524 => conv_std_logic_vector(6, 8),
21525 => conv_std_logic_vector(6, 8),
21526 => conv_std_logic_vector(7, 8),
21527 => conv_std_logic_vector(7, 8),
21528 => conv_std_logic_vector(7, 8),
21529 => conv_std_logic_vector(8, 8),
21530 => conv_std_logic_vector(8, 8),
21531 => conv_std_logic_vector(8, 8),
21532 => conv_std_logic_vector(9, 8),
21533 => conv_std_logic_vector(9, 8),
21534 => conv_std_logic_vector(9, 8),
21535 => conv_std_logic_vector(10, 8),
21536 => conv_std_logic_vector(10, 8),
21537 => conv_std_logic_vector(10, 8),
21538 => conv_std_logic_vector(11, 8),
21539 => conv_std_logic_vector(11, 8),
21540 => conv_std_logic_vector(11, 8),
21541 => conv_std_logic_vector(12, 8),
21542 => conv_std_logic_vector(12, 8),
21543 => conv_std_logic_vector(12, 8),
21544 => conv_std_logic_vector(13, 8),
21545 => conv_std_logic_vector(13, 8),
21546 => conv_std_logic_vector(13, 8),
21547 => conv_std_logic_vector(14, 8),
21548 => conv_std_logic_vector(14, 8),
21549 => conv_std_logic_vector(14, 8),
21550 => conv_std_logic_vector(15, 8),
21551 => conv_std_logic_vector(15, 8),
21552 => conv_std_logic_vector(15, 8),
21553 => conv_std_logic_vector(16, 8),
21554 => conv_std_logic_vector(16, 8),
21555 => conv_std_logic_vector(16, 8),
21556 => conv_std_logic_vector(17, 8),
21557 => conv_std_logic_vector(17, 8),
21558 => conv_std_logic_vector(17, 8),
21559 => conv_std_logic_vector(18, 8),
21560 => conv_std_logic_vector(18, 8),
21561 => conv_std_logic_vector(18, 8),
21562 => conv_std_logic_vector(19, 8),
21563 => conv_std_logic_vector(19, 8),
21564 => conv_std_logic_vector(19, 8),
21565 => conv_std_logic_vector(20, 8),
21566 => conv_std_logic_vector(20, 8),
21567 => conv_std_logic_vector(20, 8),
21568 => conv_std_logic_vector(21, 8),
21569 => conv_std_logic_vector(21, 8),
21570 => conv_std_logic_vector(21, 8),
21571 => conv_std_logic_vector(21, 8),
21572 => conv_std_logic_vector(22, 8),
21573 => conv_std_logic_vector(22, 8),
21574 => conv_std_logic_vector(22, 8),
21575 => conv_std_logic_vector(23, 8),
21576 => conv_std_logic_vector(23, 8),
21577 => conv_std_logic_vector(23, 8),
21578 => conv_std_logic_vector(24, 8),
21579 => conv_std_logic_vector(24, 8),
21580 => conv_std_logic_vector(24, 8),
21581 => conv_std_logic_vector(25, 8),
21582 => conv_std_logic_vector(25, 8),
21583 => conv_std_logic_vector(25, 8),
21584 => conv_std_logic_vector(26, 8),
21585 => conv_std_logic_vector(26, 8),
21586 => conv_std_logic_vector(26, 8),
21587 => conv_std_logic_vector(27, 8),
21588 => conv_std_logic_vector(27, 8),
21589 => conv_std_logic_vector(27, 8),
21590 => conv_std_logic_vector(28, 8),
21591 => conv_std_logic_vector(28, 8),
21592 => conv_std_logic_vector(28, 8),
21593 => conv_std_logic_vector(29, 8),
21594 => conv_std_logic_vector(29, 8),
21595 => conv_std_logic_vector(29, 8),
21596 => conv_std_logic_vector(30, 8),
21597 => conv_std_logic_vector(30, 8),
21598 => conv_std_logic_vector(30, 8),
21599 => conv_std_logic_vector(31, 8),
21600 => conv_std_logic_vector(31, 8),
21601 => conv_std_logic_vector(31, 8),
21602 => conv_std_logic_vector(32, 8),
21603 => conv_std_logic_vector(32, 8),
21604 => conv_std_logic_vector(32, 8),
21605 => conv_std_logic_vector(33, 8),
21606 => conv_std_logic_vector(33, 8),
21607 => conv_std_logic_vector(33, 8),
21608 => conv_std_logic_vector(34, 8),
21609 => conv_std_logic_vector(34, 8),
21610 => conv_std_logic_vector(34, 8),
21611 => conv_std_logic_vector(35, 8),
21612 => conv_std_logic_vector(35, 8),
21613 => conv_std_logic_vector(35, 8),
21614 => conv_std_logic_vector(36, 8),
21615 => conv_std_logic_vector(36, 8),
21616 => conv_std_logic_vector(36, 8),
21617 => conv_std_logic_vector(37, 8),
21618 => conv_std_logic_vector(37, 8),
21619 => conv_std_logic_vector(37, 8),
21620 => conv_std_logic_vector(38, 8),
21621 => conv_std_logic_vector(38, 8),
21622 => conv_std_logic_vector(38, 8),
21623 => conv_std_logic_vector(39, 8),
21624 => conv_std_logic_vector(39, 8),
21625 => conv_std_logic_vector(39, 8),
21626 => conv_std_logic_vector(40, 8),
21627 => conv_std_logic_vector(40, 8),
21628 => conv_std_logic_vector(40, 8),
21629 => conv_std_logic_vector(41, 8),
21630 => conv_std_logic_vector(41, 8),
21631 => conv_std_logic_vector(41, 8),
21632 => conv_std_logic_vector(42, 8),
21633 => conv_std_logic_vector(42, 8),
21634 => conv_std_logic_vector(42, 8),
21635 => conv_std_logic_vector(42, 8),
21636 => conv_std_logic_vector(43, 8),
21637 => conv_std_logic_vector(43, 8),
21638 => conv_std_logic_vector(43, 8),
21639 => conv_std_logic_vector(44, 8),
21640 => conv_std_logic_vector(44, 8),
21641 => conv_std_logic_vector(44, 8),
21642 => conv_std_logic_vector(45, 8),
21643 => conv_std_logic_vector(45, 8),
21644 => conv_std_logic_vector(45, 8),
21645 => conv_std_logic_vector(46, 8),
21646 => conv_std_logic_vector(46, 8),
21647 => conv_std_logic_vector(46, 8),
21648 => conv_std_logic_vector(47, 8),
21649 => conv_std_logic_vector(47, 8),
21650 => conv_std_logic_vector(47, 8),
21651 => conv_std_logic_vector(48, 8),
21652 => conv_std_logic_vector(48, 8),
21653 => conv_std_logic_vector(48, 8),
21654 => conv_std_logic_vector(49, 8),
21655 => conv_std_logic_vector(49, 8),
21656 => conv_std_logic_vector(49, 8),
21657 => conv_std_logic_vector(50, 8),
21658 => conv_std_logic_vector(50, 8),
21659 => conv_std_logic_vector(50, 8),
21660 => conv_std_logic_vector(51, 8),
21661 => conv_std_logic_vector(51, 8),
21662 => conv_std_logic_vector(51, 8),
21663 => conv_std_logic_vector(52, 8),
21664 => conv_std_logic_vector(52, 8),
21665 => conv_std_logic_vector(52, 8),
21666 => conv_std_logic_vector(53, 8),
21667 => conv_std_logic_vector(53, 8),
21668 => conv_std_logic_vector(53, 8),
21669 => conv_std_logic_vector(54, 8),
21670 => conv_std_logic_vector(54, 8),
21671 => conv_std_logic_vector(54, 8),
21672 => conv_std_logic_vector(55, 8),
21673 => conv_std_logic_vector(55, 8),
21674 => conv_std_logic_vector(55, 8),
21675 => conv_std_logic_vector(56, 8),
21676 => conv_std_logic_vector(56, 8),
21677 => conv_std_logic_vector(56, 8),
21678 => conv_std_logic_vector(57, 8),
21679 => conv_std_logic_vector(57, 8),
21680 => conv_std_logic_vector(57, 8),
21681 => conv_std_logic_vector(58, 8),
21682 => conv_std_logic_vector(58, 8),
21683 => conv_std_logic_vector(58, 8),
21684 => conv_std_logic_vector(59, 8),
21685 => conv_std_logic_vector(59, 8),
21686 => conv_std_logic_vector(59, 8),
21687 => conv_std_logic_vector(60, 8),
21688 => conv_std_logic_vector(60, 8),
21689 => conv_std_logic_vector(60, 8),
21690 => conv_std_logic_vector(61, 8),
21691 => conv_std_logic_vector(61, 8),
21692 => conv_std_logic_vector(61, 8),
21693 => conv_std_logic_vector(62, 8),
21694 => conv_std_logic_vector(62, 8),
21695 => conv_std_logic_vector(62, 8),
21696 => conv_std_logic_vector(63, 8),
21697 => conv_std_logic_vector(63, 8),
21698 => conv_std_logic_vector(63, 8),
21699 => conv_std_logic_vector(63, 8),
21700 => conv_std_logic_vector(64, 8),
21701 => conv_std_logic_vector(64, 8),
21702 => conv_std_logic_vector(64, 8),
21703 => conv_std_logic_vector(65, 8),
21704 => conv_std_logic_vector(65, 8),
21705 => conv_std_logic_vector(65, 8),
21706 => conv_std_logic_vector(66, 8),
21707 => conv_std_logic_vector(66, 8),
21708 => conv_std_logic_vector(66, 8),
21709 => conv_std_logic_vector(67, 8),
21710 => conv_std_logic_vector(67, 8),
21711 => conv_std_logic_vector(67, 8),
21712 => conv_std_logic_vector(68, 8),
21713 => conv_std_logic_vector(68, 8),
21714 => conv_std_logic_vector(68, 8),
21715 => conv_std_logic_vector(69, 8),
21716 => conv_std_logic_vector(69, 8),
21717 => conv_std_logic_vector(69, 8),
21718 => conv_std_logic_vector(70, 8),
21719 => conv_std_logic_vector(70, 8),
21720 => conv_std_logic_vector(70, 8),
21721 => conv_std_logic_vector(71, 8),
21722 => conv_std_logic_vector(71, 8),
21723 => conv_std_logic_vector(71, 8),
21724 => conv_std_logic_vector(72, 8),
21725 => conv_std_logic_vector(72, 8),
21726 => conv_std_logic_vector(72, 8),
21727 => conv_std_logic_vector(73, 8),
21728 => conv_std_logic_vector(73, 8),
21729 => conv_std_logic_vector(73, 8),
21730 => conv_std_logic_vector(74, 8),
21731 => conv_std_logic_vector(74, 8),
21732 => conv_std_logic_vector(74, 8),
21733 => conv_std_logic_vector(75, 8),
21734 => conv_std_logic_vector(75, 8),
21735 => conv_std_logic_vector(75, 8),
21736 => conv_std_logic_vector(76, 8),
21737 => conv_std_logic_vector(76, 8),
21738 => conv_std_logic_vector(76, 8),
21739 => conv_std_logic_vector(77, 8),
21740 => conv_std_logic_vector(77, 8),
21741 => conv_std_logic_vector(77, 8),
21742 => conv_std_logic_vector(78, 8),
21743 => conv_std_logic_vector(78, 8),
21744 => conv_std_logic_vector(78, 8),
21745 => conv_std_logic_vector(79, 8),
21746 => conv_std_logic_vector(79, 8),
21747 => conv_std_logic_vector(79, 8),
21748 => conv_std_logic_vector(80, 8),
21749 => conv_std_logic_vector(80, 8),
21750 => conv_std_logic_vector(80, 8),
21751 => conv_std_logic_vector(81, 8),
21752 => conv_std_logic_vector(81, 8),
21753 => conv_std_logic_vector(81, 8),
21754 => conv_std_logic_vector(82, 8),
21755 => conv_std_logic_vector(82, 8),
21756 => conv_std_logic_vector(82, 8),
21757 => conv_std_logic_vector(83, 8),
21758 => conv_std_logic_vector(83, 8),
21759 => conv_std_logic_vector(83, 8),
21760 => conv_std_logic_vector(0, 8),
21761 => conv_std_logic_vector(0, 8),
21762 => conv_std_logic_vector(0, 8),
21763 => conv_std_logic_vector(0, 8),
21764 => conv_std_logic_vector(1, 8),
21765 => conv_std_logic_vector(1, 8),
21766 => conv_std_logic_vector(1, 8),
21767 => conv_std_logic_vector(2, 8),
21768 => conv_std_logic_vector(2, 8),
21769 => conv_std_logic_vector(2, 8),
21770 => conv_std_logic_vector(3, 8),
21771 => conv_std_logic_vector(3, 8),
21772 => conv_std_logic_vector(3, 8),
21773 => conv_std_logic_vector(4, 8),
21774 => conv_std_logic_vector(4, 8),
21775 => conv_std_logic_vector(4, 8),
21776 => conv_std_logic_vector(5, 8),
21777 => conv_std_logic_vector(5, 8),
21778 => conv_std_logic_vector(5, 8),
21779 => conv_std_logic_vector(6, 8),
21780 => conv_std_logic_vector(6, 8),
21781 => conv_std_logic_vector(6, 8),
21782 => conv_std_logic_vector(7, 8),
21783 => conv_std_logic_vector(7, 8),
21784 => conv_std_logic_vector(7, 8),
21785 => conv_std_logic_vector(8, 8),
21786 => conv_std_logic_vector(8, 8),
21787 => conv_std_logic_vector(8, 8),
21788 => conv_std_logic_vector(9, 8),
21789 => conv_std_logic_vector(9, 8),
21790 => conv_std_logic_vector(9, 8),
21791 => conv_std_logic_vector(10, 8),
21792 => conv_std_logic_vector(10, 8),
21793 => conv_std_logic_vector(10, 8),
21794 => conv_std_logic_vector(11, 8),
21795 => conv_std_logic_vector(11, 8),
21796 => conv_std_logic_vector(11, 8),
21797 => conv_std_logic_vector(12, 8),
21798 => conv_std_logic_vector(12, 8),
21799 => conv_std_logic_vector(12, 8),
21800 => conv_std_logic_vector(13, 8),
21801 => conv_std_logic_vector(13, 8),
21802 => conv_std_logic_vector(13, 8),
21803 => conv_std_logic_vector(14, 8),
21804 => conv_std_logic_vector(14, 8),
21805 => conv_std_logic_vector(14, 8),
21806 => conv_std_logic_vector(15, 8),
21807 => conv_std_logic_vector(15, 8),
21808 => conv_std_logic_vector(15, 8),
21809 => conv_std_logic_vector(16, 8),
21810 => conv_std_logic_vector(16, 8),
21811 => conv_std_logic_vector(16, 8),
21812 => conv_std_logic_vector(17, 8),
21813 => conv_std_logic_vector(17, 8),
21814 => conv_std_logic_vector(17, 8),
21815 => conv_std_logic_vector(18, 8),
21816 => conv_std_logic_vector(18, 8),
21817 => conv_std_logic_vector(18, 8),
21818 => conv_std_logic_vector(19, 8),
21819 => conv_std_logic_vector(19, 8),
21820 => conv_std_logic_vector(19, 8),
21821 => conv_std_logic_vector(20, 8),
21822 => conv_std_logic_vector(20, 8),
21823 => conv_std_logic_vector(20, 8),
21824 => conv_std_logic_vector(21, 8),
21825 => conv_std_logic_vector(21, 8),
21826 => conv_std_logic_vector(21, 8),
21827 => conv_std_logic_vector(22, 8),
21828 => conv_std_logic_vector(22, 8),
21829 => conv_std_logic_vector(22, 8),
21830 => conv_std_logic_vector(23, 8),
21831 => conv_std_logic_vector(23, 8),
21832 => conv_std_logic_vector(23, 8),
21833 => conv_std_logic_vector(24, 8),
21834 => conv_std_logic_vector(24, 8),
21835 => conv_std_logic_vector(24, 8),
21836 => conv_std_logic_vector(25, 8),
21837 => conv_std_logic_vector(25, 8),
21838 => conv_std_logic_vector(25, 8),
21839 => conv_std_logic_vector(26, 8),
21840 => conv_std_logic_vector(26, 8),
21841 => conv_std_logic_vector(26, 8),
21842 => conv_std_logic_vector(27, 8),
21843 => conv_std_logic_vector(27, 8),
21844 => conv_std_logic_vector(27, 8),
21845 => conv_std_logic_vector(28, 8),
21846 => conv_std_logic_vector(28, 8),
21847 => conv_std_logic_vector(28, 8),
21848 => conv_std_logic_vector(29, 8),
21849 => conv_std_logic_vector(29, 8),
21850 => conv_std_logic_vector(29, 8),
21851 => conv_std_logic_vector(30, 8),
21852 => conv_std_logic_vector(30, 8),
21853 => conv_std_logic_vector(30, 8),
21854 => conv_std_logic_vector(31, 8),
21855 => conv_std_logic_vector(31, 8),
21856 => conv_std_logic_vector(31, 8),
21857 => conv_std_logic_vector(32, 8),
21858 => conv_std_logic_vector(32, 8),
21859 => conv_std_logic_vector(32, 8),
21860 => conv_std_logic_vector(33, 8),
21861 => conv_std_logic_vector(33, 8),
21862 => conv_std_logic_vector(33, 8),
21863 => conv_std_logic_vector(34, 8),
21864 => conv_std_logic_vector(34, 8),
21865 => conv_std_logic_vector(34, 8),
21866 => conv_std_logic_vector(35, 8),
21867 => conv_std_logic_vector(35, 8),
21868 => conv_std_logic_vector(35, 8),
21869 => conv_std_logic_vector(36, 8),
21870 => conv_std_logic_vector(36, 8),
21871 => conv_std_logic_vector(36, 8),
21872 => conv_std_logic_vector(37, 8),
21873 => conv_std_logic_vector(37, 8),
21874 => conv_std_logic_vector(37, 8),
21875 => conv_std_logic_vector(38, 8),
21876 => conv_std_logic_vector(38, 8),
21877 => conv_std_logic_vector(38, 8),
21878 => conv_std_logic_vector(39, 8),
21879 => conv_std_logic_vector(39, 8),
21880 => conv_std_logic_vector(39, 8),
21881 => conv_std_logic_vector(40, 8),
21882 => conv_std_logic_vector(40, 8),
21883 => conv_std_logic_vector(40, 8),
21884 => conv_std_logic_vector(41, 8),
21885 => conv_std_logic_vector(41, 8),
21886 => conv_std_logic_vector(41, 8),
21887 => conv_std_logic_vector(42, 8),
21888 => conv_std_logic_vector(42, 8),
21889 => conv_std_logic_vector(42, 8),
21890 => conv_std_logic_vector(43, 8),
21891 => conv_std_logic_vector(43, 8),
21892 => conv_std_logic_vector(43, 8),
21893 => conv_std_logic_vector(44, 8),
21894 => conv_std_logic_vector(44, 8),
21895 => conv_std_logic_vector(44, 8),
21896 => conv_std_logic_vector(45, 8),
21897 => conv_std_logic_vector(45, 8),
21898 => conv_std_logic_vector(45, 8),
21899 => conv_std_logic_vector(46, 8),
21900 => conv_std_logic_vector(46, 8),
21901 => conv_std_logic_vector(46, 8),
21902 => conv_std_logic_vector(47, 8),
21903 => conv_std_logic_vector(47, 8),
21904 => conv_std_logic_vector(47, 8),
21905 => conv_std_logic_vector(48, 8),
21906 => conv_std_logic_vector(48, 8),
21907 => conv_std_logic_vector(48, 8),
21908 => conv_std_logic_vector(49, 8),
21909 => conv_std_logic_vector(49, 8),
21910 => conv_std_logic_vector(49, 8),
21911 => conv_std_logic_vector(50, 8),
21912 => conv_std_logic_vector(50, 8),
21913 => conv_std_logic_vector(50, 8),
21914 => conv_std_logic_vector(51, 8),
21915 => conv_std_logic_vector(51, 8),
21916 => conv_std_logic_vector(51, 8),
21917 => conv_std_logic_vector(52, 8),
21918 => conv_std_logic_vector(52, 8),
21919 => conv_std_logic_vector(52, 8),
21920 => conv_std_logic_vector(53, 8),
21921 => conv_std_logic_vector(53, 8),
21922 => conv_std_logic_vector(53, 8),
21923 => conv_std_logic_vector(54, 8),
21924 => conv_std_logic_vector(54, 8),
21925 => conv_std_logic_vector(54, 8),
21926 => conv_std_logic_vector(55, 8),
21927 => conv_std_logic_vector(55, 8),
21928 => conv_std_logic_vector(55, 8),
21929 => conv_std_logic_vector(56, 8),
21930 => conv_std_logic_vector(56, 8),
21931 => conv_std_logic_vector(56, 8),
21932 => conv_std_logic_vector(57, 8),
21933 => conv_std_logic_vector(57, 8),
21934 => conv_std_logic_vector(57, 8),
21935 => conv_std_logic_vector(58, 8),
21936 => conv_std_logic_vector(58, 8),
21937 => conv_std_logic_vector(58, 8),
21938 => conv_std_logic_vector(59, 8),
21939 => conv_std_logic_vector(59, 8),
21940 => conv_std_logic_vector(59, 8),
21941 => conv_std_logic_vector(60, 8),
21942 => conv_std_logic_vector(60, 8),
21943 => conv_std_logic_vector(60, 8),
21944 => conv_std_logic_vector(61, 8),
21945 => conv_std_logic_vector(61, 8),
21946 => conv_std_logic_vector(61, 8),
21947 => conv_std_logic_vector(62, 8),
21948 => conv_std_logic_vector(62, 8),
21949 => conv_std_logic_vector(62, 8),
21950 => conv_std_logic_vector(63, 8),
21951 => conv_std_logic_vector(63, 8),
21952 => conv_std_logic_vector(63, 8),
21953 => conv_std_logic_vector(64, 8),
21954 => conv_std_logic_vector(64, 8),
21955 => conv_std_logic_vector(64, 8),
21956 => conv_std_logic_vector(65, 8),
21957 => conv_std_logic_vector(65, 8),
21958 => conv_std_logic_vector(65, 8),
21959 => conv_std_logic_vector(66, 8),
21960 => conv_std_logic_vector(66, 8),
21961 => conv_std_logic_vector(66, 8),
21962 => conv_std_logic_vector(67, 8),
21963 => conv_std_logic_vector(67, 8),
21964 => conv_std_logic_vector(67, 8),
21965 => conv_std_logic_vector(68, 8),
21966 => conv_std_logic_vector(68, 8),
21967 => conv_std_logic_vector(68, 8),
21968 => conv_std_logic_vector(69, 8),
21969 => conv_std_logic_vector(69, 8),
21970 => conv_std_logic_vector(69, 8),
21971 => conv_std_logic_vector(70, 8),
21972 => conv_std_logic_vector(70, 8),
21973 => conv_std_logic_vector(70, 8),
21974 => conv_std_logic_vector(71, 8),
21975 => conv_std_logic_vector(71, 8),
21976 => conv_std_logic_vector(71, 8),
21977 => conv_std_logic_vector(72, 8),
21978 => conv_std_logic_vector(72, 8),
21979 => conv_std_logic_vector(72, 8),
21980 => conv_std_logic_vector(73, 8),
21981 => conv_std_logic_vector(73, 8),
21982 => conv_std_logic_vector(73, 8),
21983 => conv_std_logic_vector(74, 8),
21984 => conv_std_logic_vector(74, 8),
21985 => conv_std_logic_vector(74, 8),
21986 => conv_std_logic_vector(75, 8),
21987 => conv_std_logic_vector(75, 8),
21988 => conv_std_logic_vector(75, 8),
21989 => conv_std_logic_vector(76, 8),
21990 => conv_std_logic_vector(76, 8),
21991 => conv_std_logic_vector(76, 8),
21992 => conv_std_logic_vector(77, 8),
21993 => conv_std_logic_vector(77, 8),
21994 => conv_std_logic_vector(77, 8),
21995 => conv_std_logic_vector(78, 8),
21996 => conv_std_logic_vector(78, 8),
21997 => conv_std_logic_vector(78, 8),
21998 => conv_std_logic_vector(79, 8),
21999 => conv_std_logic_vector(79, 8),
22000 => conv_std_logic_vector(79, 8),
22001 => conv_std_logic_vector(80, 8),
22002 => conv_std_logic_vector(80, 8),
22003 => conv_std_logic_vector(80, 8),
22004 => conv_std_logic_vector(81, 8),
22005 => conv_std_logic_vector(81, 8),
22006 => conv_std_logic_vector(81, 8),
22007 => conv_std_logic_vector(82, 8),
22008 => conv_std_logic_vector(82, 8),
22009 => conv_std_logic_vector(82, 8),
22010 => conv_std_logic_vector(83, 8),
22011 => conv_std_logic_vector(83, 8),
22012 => conv_std_logic_vector(83, 8),
22013 => conv_std_logic_vector(84, 8),
22014 => conv_std_logic_vector(84, 8),
22015 => conv_std_logic_vector(84, 8),
22016 => conv_std_logic_vector(0, 8),
22017 => conv_std_logic_vector(0, 8),
22018 => conv_std_logic_vector(0, 8),
22019 => conv_std_logic_vector(1, 8),
22020 => conv_std_logic_vector(1, 8),
22021 => conv_std_logic_vector(1, 8),
22022 => conv_std_logic_vector(2, 8),
22023 => conv_std_logic_vector(2, 8),
22024 => conv_std_logic_vector(2, 8),
22025 => conv_std_logic_vector(3, 8),
22026 => conv_std_logic_vector(3, 8),
22027 => conv_std_logic_vector(3, 8),
22028 => conv_std_logic_vector(4, 8),
22029 => conv_std_logic_vector(4, 8),
22030 => conv_std_logic_vector(4, 8),
22031 => conv_std_logic_vector(5, 8),
22032 => conv_std_logic_vector(5, 8),
22033 => conv_std_logic_vector(5, 8),
22034 => conv_std_logic_vector(6, 8),
22035 => conv_std_logic_vector(6, 8),
22036 => conv_std_logic_vector(6, 8),
22037 => conv_std_logic_vector(7, 8),
22038 => conv_std_logic_vector(7, 8),
22039 => conv_std_logic_vector(7, 8),
22040 => conv_std_logic_vector(8, 8),
22041 => conv_std_logic_vector(8, 8),
22042 => conv_std_logic_vector(8, 8),
22043 => conv_std_logic_vector(9, 8),
22044 => conv_std_logic_vector(9, 8),
22045 => conv_std_logic_vector(9, 8),
22046 => conv_std_logic_vector(10, 8),
22047 => conv_std_logic_vector(10, 8),
22048 => conv_std_logic_vector(10, 8),
22049 => conv_std_logic_vector(11, 8),
22050 => conv_std_logic_vector(11, 8),
22051 => conv_std_logic_vector(11, 8),
22052 => conv_std_logic_vector(12, 8),
22053 => conv_std_logic_vector(12, 8),
22054 => conv_std_logic_vector(12, 8),
22055 => conv_std_logic_vector(13, 8),
22056 => conv_std_logic_vector(13, 8),
22057 => conv_std_logic_vector(13, 8),
22058 => conv_std_logic_vector(14, 8),
22059 => conv_std_logic_vector(14, 8),
22060 => conv_std_logic_vector(14, 8),
22061 => conv_std_logic_vector(15, 8),
22062 => conv_std_logic_vector(15, 8),
22063 => conv_std_logic_vector(15, 8),
22064 => conv_std_logic_vector(16, 8),
22065 => conv_std_logic_vector(16, 8),
22066 => conv_std_logic_vector(16, 8),
22067 => conv_std_logic_vector(17, 8),
22068 => conv_std_logic_vector(17, 8),
22069 => conv_std_logic_vector(17, 8),
22070 => conv_std_logic_vector(18, 8),
22071 => conv_std_logic_vector(18, 8),
22072 => conv_std_logic_vector(18, 8),
22073 => conv_std_logic_vector(19, 8),
22074 => conv_std_logic_vector(19, 8),
22075 => conv_std_logic_vector(19, 8),
22076 => conv_std_logic_vector(20, 8),
22077 => conv_std_logic_vector(20, 8),
22078 => conv_std_logic_vector(20, 8),
22079 => conv_std_logic_vector(21, 8),
22080 => conv_std_logic_vector(21, 8),
22081 => conv_std_logic_vector(21, 8),
22082 => conv_std_logic_vector(22, 8),
22083 => conv_std_logic_vector(22, 8),
22084 => conv_std_logic_vector(22, 8),
22085 => conv_std_logic_vector(23, 8),
22086 => conv_std_logic_vector(23, 8),
22087 => conv_std_logic_vector(23, 8),
22088 => conv_std_logic_vector(24, 8),
22089 => conv_std_logic_vector(24, 8),
22090 => conv_std_logic_vector(24, 8),
22091 => conv_std_logic_vector(25, 8),
22092 => conv_std_logic_vector(25, 8),
22093 => conv_std_logic_vector(25, 8),
22094 => conv_std_logic_vector(26, 8),
22095 => conv_std_logic_vector(26, 8),
22096 => conv_std_logic_vector(26, 8),
22097 => conv_std_logic_vector(27, 8),
22098 => conv_std_logic_vector(27, 8),
22099 => conv_std_logic_vector(27, 8),
22100 => conv_std_logic_vector(28, 8),
22101 => conv_std_logic_vector(28, 8),
22102 => conv_std_logic_vector(28, 8),
22103 => conv_std_logic_vector(29, 8),
22104 => conv_std_logic_vector(29, 8),
22105 => conv_std_logic_vector(29, 8),
22106 => conv_std_logic_vector(30, 8),
22107 => conv_std_logic_vector(30, 8),
22108 => conv_std_logic_vector(30, 8),
22109 => conv_std_logic_vector(31, 8),
22110 => conv_std_logic_vector(31, 8),
22111 => conv_std_logic_vector(31, 8),
22112 => conv_std_logic_vector(32, 8),
22113 => conv_std_logic_vector(32, 8),
22114 => conv_std_logic_vector(32, 8),
22115 => conv_std_logic_vector(33, 8),
22116 => conv_std_logic_vector(33, 8),
22117 => conv_std_logic_vector(33, 8),
22118 => conv_std_logic_vector(34, 8),
22119 => conv_std_logic_vector(34, 8),
22120 => conv_std_logic_vector(34, 8),
22121 => conv_std_logic_vector(35, 8),
22122 => conv_std_logic_vector(35, 8),
22123 => conv_std_logic_vector(35, 8),
22124 => conv_std_logic_vector(36, 8),
22125 => conv_std_logic_vector(36, 8),
22126 => conv_std_logic_vector(36, 8),
22127 => conv_std_logic_vector(37, 8),
22128 => conv_std_logic_vector(37, 8),
22129 => conv_std_logic_vector(37, 8),
22130 => conv_std_logic_vector(38, 8),
22131 => conv_std_logic_vector(38, 8),
22132 => conv_std_logic_vector(38, 8),
22133 => conv_std_logic_vector(39, 8),
22134 => conv_std_logic_vector(39, 8),
22135 => conv_std_logic_vector(39, 8),
22136 => conv_std_logic_vector(40, 8),
22137 => conv_std_logic_vector(40, 8),
22138 => conv_std_logic_vector(40, 8),
22139 => conv_std_logic_vector(41, 8),
22140 => conv_std_logic_vector(41, 8),
22141 => conv_std_logic_vector(41, 8),
22142 => conv_std_logic_vector(42, 8),
22143 => conv_std_logic_vector(42, 8),
22144 => conv_std_logic_vector(43, 8),
22145 => conv_std_logic_vector(43, 8),
22146 => conv_std_logic_vector(43, 8),
22147 => conv_std_logic_vector(44, 8),
22148 => conv_std_logic_vector(44, 8),
22149 => conv_std_logic_vector(44, 8),
22150 => conv_std_logic_vector(45, 8),
22151 => conv_std_logic_vector(45, 8),
22152 => conv_std_logic_vector(45, 8),
22153 => conv_std_logic_vector(46, 8),
22154 => conv_std_logic_vector(46, 8),
22155 => conv_std_logic_vector(46, 8),
22156 => conv_std_logic_vector(47, 8),
22157 => conv_std_logic_vector(47, 8),
22158 => conv_std_logic_vector(47, 8),
22159 => conv_std_logic_vector(48, 8),
22160 => conv_std_logic_vector(48, 8),
22161 => conv_std_logic_vector(48, 8),
22162 => conv_std_logic_vector(49, 8),
22163 => conv_std_logic_vector(49, 8),
22164 => conv_std_logic_vector(49, 8),
22165 => conv_std_logic_vector(50, 8),
22166 => conv_std_logic_vector(50, 8),
22167 => conv_std_logic_vector(50, 8),
22168 => conv_std_logic_vector(51, 8),
22169 => conv_std_logic_vector(51, 8),
22170 => conv_std_logic_vector(51, 8),
22171 => conv_std_logic_vector(52, 8),
22172 => conv_std_logic_vector(52, 8),
22173 => conv_std_logic_vector(52, 8),
22174 => conv_std_logic_vector(53, 8),
22175 => conv_std_logic_vector(53, 8),
22176 => conv_std_logic_vector(53, 8),
22177 => conv_std_logic_vector(54, 8),
22178 => conv_std_logic_vector(54, 8),
22179 => conv_std_logic_vector(54, 8),
22180 => conv_std_logic_vector(55, 8),
22181 => conv_std_logic_vector(55, 8),
22182 => conv_std_logic_vector(55, 8),
22183 => conv_std_logic_vector(56, 8),
22184 => conv_std_logic_vector(56, 8),
22185 => conv_std_logic_vector(56, 8),
22186 => conv_std_logic_vector(57, 8),
22187 => conv_std_logic_vector(57, 8),
22188 => conv_std_logic_vector(57, 8),
22189 => conv_std_logic_vector(58, 8),
22190 => conv_std_logic_vector(58, 8),
22191 => conv_std_logic_vector(58, 8),
22192 => conv_std_logic_vector(59, 8),
22193 => conv_std_logic_vector(59, 8),
22194 => conv_std_logic_vector(59, 8),
22195 => conv_std_logic_vector(60, 8),
22196 => conv_std_logic_vector(60, 8),
22197 => conv_std_logic_vector(60, 8),
22198 => conv_std_logic_vector(61, 8),
22199 => conv_std_logic_vector(61, 8),
22200 => conv_std_logic_vector(61, 8),
22201 => conv_std_logic_vector(62, 8),
22202 => conv_std_logic_vector(62, 8),
22203 => conv_std_logic_vector(62, 8),
22204 => conv_std_logic_vector(63, 8),
22205 => conv_std_logic_vector(63, 8),
22206 => conv_std_logic_vector(63, 8),
22207 => conv_std_logic_vector(64, 8),
22208 => conv_std_logic_vector(64, 8),
22209 => conv_std_logic_vector(64, 8),
22210 => conv_std_logic_vector(65, 8),
22211 => conv_std_logic_vector(65, 8),
22212 => conv_std_logic_vector(65, 8),
22213 => conv_std_logic_vector(66, 8),
22214 => conv_std_logic_vector(66, 8),
22215 => conv_std_logic_vector(66, 8),
22216 => conv_std_logic_vector(67, 8),
22217 => conv_std_logic_vector(67, 8),
22218 => conv_std_logic_vector(67, 8),
22219 => conv_std_logic_vector(68, 8),
22220 => conv_std_logic_vector(68, 8),
22221 => conv_std_logic_vector(68, 8),
22222 => conv_std_logic_vector(69, 8),
22223 => conv_std_logic_vector(69, 8),
22224 => conv_std_logic_vector(69, 8),
22225 => conv_std_logic_vector(70, 8),
22226 => conv_std_logic_vector(70, 8),
22227 => conv_std_logic_vector(70, 8),
22228 => conv_std_logic_vector(71, 8),
22229 => conv_std_logic_vector(71, 8),
22230 => conv_std_logic_vector(71, 8),
22231 => conv_std_logic_vector(72, 8),
22232 => conv_std_logic_vector(72, 8),
22233 => conv_std_logic_vector(72, 8),
22234 => conv_std_logic_vector(73, 8),
22235 => conv_std_logic_vector(73, 8),
22236 => conv_std_logic_vector(73, 8),
22237 => conv_std_logic_vector(74, 8),
22238 => conv_std_logic_vector(74, 8),
22239 => conv_std_logic_vector(74, 8),
22240 => conv_std_logic_vector(75, 8),
22241 => conv_std_logic_vector(75, 8),
22242 => conv_std_logic_vector(75, 8),
22243 => conv_std_logic_vector(76, 8),
22244 => conv_std_logic_vector(76, 8),
22245 => conv_std_logic_vector(76, 8),
22246 => conv_std_logic_vector(77, 8),
22247 => conv_std_logic_vector(77, 8),
22248 => conv_std_logic_vector(77, 8),
22249 => conv_std_logic_vector(78, 8),
22250 => conv_std_logic_vector(78, 8),
22251 => conv_std_logic_vector(78, 8),
22252 => conv_std_logic_vector(79, 8),
22253 => conv_std_logic_vector(79, 8),
22254 => conv_std_logic_vector(79, 8),
22255 => conv_std_logic_vector(80, 8),
22256 => conv_std_logic_vector(80, 8),
22257 => conv_std_logic_vector(80, 8),
22258 => conv_std_logic_vector(81, 8),
22259 => conv_std_logic_vector(81, 8),
22260 => conv_std_logic_vector(81, 8),
22261 => conv_std_logic_vector(82, 8),
22262 => conv_std_logic_vector(82, 8),
22263 => conv_std_logic_vector(82, 8),
22264 => conv_std_logic_vector(83, 8),
22265 => conv_std_logic_vector(83, 8),
22266 => conv_std_logic_vector(83, 8),
22267 => conv_std_logic_vector(84, 8),
22268 => conv_std_logic_vector(84, 8),
22269 => conv_std_logic_vector(84, 8),
22270 => conv_std_logic_vector(85, 8),
22271 => conv_std_logic_vector(85, 8),
22272 => conv_std_logic_vector(0, 8),
22273 => conv_std_logic_vector(0, 8),
22274 => conv_std_logic_vector(0, 8),
22275 => conv_std_logic_vector(1, 8),
22276 => conv_std_logic_vector(1, 8),
22277 => conv_std_logic_vector(1, 8),
22278 => conv_std_logic_vector(2, 8),
22279 => conv_std_logic_vector(2, 8),
22280 => conv_std_logic_vector(2, 8),
22281 => conv_std_logic_vector(3, 8),
22282 => conv_std_logic_vector(3, 8),
22283 => conv_std_logic_vector(3, 8),
22284 => conv_std_logic_vector(4, 8),
22285 => conv_std_logic_vector(4, 8),
22286 => conv_std_logic_vector(4, 8),
22287 => conv_std_logic_vector(5, 8),
22288 => conv_std_logic_vector(5, 8),
22289 => conv_std_logic_vector(5, 8),
22290 => conv_std_logic_vector(6, 8),
22291 => conv_std_logic_vector(6, 8),
22292 => conv_std_logic_vector(6, 8),
22293 => conv_std_logic_vector(7, 8),
22294 => conv_std_logic_vector(7, 8),
22295 => conv_std_logic_vector(7, 8),
22296 => conv_std_logic_vector(8, 8),
22297 => conv_std_logic_vector(8, 8),
22298 => conv_std_logic_vector(8, 8),
22299 => conv_std_logic_vector(9, 8),
22300 => conv_std_logic_vector(9, 8),
22301 => conv_std_logic_vector(9, 8),
22302 => conv_std_logic_vector(10, 8),
22303 => conv_std_logic_vector(10, 8),
22304 => conv_std_logic_vector(10, 8),
22305 => conv_std_logic_vector(11, 8),
22306 => conv_std_logic_vector(11, 8),
22307 => conv_std_logic_vector(11, 8),
22308 => conv_std_logic_vector(12, 8),
22309 => conv_std_logic_vector(12, 8),
22310 => conv_std_logic_vector(12, 8),
22311 => conv_std_logic_vector(13, 8),
22312 => conv_std_logic_vector(13, 8),
22313 => conv_std_logic_vector(13, 8),
22314 => conv_std_logic_vector(14, 8),
22315 => conv_std_logic_vector(14, 8),
22316 => conv_std_logic_vector(14, 8),
22317 => conv_std_logic_vector(15, 8),
22318 => conv_std_logic_vector(15, 8),
22319 => conv_std_logic_vector(15, 8),
22320 => conv_std_logic_vector(16, 8),
22321 => conv_std_logic_vector(16, 8),
22322 => conv_std_logic_vector(16, 8),
22323 => conv_std_logic_vector(17, 8),
22324 => conv_std_logic_vector(17, 8),
22325 => conv_std_logic_vector(18, 8),
22326 => conv_std_logic_vector(18, 8),
22327 => conv_std_logic_vector(18, 8),
22328 => conv_std_logic_vector(19, 8),
22329 => conv_std_logic_vector(19, 8),
22330 => conv_std_logic_vector(19, 8),
22331 => conv_std_logic_vector(20, 8),
22332 => conv_std_logic_vector(20, 8),
22333 => conv_std_logic_vector(20, 8),
22334 => conv_std_logic_vector(21, 8),
22335 => conv_std_logic_vector(21, 8),
22336 => conv_std_logic_vector(21, 8),
22337 => conv_std_logic_vector(22, 8),
22338 => conv_std_logic_vector(22, 8),
22339 => conv_std_logic_vector(22, 8),
22340 => conv_std_logic_vector(23, 8),
22341 => conv_std_logic_vector(23, 8),
22342 => conv_std_logic_vector(23, 8),
22343 => conv_std_logic_vector(24, 8),
22344 => conv_std_logic_vector(24, 8),
22345 => conv_std_logic_vector(24, 8),
22346 => conv_std_logic_vector(25, 8),
22347 => conv_std_logic_vector(25, 8),
22348 => conv_std_logic_vector(25, 8),
22349 => conv_std_logic_vector(26, 8),
22350 => conv_std_logic_vector(26, 8),
22351 => conv_std_logic_vector(26, 8),
22352 => conv_std_logic_vector(27, 8),
22353 => conv_std_logic_vector(27, 8),
22354 => conv_std_logic_vector(27, 8),
22355 => conv_std_logic_vector(28, 8),
22356 => conv_std_logic_vector(28, 8),
22357 => conv_std_logic_vector(28, 8),
22358 => conv_std_logic_vector(29, 8),
22359 => conv_std_logic_vector(29, 8),
22360 => conv_std_logic_vector(29, 8),
22361 => conv_std_logic_vector(30, 8),
22362 => conv_std_logic_vector(30, 8),
22363 => conv_std_logic_vector(30, 8),
22364 => conv_std_logic_vector(31, 8),
22365 => conv_std_logic_vector(31, 8),
22366 => conv_std_logic_vector(31, 8),
22367 => conv_std_logic_vector(32, 8),
22368 => conv_std_logic_vector(32, 8),
22369 => conv_std_logic_vector(32, 8),
22370 => conv_std_logic_vector(33, 8),
22371 => conv_std_logic_vector(33, 8),
22372 => conv_std_logic_vector(33, 8),
22373 => conv_std_logic_vector(34, 8),
22374 => conv_std_logic_vector(34, 8),
22375 => conv_std_logic_vector(35, 8),
22376 => conv_std_logic_vector(35, 8),
22377 => conv_std_logic_vector(35, 8),
22378 => conv_std_logic_vector(36, 8),
22379 => conv_std_logic_vector(36, 8),
22380 => conv_std_logic_vector(36, 8),
22381 => conv_std_logic_vector(37, 8),
22382 => conv_std_logic_vector(37, 8),
22383 => conv_std_logic_vector(37, 8),
22384 => conv_std_logic_vector(38, 8),
22385 => conv_std_logic_vector(38, 8),
22386 => conv_std_logic_vector(38, 8),
22387 => conv_std_logic_vector(39, 8),
22388 => conv_std_logic_vector(39, 8),
22389 => conv_std_logic_vector(39, 8),
22390 => conv_std_logic_vector(40, 8),
22391 => conv_std_logic_vector(40, 8),
22392 => conv_std_logic_vector(40, 8),
22393 => conv_std_logic_vector(41, 8),
22394 => conv_std_logic_vector(41, 8),
22395 => conv_std_logic_vector(41, 8),
22396 => conv_std_logic_vector(42, 8),
22397 => conv_std_logic_vector(42, 8),
22398 => conv_std_logic_vector(42, 8),
22399 => conv_std_logic_vector(43, 8),
22400 => conv_std_logic_vector(43, 8),
22401 => conv_std_logic_vector(43, 8),
22402 => conv_std_logic_vector(44, 8),
22403 => conv_std_logic_vector(44, 8),
22404 => conv_std_logic_vector(44, 8),
22405 => conv_std_logic_vector(45, 8),
22406 => conv_std_logic_vector(45, 8),
22407 => conv_std_logic_vector(45, 8),
22408 => conv_std_logic_vector(46, 8),
22409 => conv_std_logic_vector(46, 8),
22410 => conv_std_logic_vector(46, 8),
22411 => conv_std_logic_vector(47, 8),
22412 => conv_std_logic_vector(47, 8),
22413 => conv_std_logic_vector(47, 8),
22414 => conv_std_logic_vector(48, 8),
22415 => conv_std_logic_vector(48, 8),
22416 => conv_std_logic_vector(48, 8),
22417 => conv_std_logic_vector(49, 8),
22418 => conv_std_logic_vector(49, 8),
22419 => conv_std_logic_vector(49, 8),
22420 => conv_std_logic_vector(50, 8),
22421 => conv_std_logic_vector(50, 8),
22422 => conv_std_logic_vector(50, 8),
22423 => conv_std_logic_vector(51, 8),
22424 => conv_std_logic_vector(51, 8),
22425 => conv_std_logic_vector(51, 8),
22426 => conv_std_logic_vector(52, 8),
22427 => conv_std_logic_vector(52, 8),
22428 => conv_std_logic_vector(53, 8),
22429 => conv_std_logic_vector(53, 8),
22430 => conv_std_logic_vector(53, 8),
22431 => conv_std_logic_vector(54, 8),
22432 => conv_std_logic_vector(54, 8),
22433 => conv_std_logic_vector(54, 8),
22434 => conv_std_logic_vector(55, 8),
22435 => conv_std_logic_vector(55, 8),
22436 => conv_std_logic_vector(55, 8),
22437 => conv_std_logic_vector(56, 8),
22438 => conv_std_logic_vector(56, 8),
22439 => conv_std_logic_vector(56, 8),
22440 => conv_std_logic_vector(57, 8),
22441 => conv_std_logic_vector(57, 8),
22442 => conv_std_logic_vector(57, 8),
22443 => conv_std_logic_vector(58, 8),
22444 => conv_std_logic_vector(58, 8),
22445 => conv_std_logic_vector(58, 8),
22446 => conv_std_logic_vector(59, 8),
22447 => conv_std_logic_vector(59, 8),
22448 => conv_std_logic_vector(59, 8),
22449 => conv_std_logic_vector(60, 8),
22450 => conv_std_logic_vector(60, 8),
22451 => conv_std_logic_vector(60, 8),
22452 => conv_std_logic_vector(61, 8),
22453 => conv_std_logic_vector(61, 8),
22454 => conv_std_logic_vector(61, 8),
22455 => conv_std_logic_vector(62, 8),
22456 => conv_std_logic_vector(62, 8),
22457 => conv_std_logic_vector(62, 8),
22458 => conv_std_logic_vector(63, 8),
22459 => conv_std_logic_vector(63, 8),
22460 => conv_std_logic_vector(63, 8),
22461 => conv_std_logic_vector(64, 8),
22462 => conv_std_logic_vector(64, 8),
22463 => conv_std_logic_vector(64, 8),
22464 => conv_std_logic_vector(65, 8),
22465 => conv_std_logic_vector(65, 8),
22466 => conv_std_logic_vector(65, 8),
22467 => conv_std_logic_vector(66, 8),
22468 => conv_std_logic_vector(66, 8),
22469 => conv_std_logic_vector(66, 8),
22470 => conv_std_logic_vector(67, 8),
22471 => conv_std_logic_vector(67, 8),
22472 => conv_std_logic_vector(67, 8),
22473 => conv_std_logic_vector(68, 8),
22474 => conv_std_logic_vector(68, 8),
22475 => conv_std_logic_vector(68, 8),
22476 => conv_std_logic_vector(69, 8),
22477 => conv_std_logic_vector(69, 8),
22478 => conv_std_logic_vector(70, 8),
22479 => conv_std_logic_vector(70, 8),
22480 => conv_std_logic_vector(70, 8),
22481 => conv_std_logic_vector(71, 8),
22482 => conv_std_logic_vector(71, 8),
22483 => conv_std_logic_vector(71, 8),
22484 => conv_std_logic_vector(72, 8),
22485 => conv_std_logic_vector(72, 8),
22486 => conv_std_logic_vector(72, 8),
22487 => conv_std_logic_vector(73, 8),
22488 => conv_std_logic_vector(73, 8),
22489 => conv_std_logic_vector(73, 8),
22490 => conv_std_logic_vector(74, 8),
22491 => conv_std_logic_vector(74, 8),
22492 => conv_std_logic_vector(74, 8),
22493 => conv_std_logic_vector(75, 8),
22494 => conv_std_logic_vector(75, 8),
22495 => conv_std_logic_vector(75, 8),
22496 => conv_std_logic_vector(76, 8),
22497 => conv_std_logic_vector(76, 8),
22498 => conv_std_logic_vector(76, 8),
22499 => conv_std_logic_vector(77, 8),
22500 => conv_std_logic_vector(77, 8),
22501 => conv_std_logic_vector(77, 8),
22502 => conv_std_logic_vector(78, 8),
22503 => conv_std_logic_vector(78, 8),
22504 => conv_std_logic_vector(78, 8),
22505 => conv_std_logic_vector(79, 8),
22506 => conv_std_logic_vector(79, 8),
22507 => conv_std_logic_vector(79, 8),
22508 => conv_std_logic_vector(80, 8),
22509 => conv_std_logic_vector(80, 8),
22510 => conv_std_logic_vector(80, 8),
22511 => conv_std_logic_vector(81, 8),
22512 => conv_std_logic_vector(81, 8),
22513 => conv_std_logic_vector(81, 8),
22514 => conv_std_logic_vector(82, 8),
22515 => conv_std_logic_vector(82, 8),
22516 => conv_std_logic_vector(82, 8),
22517 => conv_std_logic_vector(83, 8),
22518 => conv_std_logic_vector(83, 8),
22519 => conv_std_logic_vector(83, 8),
22520 => conv_std_logic_vector(84, 8),
22521 => conv_std_logic_vector(84, 8),
22522 => conv_std_logic_vector(84, 8),
22523 => conv_std_logic_vector(85, 8),
22524 => conv_std_logic_vector(85, 8),
22525 => conv_std_logic_vector(85, 8),
22526 => conv_std_logic_vector(86, 8),
22527 => conv_std_logic_vector(86, 8),
22528 => conv_std_logic_vector(0, 8),
22529 => conv_std_logic_vector(0, 8),
22530 => conv_std_logic_vector(0, 8),
22531 => conv_std_logic_vector(1, 8),
22532 => conv_std_logic_vector(1, 8),
22533 => conv_std_logic_vector(1, 8),
22534 => conv_std_logic_vector(2, 8),
22535 => conv_std_logic_vector(2, 8),
22536 => conv_std_logic_vector(2, 8),
22537 => conv_std_logic_vector(3, 8),
22538 => conv_std_logic_vector(3, 8),
22539 => conv_std_logic_vector(3, 8),
22540 => conv_std_logic_vector(4, 8),
22541 => conv_std_logic_vector(4, 8),
22542 => conv_std_logic_vector(4, 8),
22543 => conv_std_logic_vector(5, 8),
22544 => conv_std_logic_vector(5, 8),
22545 => conv_std_logic_vector(5, 8),
22546 => conv_std_logic_vector(6, 8),
22547 => conv_std_logic_vector(6, 8),
22548 => conv_std_logic_vector(6, 8),
22549 => conv_std_logic_vector(7, 8),
22550 => conv_std_logic_vector(7, 8),
22551 => conv_std_logic_vector(7, 8),
22552 => conv_std_logic_vector(8, 8),
22553 => conv_std_logic_vector(8, 8),
22554 => conv_std_logic_vector(8, 8),
22555 => conv_std_logic_vector(9, 8),
22556 => conv_std_logic_vector(9, 8),
22557 => conv_std_logic_vector(9, 8),
22558 => conv_std_logic_vector(10, 8),
22559 => conv_std_logic_vector(10, 8),
22560 => conv_std_logic_vector(11, 8),
22561 => conv_std_logic_vector(11, 8),
22562 => conv_std_logic_vector(11, 8),
22563 => conv_std_logic_vector(12, 8),
22564 => conv_std_logic_vector(12, 8),
22565 => conv_std_logic_vector(12, 8),
22566 => conv_std_logic_vector(13, 8),
22567 => conv_std_logic_vector(13, 8),
22568 => conv_std_logic_vector(13, 8),
22569 => conv_std_logic_vector(14, 8),
22570 => conv_std_logic_vector(14, 8),
22571 => conv_std_logic_vector(14, 8),
22572 => conv_std_logic_vector(15, 8),
22573 => conv_std_logic_vector(15, 8),
22574 => conv_std_logic_vector(15, 8),
22575 => conv_std_logic_vector(16, 8),
22576 => conv_std_logic_vector(16, 8),
22577 => conv_std_logic_vector(16, 8),
22578 => conv_std_logic_vector(17, 8),
22579 => conv_std_logic_vector(17, 8),
22580 => conv_std_logic_vector(17, 8),
22581 => conv_std_logic_vector(18, 8),
22582 => conv_std_logic_vector(18, 8),
22583 => conv_std_logic_vector(18, 8),
22584 => conv_std_logic_vector(19, 8),
22585 => conv_std_logic_vector(19, 8),
22586 => conv_std_logic_vector(19, 8),
22587 => conv_std_logic_vector(20, 8),
22588 => conv_std_logic_vector(20, 8),
22589 => conv_std_logic_vector(20, 8),
22590 => conv_std_logic_vector(21, 8),
22591 => conv_std_logic_vector(21, 8),
22592 => conv_std_logic_vector(22, 8),
22593 => conv_std_logic_vector(22, 8),
22594 => conv_std_logic_vector(22, 8),
22595 => conv_std_logic_vector(23, 8),
22596 => conv_std_logic_vector(23, 8),
22597 => conv_std_logic_vector(23, 8),
22598 => conv_std_logic_vector(24, 8),
22599 => conv_std_logic_vector(24, 8),
22600 => conv_std_logic_vector(24, 8),
22601 => conv_std_logic_vector(25, 8),
22602 => conv_std_logic_vector(25, 8),
22603 => conv_std_logic_vector(25, 8),
22604 => conv_std_logic_vector(26, 8),
22605 => conv_std_logic_vector(26, 8),
22606 => conv_std_logic_vector(26, 8),
22607 => conv_std_logic_vector(27, 8),
22608 => conv_std_logic_vector(27, 8),
22609 => conv_std_logic_vector(27, 8),
22610 => conv_std_logic_vector(28, 8),
22611 => conv_std_logic_vector(28, 8),
22612 => conv_std_logic_vector(28, 8),
22613 => conv_std_logic_vector(29, 8),
22614 => conv_std_logic_vector(29, 8),
22615 => conv_std_logic_vector(29, 8),
22616 => conv_std_logic_vector(30, 8),
22617 => conv_std_logic_vector(30, 8),
22618 => conv_std_logic_vector(30, 8),
22619 => conv_std_logic_vector(31, 8),
22620 => conv_std_logic_vector(31, 8),
22621 => conv_std_logic_vector(31, 8),
22622 => conv_std_logic_vector(32, 8),
22623 => conv_std_logic_vector(32, 8),
22624 => conv_std_logic_vector(33, 8),
22625 => conv_std_logic_vector(33, 8),
22626 => conv_std_logic_vector(33, 8),
22627 => conv_std_logic_vector(34, 8),
22628 => conv_std_logic_vector(34, 8),
22629 => conv_std_logic_vector(34, 8),
22630 => conv_std_logic_vector(35, 8),
22631 => conv_std_logic_vector(35, 8),
22632 => conv_std_logic_vector(35, 8),
22633 => conv_std_logic_vector(36, 8),
22634 => conv_std_logic_vector(36, 8),
22635 => conv_std_logic_vector(36, 8),
22636 => conv_std_logic_vector(37, 8),
22637 => conv_std_logic_vector(37, 8),
22638 => conv_std_logic_vector(37, 8),
22639 => conv_std_logic_vector(38, 8),
22640 => conv_std_logic_vector(38, 8),
22641 => conv_std_logic_vector(38, 8),
22642 => conv_std_logic_vector(39, 8),
22643 => conv_std_logic_vector(39, 8),
22644 => conv_std_logic_vector(39, 8),
22645 => conv_std_logic_vector(40, 8),
22646 => conv_std_logic_vector(40, 8),
22647 => conv_std_logic_vector(40, 8),
22648 => conv_std_logic_vector(41, 8),
22649 => conv_std_logic_vector(41, 8),
22650 => conv_std_logic_vector(41, 8),
22651 => conv_std_logic_vector(42, 8),
22652 => conv_std_logic_vector(42, 8),
22653 => conv_std_logic_vector(42, 8),
22654 => conv_std_logic_vector(43, 8),
22655 => conv_std_logic_vector(43, 8),
22656 => conv_std_logic_vector(44, 8),
22657 => conv_std_logic_vector(44, 8),
22658 => conv_std_logic_vector(44, 8),
22659 => conv_std_logic_vector(45, 8),
22660 => conv_std_logic_vector(45, 8),
22661 => conv_std_logic_vector(45, 8),
22662 => conv_std_logic_vector(46, 8),
22663 => conv_std_logic_vector(46, 8),
22664 => conv_std_logic_vector(46, 8),
22665 => conv_std_logic_vector(47, 8),
22666 => conv_std_logic_vector(47, 8),
22667 => conv_std_logic_vector(47, 8),
22668 => conv_std_logic_vector(48, 8),
22669 => conv_std_logic_vector(48, 8),
22670 => conv_std_logic_vector(48, 8),
22671 => conv_std_logic_vector(49, 8),
22672 => conv_std_logic_vector(49, 8),
22673 => conv_std_logic_vector(49, 8),
22674 => conv_std_logic_vector(50, 8),
22675 => conv_std_logic_vector(50, 8),
22676 => conv_std_logic_vector(50, 8),
22677 => conv_std_logic_vector(51, 8),
22678 => conv_std_logic_vector(51, 8),
22679 => conv_std_logic_vector(51, 8),
22680 => conv_std_logic_vector(52, 8),
22681 => conv_std_logic_vector(52, 8),
22682 => conv_std_logic_vector(52, 8),
22683 => conv_std_logic_vector(53, 8),
22684 => conv_std_logic_vector(53, 8),
22685 => conv_std_logic_vector(53, 8),
22686 => conv_std_logic_vector(54, 8),
22687 => conv_std_logic_vector(54, 8),
22688 => conv_std_logic_vector(55, 8),
22689 => conv_std_logic_vector(55, 8),
22690 => conv_std_logic_vector(55, 8),
22691 => conv_std_logic_vector(56, 8),
22692 => conv_std_logic_vector(56, 8),
22693 => conv_std_logic_vector(56, 8),
22694 => conv_std_logic_vector(57, 8),
22695 => conv_std_logic_vector(57, 8),
22696 => conv_std_logic_vector(57, 8),
22697 => conv_std_logic_vector(58, 8),
22698 => conv_std_logic_vector(58, 8),
22699 => conv_std_logic_vector(58, 8),
22700 => conv_std_logic_vector(59, 8),
22701 => conv_std_logic_vector(59, 8),
22702 => conv_std_logic_vector(59, 8),
22703 => conv_std_logic_vector(60, 8),
22704 => conv_std_logic_vector(60, 8),
22705 => conv_std_logic_vector(60, 8),
22706 => conv_std_logic_vector(61, 8),
22707 => conv_std_logic_vector(61, 8),
22708 => conv_std_logic_vector(61, 8),
22709 => conv_std_logic_vector(62, 8),
22710 => conv_std_logic_vector(62, 8),
22711 => conv_std_logic_vector(62, 8),
22712 => conv_std_logic_vector(63, 8),
22713 => conv_std_logic_vector(63, 8),
22714 => conv_std_logic_vector(63, 8),
22715 => conv_std_logic_vector(64, 8),
22716 => conv_std_logic_vector(64, 8),
22717 => conv_std_logic_vector(64, 8),
22718 => conv_std_logic_vector(65, 8),
22719 => conv_std_logic_vector(65, 8),
22720 => conv_std_logic_vector(66, 8),
22721 => conv_std_logic_vector(66, 8),
22722 => conv_std_logic_vector(66, 8),
22723 => conv_std_logic_vector(67, 8),
22724 => conv_std_logic_vector(67, 8),
22725 => conv_std_logic_vector(67, 8),
22726 => conv_std_logic_vector(68, 8),
22727 => conv_std_logic_vector(68, 8),
22728 => conv_std_logic_vector(68, 8),
22729 => conv_std_logic_vector(69, 8),
22730 => conv_std_logic_vector(69, 8),
22731 => conv_std_logic_vector(69, 8),
22732 => conv_std_logic_vector(70, 8),
22733 => conv_std_logic_vector(70, 8),
22734 => conv_std_logic_vector(70, 8),
22735 => conv_std_logic_vector(71, 8),
22736 => conv_std_logic_vector(71, 8),
22737 => conv_std_logic_vector(71, 8),
22738 => conv_std_logic_vector(72, 8),
22739 => conv_std_logic_vector(72, 8),
22740 => conv_std_logic_vector(72, 8),
22741 => conv_std_logic_vector(73, 8),
22742 => conv_std_logic_vector(73, 8),
22743 => conv_std_logic_vector(73, 8),
22744 => conv_std_logic_vector(74, 8),
22745 => conv_std_logic_vector(74, 8),
22746 => conv_std_logic_vector(74, 8),
22747 => conv_std_logic_vector(75, 8),
22748 => conv_std_logic_vector(75, 8),
22749 => conv_std_logic_vector(75, 8),
22750 => conv_std_logic_vector(76, 8),
22751 => conv_std_logic_vector(76, 8),
22752 => conv_std_logic_vector(77, 8),
22753 => conv_std_logic_vector(77, 8),
22754 => conv_std_logic_vector(77, 8),
22755 => conv_std_logic_vector(78, 8),
22756 => conv_std_logic_vector(78, 8),
22757 => conv_std_logic_vector(78, 8),
22758 => conv_std_logic_vector(79, 8),
22759 => conv_std_logic_vector(79, 8),
22760 => conv_std_logic_vector(79, 8),
22761 => conv_std_logic_vector(80, 8),
22762 => conv_std_logic_vector(80, 8),
22763 => conv_std_logic_vector(80, 8),
22764 => conv_std_logic_vector(81, 8),
22765 => conv_std_logic_vector(81, 8),
22766 => conv_std_logic_vector(81, 8),
22767 => conv_std_logic_vector(82, 8),
22768 => conv_std_logic_vector(82, 8),
22769 => conv_std_logic_vector(82, 8),
22770 => conv_std_logic_vector(83, 8),
22771 => conv_std_logic_vector(83, 8),
22772 => conv_std_logic_vector(83, 8),
22773 => conv_std_logic_vector(84, 8),
22774 => conv_std_logic_vector(84, 8),
22775 => conv_std_logic_vector(84, 8),
22776 => conv_std_logic_vector(85, 8),
22777 => conv_std_logic_vector(85, 8),
22778 => conv_std_logic_vector(85, 8),
22779 => conv_std_logic_vector(86, 8),
22780 => conv_std_logic_vector(86, 8),
22781 => conv_std_logic_vector(86, 8),
22782 => conv_std_logic_vector(87, 8),
22783 => conv_std_logic_vector(87, 8),
22784 => conv_std_logic_vector(0, 8),
22785 => conv_std_logic_vector(0, 8),
22786 => conv_std_logic_vector(0, 8),
22787 => conv_std_logic_vector(1, 8),
22788 => conv_std_logic_vector(1, 8),
22789 => conv_std_logic_vector(1, 8),
22790 => conv_std_logic_vector(2, 8),
22791 => conv_std_logic_vector(2, 8),
22792 => conv_std_logic_vector(2, 8),
22793 => conv_std_logic_vector(3, 8),
22794 => conv_std_logic_vector(3, 8),
22795 => conv_std_logic_vector(3, 8),
22796 => conv_std_logic_vector(4, 8),
22797 => conv_std_logic_vector(4, 8),
22798 => conv_std_logic_vector(4, 8),
22799 => conv_std_logic_vector(5, 8),
22800 => conv_std_logic_vector(5, 8),
22801 => conv_std_logic_vector(5, 8),
22802 => conv_std_logic_vector(6, 8),
22803 => conv_std_logic_vector(6, 8),
22804 => conv_std_logic_vector(6, 8),
22805 => conv_std_logic_vector(7, 8),
22806 => conv_std_logic_vector(7, 8),
22807 => conv_std_logic_vector(7, 8),
22808 => conv_std_logic_vector(8, 8),
22809 => conv_std_logic_vector(8, 8),
22810 => conv_std_logic_vector(9, 8),
22811 => conv_std_logic_vector(9, 8),
22812 => conv_std_logic_vector(9, 8),
22813 => conv_std_logic_vector(10, 8),
22814 => conv_std_logic_vector(10, 8),
22815 => conv_std_logic_vector(10, 8),
22816 => conv_std_logic_vector(11, 8),
22817 => conv_std_logic_vector(11, 8),
22818 => conv_std_logic_vector(11, 8),
22819 => conv_std_logic_vector(12, 8),
22820 => conv_std_logic_vector(12, 8),
22821 => conv_std_logic_vector(12, 8),
22822 => conv_std_logic_vector(13, 8),
22823 => conv_std_logic_vector(13, 8),
22824 => conv_std_logic_vector(13, 8),
22825 => conv_std_logic_vector(14, 8),
22826 => conv_std_logic_vector(14, 8),
22827 => conv_std_logic_vector(14, 8),
22828 => conv_std_logic_vector(15, 8),
22829 => conv_std_logic_vector(15, 8),
22830 => conv_std_logic_vector(15, 8),
22831 => conv_std_logic_vector(16, 8),
22832 => conv_std_logic_vector(16, 8),
22833 => conv_std_logic_vector(17, 8),
22834 => conv_std_logic_vector(17, 8),
22835 => conv_std_logic_vector(17, 8),
22836 => conv_std_logic_vector(18, 8),
22837 => conv_std_logic_vector(18, 8),
22838 => conv_std_logic_vector(18, 8),
22839 => conv_std_logic_vector(19, 8),
22840 => conv_std_logic_vector(19, 8),
22841 => conv_std_logic_vector(19, 8),
22842 => conv_std_logic_vector(20, 8),
22843 => conv_std_logic_vector(20, 8),
22844 => conv_std_logic_vector(20, 8),
22845 => conv_std_logic_vector(21, 8),
22846 => conv_std_logic_vector(21, 8),
22847 => conv_std_logic_vector(21, 8),
22848 => conv_std_logic_vector(22, 8),
22849 => conv_std_logic_vector(22, 8),
22850 => conv_std_logic_vector(22, 8),
22851 => conv_std_logic_vector(23, 8),
22852 => conv_std_logic_vector(23, 8),
22853 => conv_std_logic_vector(23, 8),
22854 => conv_std_logic_vector(24, 8),
22855 => conv_std_logic_vector(24, 8),
22856 => conv_std_logic_vector(25, 8),
22857 => conv_std_logic_vector(25, 8),
22858 => conv_std_logic_vector(25, 8),
22859 => conv_std_logic_vector(26, 8),
22860 => conv_std_logic_vector(26, 8),
22861 => conv_std_logic_vector(26, 8),
22862 => conv_std_logic_vector(27, 8),
22863 => conv_std_logic_vector(27, 8),
22864 => conv_std_logic_vector(27, 8),
22865 => conv_std_logic_vector(28, 8),
22866 => conv_std_logic_vector(28, 8),
22867 => conv_std_logic_vector(28, 8),
22868 => conv_std_logic_vector(29, 8),
22869 => conv_std_logic_vector(29, 8),
22870 => conv_std_logic_vector(29, 8),
22871 => conv_std_logic_vector(30, 8),
22872 => conv_std_logic_vector(30, 8),
22873 => conv_std_logic_vector(30, 8),
22874 => conv_std_logic_vector(31, 8),
22875 => conv_std_logic_vector(31, 8),
22876 => conv_std_logic_vector(31, 8),
22877 => conv_std_logic_vector(32, 8),
22878 => conv_std_logic_vector(32, 8),
22879 => conv_std_logic_vector(33, 8),
22880 => conv_std_logic_vector(33, 8),
22881 => conv_std_logic_vector(33, 8),
22882 => conv_std_logic_vector(34, 8),
22883 => conv_std_logic_vector(34, 8),
22884 => conv_std_logic_vector(34, 8),
22885 => conv_std_logic_vector(35, 8),
22886 => conv_std_logic_vector(35, 8),
22887 => conv_std_logic_vector(35, 8),
22888 => conv_std_logic_vector(36, 8),
22889 => conv_std_logic_vector(36, 8),
22890 => conv_std_logic_vector(36, 8),
22891 => conv_std_logic_vector(37, 8),
22892 => conv_std_logic_vector(37, 8),
22893 => conv_std_logic_vector(37, 8),
22894 => conv_std_logic_vector(38, 8),
22895 => conv_std_logic_vector(38, 8),
22896 => conv_std_logic_vector(38, 8),
22897 => conv_std_logic_vector(39, 8),
22898 => conv_std_logic_vector(39, 8),
22899 => conv_std_logic_vector(39, 8),
22900 => conv_std_logic_vector(40, 8),
22901 => conv_std_logic_vector(40, 8),
22902 => conv_std_logic_vector(41, 8),
22903 => conv_std_logic_vector(41, 8),
22904 => conv_std_logic_vector(41, 8),
22905 => conv_std_logic_vector(42, 8),
22906 => conv_std_logic_vector(42, 8),
22907 => conv_std_logic_vector(42, 8),
22908 => conv_std_logic_vector(43, 8),
22909 => conv_std_logic_vector(43, 8),
22910 => conv_std_logic_vector(43, 8),
22911 => conv_std_logic_vector(44, 8),
22912 => conv_std_logic_vector(44, 8),
22913 => conv_std_logic_vector(44, 8),
22914 => conv_std_logic_vector(45, 8),
22915 => conv_std_logic_vector(45, 8),
22916 => conv_std_logic_vector(45, 8),
22917 => conv_std_logic_vector(46, 8),
22918 => conv_std_logic_vector(46, 8),
22919 => conv_std_logic_vector(46, 8),
22920 => conv_std_logic_vector(47, 8),
22921 => conv_std_logic_vector(47, 8),
22922 => conv_std_logic_vector(47, 8),
22923 => conv_std_logic_vector(48, 8),
22924 => conv_std_logic_vector(48, 8),
22925 => conv_std_logic_vector(49, 8),
22926 => conv_std_logic_vector(49, 8),
22927 => conv_std_logic_vector(49, 8),
22928 => conv_std_logic_vector(50, 8),
22929 => conv_std_logic_vector(50, 8),
22930 => conv_std_logic_vector(50, 8),
22931 => conv_std_logic_vector(51, 8),
22932 => conv_std_logic_vector(51, 8),
22933 => conv_std_logic_vector(51, 8),
22934 => conv_std_logic_vector(52, 8),
22935 => conv_std_logic_vector(52, 8),
22936 => conv_std_logic_vector(52, 8),
22937 => conv_std_logic_vector(53, 8),
22938 => conv_std_logic_vector(53, 8),
22939 => conv_std_logic_vector(53, 8),
22940 => conv_std_logic_vector(54, 8),
22941 => conv_std_logic_vector(54, 8),
22942 => conv_std_logic_vector(54, 8),
22943 => conv_std_logic_vector(55, 8),
22944 => conv_std_logic_vector(55, 8),
22945 => conv_std_logic_vector(55, 8),
22946 => conv_std_logic_vector(56, 8),
22947 => conv_std_logic_vector(56, 8),
22948 => conv_std_logic_vector(57, 8),
22949 => conv_std_logic_vector(57, 8),
22950 => conv_std_logic_vector(57, 8),
22951 => conv_std_logic_vector(58, 8),
22952 => conv_std_logic_vector(58, 8),
22953 => conv_std_logic_vector(58, 8),
22954 => conv_std_logic_vector(59, 8),
22955 => conv_std_logic_vector(59, 8),
22956 => conv_std_logic_vector(59, 8),
22957 => conv_std_logic_vector(60, 8),
22958 => conv_std_logic_vector(60, 8),
22959 => conv_std_logic_vector(60, 8),
22960 => conv_std_logic_vector(61, 8),
22961 => conv_std_logic_vector(61, 8),
22962 => conv_std_logic_vector(61, 8),
22963 => conv_std_logic_vector(62, 8),
22964 => conv_std_logic_vector(62, 8),
22965 => conv_std_logic_vector(62, 8),
22966 => conv_std_logic_vector(63, 8),
22967 => conv_std_logic_vector(63, 8),
22968 => conv_std_logic_vector(63, 8),
22969 => conv_std_logic_vector(64, 8),
22970 => conv_std_logic_vector(64, 8),
22971 => conv_std_logic_vector(65, 8),
22972 => conv_std_logic_vector(65, 8),
22973 => conv_std_logic_vector(65, 8),
22974 => conv_std_logic_vector(66, 8),
22975 => conv_std_logic_vector(66, 8),
22976 => conv_std_logic_vector(66, 8),
22977 => conv_std_logic_vector(67, 8),
22978 => conv_std_logic_vector(67, 8),
22979 => conv_std_logic_vector(67, 8),
22980 => conv_std_logic_vector(68, 8),
22981 => conv_std_logic_vector(68, 8),
22982 => conv_std_logic_vector(68, 8),
22983 => conv_std_logic_vector(69, 8),
22984 => conv_std_logic_vector(69, 8),
22985 => conv_std_logic_vector(69, 8),
22986 => conv_std_logic_vector(70, 8),
22987 => conv_std_logic_vector(70, 8),
22988 => conv_std_logic_vector(70, 8),
22989 => conv_std_logic_vector(71, 8),
22990 => conv_std_logic_vector(71, 8),
22991 => conv_std_logic_vector(71, 8),
22992 => conv_std_logic_vector(72, 8),
22993 => conv_std_logic_vector(72, 8),
22994 => conv_std_logic_vector(73, 8),
22995 => conv_std_logic_vector(73, 8),
22996 => conv_std_logic_vector(73, 8),
22997 => conv_std_logic_vector(74, 8),
22998 => conv_std_logic_vector(74, 8),
22999 => conv_std_logic_vector(74, 8),
23000 => conv_std_logic_vector(75, 8),
23001 => conv_std_logic_vector(75, 8),
23002 => conv_std_logic_vector(75, 8),
23003 => conv_std_logic_vector(76, 8),
23004 => conv_std_logic_vector(76, 8),
23005 => conv_std_logic_vector(76, 8),
23006 => conv_std_logic_vector(77, 8),
23007 => conv_std_logic_vector(77, 8),
23008 => conv_std_logic_vector(77, 8),
23009 => conv_std_logic_vector(78, 8),
23010 => conv_std_logic_vector(78, 8),
23011 => conv_std_logic_vector(78, 8),
23012 => conv_std_logic_vector(79, 8),
23013 => conv_std_logic_vector(79, 8),
23014 => conv_std_logic_vector(79, 8),
23015 => conv_std_logic_vector(80, 8),
23016 => conv_std_logic_vector(80, 8),
23017 => conv_std_logic_vector(81, 8),
23018 => conv_std_logic_vector(81, 8),
23019 => conv_std_logic_vector(81, 8),
23020 => conv_std_logic_vector(82, 8),
23021 => conv_std_logic_vector(82, 8),
23022 => conv_std_logic_vector(82, 8),
23023 => conv_std_logic_vector(83, 8),
23024 => conv_std_logic_vector(83, 8),
23025 => conv_std_logic_vector(83, 8),
23026 => conv_std_logic_vector(84, 8),
23027 => conv_std_logic_vector(84, 8),
23028 => conv_std_logic_vector(84, 8),
23029 => conv_std_logic_vector(85, 8),
23030 => conv_std_logic_vector(85, 8),
23031 => conv_std_logic_vector(85, 8),
23032 => conv_std_logic_vector(86, 8),
23033 => conv_std_logic_vector(86, 8),
23034 => conv_std_logic_vector(86, 8),
23035 => conv_std_logic_vector(87, 8),
23036 => conv_std_logic_vector(87, 8),
23037 => conv_std_logic_vector(87, 8),
23038 => conv_std_logic_vector(88, 8),
23039 => conv_std_logic_vector(88, 8),
23040 => conv_std_logic_vector(0, 8),
23041 => conv_std_logic_vector(0, 8),
23042 => conv_std_logic_vector(0, 8),
23043 => conv_std_logic_vector(1, 8),
23044 => conv_std_logic_vector(1, 8),
23045 => conv_std_logic_vector(1, 8),
23046 => conv_std_logic_vector(2, 8),
23047 => conv_std_logic_vector(2, 8),
23048 => conv_std_logic_vector(2, 8),
23049 => conv_std_logic_vector(3, 8),
23050 => conv_std_logic_vector(3, 8),
23051 => conv_std_logic_vector(3, 8),
23052 => conv_std_logic_vector(4, 8),
23053 => conv_std_logic_vector(4, 8),
23054 => conv_std_logic_vector(4, 8),
23055 => conv_std_logic_vector(5, 8),
23056 => conv_std_logic_vector(5, 8),
23057 => conv_std_logic_vector(5, 8),
23058 => conv_std_logic_vector(6, 8),
23059 => conv_std_logic_vector(6, 8),
23060 => conv_std_logic_vector(7, 8),
23061 => conv_std_logic_vector(7, 8),
23062 => conv_std_logic_vector(7, 8),
23063 => conv_std_logic_vector(8, 8),
23064 => conv_std_logic_vector(8, 8),
23065 => conv_std_logic_vector(8, 8),
23066 => conv_std_logic_vector(9, 8),
23067 => conv_std_logic_vector(9, 8),
23068 => conv_std_logic_vector(9, 8),
23069 => conv_std_logic_vector(10, 8),
23070 => conv_std_logic_vector(10, 8),
23071 => conv_std_logic_vector(10, 8),
23072 => conv_std_logic_vector(11, 8),
23073 => conv_std_logic_vector(11, 8),
23074 => conv_std_logic_vector(11, 8),
23075 => conv_std_logic_vector(12, 8),
23076 => conv_std_logic_vector(12, 8),
23077 => conv_std_logic_vector(13, 8),
23078 => conv_std_logic_vector(13, 8),
23079 => conv_std_logic_vector(13, 8),
23080 => conv_std_logic_vector(14, 8),
23081 => conv_std_logic_vector(14, 8),
23082 => conv_std_logic_vector(14, 8),
23083 => conv_std_logic_vector(15, 8),
23084 => conv_std_logic_vector(15, 8),
23085 => conv_std_logic_vector(15, 8),
23086 => conv_std_logic_vector(16, 8),
23087 => conv_std_logic_vector(16, 8),
23088 => conv_std_logic_vector(16, 8),
23089 => conv_std_logic_vector(17, 8),
23090 => conv_std_logic_vector(17, 8),
23091 => conv_std_logic_vector(17, 8),
23092 => conv_std_logic_vector(18, 8),
23093 => conv_std_logic_vector(18, 8),
23094 => conv_std_logic_vector(18, 8),
23095 => conv_std_logic_vector(19, 8),
23096 => conv_std_logic_vector(19, 8),
23097 => conv_std_logic_vector(20, 8),
23098 => conv_std_logic_vector(20, 8),
23099 => conv_std_logic_vector(20, 8),
23100 => conv_std_logic_vector(21, 8),
23101 => conv_std_logic_vector(21, 8),
23102 => conv_std_logic_vector(21, 8),
23103 => conv_std_logic_vector(22, 8),
23104 => conv_std_logic_vector(22, 8),
23105 => conv_std_logic_vector(22, 8),
23106 => conv_std_logic_vector(23, 8),
23107 => conv_std_logic_vector(23, 8),
23108 => conv_std_logic_vector(23, 8),
23109 => conv_std_logic_vector(24, 8),
23110 => conv_std_logic_vector(24, 8),
23111 => conv_std_logic_vector(24, 8),
23112 => conv_std_logic_vector(25, 8),
23113 => conv_std_logic_vector(25, 8),
23114 => conv_std_logic_vector(26, 8),
23115 => conv_std_logic_vector(26, 8),
23116 => conv_std_logic_vector(26, 8),
23117 => conv_std_logic_vector(27, 8),
23118 => conv_std_logic_vector(27, 8),
23119 => conv_std_logic_vector(27, 8),
23120 => conv_std_logic_vector(28, 8),
23121 => conv_std_logic_vector(28, 8),
23122 => conv_std_logic_vector(28, 8),
23123 => conv_std_logic_vector(29, 8),
23124 => conv_std_logic_vector(29, 8),
23125 => conv_std_logic_vector(29, 8),
23126 => conv_std_logic_vector(30, 8),
23127 => conv_std_logic_vector(30, 8),
23128 => conv_std_logic_vector(30, 8),
23129 => conv_std_logic_vector(31, 8),
23130 => conv_std_logic_vector(31, 8),
23131 => conv_std_logic_vector(31, 8),
23132 => conv_std_logic_vector(32, 8),
23133 => conv_std_logic_vector(32, 8),
23134 => conv_std_logic_vector(33, 8),
23135 => conv_std_logic_vector(33, 8),
23136 => conv_std_logic_vector(33, 8),
23137 => conv_std_logic_vector(34, 8),
23138 => conv_std_logic_vector(34, 8),
23139 => conv_std_logic_vector(34, 8),
23140 => conv_std_logic_vector(35, 8),
23141 => conv_std_logic_vector(35, 8),
23142 => conv_std_logic_vector(35, 8),
23143 => conv_std_logic_vector(36, 8),
23144 => conv_std_logic_vector(36, 8),
23145 => conv_std_logic_vector(36, 8),
23146 => conv_std_logic_vector(37, 8),
23147 => conv_std_logic_vector(37, 8),
23148 => conv_std_logic_vector(37, 8),
23149 => conv_std_logic_vector(38, 8),
23150 => conv_std_logic_vector(38, 8),
23151 => conv_std_logic_vector(39, 8),
23152 => conv_std_logic_vector(39, 8),
23153 => conv_std_logic_vector(39, 8),
23154 => conv_std_logic_vector(40, 8),
23155 => conv_std_logic_vector(40, 8),
23156 => conv_std_logic_vector(40, 8),
23157 => conv_std_logic_vector(41, 8),
23158 => conv_std_logic_vector(41, 8),
23159 => conv_std_logic_vector(41, 8),
23160 => conv_std_logic_vector(42, 8),
23161 => conv_std_logic_vector(42, 8),
23162 => conv_std_logic_vector(42, 8),
23163 => conv_std_logic_vector(43, 8),
23164 => conv_std_logic_vector(43, 8),
23165 => conv_std_logic_vector(43, 8),
23166 => conv_std_logic_vector(44, 8),
23167 => conv_std_logic_vector(44, 8),
23168 => conv_std_logic_vector(45, 8),
23169 => conv_std_logic_vector(45, 8),
23170 => conv_std_logic_vector(45, 8),
23171 => conv_std_logic_vector(46, 8),
23172 => conv_std_logic_vector(46, 8),
23173 => conv_std_logic_vector(46, 8),
23174 => conv_std_logic_vector(47, 8),
23175 => conv_std_logic_vector(47, 8),
23176 => conv_std_logic_vector(47, 8),
23177 => conv_std_logic_vector(48, 8),
23178 => conv_std_logic_vector(48, 8),
23179 => conv_std_logic_vector(48, 8),
23180 => conv_std_logic_vector(49, 8),
23181 => conv_std_logic_vector(49, 8),
23182 => conv_std_logic_vector(49, 8),
23183 => conv_std_logic_vector(50, 8),
23184 => conv_std_logic_vector(50, 8),
23185 => conv_std_logic_vector(50, 8),
23186 => conv_std_logic_vector(51, 8),
23187 => conv_std_logic_vector(51, 8),
23188 => conv_std_logic_vector(52, 8),
23189 => conv_std_logic_vector(52, 8),
23190 => conv_std_logic_vector(52, 8),
23191 => conv_std_logic_vector(53, 8),
23192 => conv_std_logic_vector(53, 8),
23193 => conv_std_logic_vector(53, 8),
23194 => conv_std_logic_vector(54, 8),
23195 => conv_std_logic_vector(54, 8),
23196 => conv_std_logic_vector(54, 8),
23197 => conv_std_logic_vector(55, 8),
23198 => conv_std_logic_vector(55, 8),
23199 => conv_std_logic_vector(55, 8),
23200 => conv_std_logic_vector(56, 8),
23201 => conv_std_logic_vector(56, 8),
23202 => conv_std_logic_vector(56, 8),
23203 => conv_std_logic_vector(57, 8),
23204 => conv_std_logic_vector(57, 8),
23205 => conv_std_logic_vector(58, 8),
23206 => conv_std_logic_vector(58, 8),
23207 => conv_std_logic_vector(58, 8),
23208 => conv_std_logic_vector(59, 8),
23209 => conv_std_logic_vector(59, 8),
23210 => conv_std_logic_vector(59, 8),
23211 => conv_std_logic_vector(60, 8),
23212 => conv_std_logic_vector(60, 8),
23213 => conv_std_logic_vector(60, 8),
23214 => conv_std_logic_vector(61, 8),
23215 => conv_std_logic_vector(61, 8),
23216 => conv_std_logic_vector(61, 8),
23217 => conv_std_logic_vector(62, 8),
23218 => conv_std_logic_vector(62, 8),
23219 => conv_std_logic_vector(62, 8),
23220 => conv_std_logic_vector(63, 8),
23221 => conv_std_logic_vector(63, 8),
23222 => conv_std_logic_vector(63, 8),
23223 => conv_std_logic_vector(64, 8),
23224 => conv_std_logic_vector(64, 8),
23225 => conv_std_logic_vector(65, 8),
23226 => conv_std_logic_vector(65, 8),
23227 => conv_std_logic_vector(65, 8),
23228 => conv_std_logic_vector(66, 8),
23229 => conv_std_logic_vector(66, 8),
23230 => conv_std_logic_vector(66, 8),
23231 => conv_std_logic_vector(67, 8),
23232 => conv_std_logic_vector(67, 8),
23233 => conv_std_logic_vector(67, 8),
23234 => conv_std_logic_vector(68, 8),
23235 => conv_std_logic_vector(68, 8),
23236 => conv_std_logic_vector(68, 8),
23237 => conv_std_logic_vector(69, 8),
23238 => conv_std_logic_vector(69, 8),
23239 => conv_std_logic_vector(69, 8),
23240 => conv_std_logic_vector(70, 8),
23241 => conv_std_logic_vector(70, 8),
23242 => conv_std_logic_vector(71, 8),
23243 => conv_std_logic_vector(71, 8),
23244 => conv_std_logic_vector(71, 8),
23245 => conv_std_logic_vector(72, 8),
23246 => conv_std_logic_vector(72, 8),
23247 => conv_std_logic_vector(72, 8),
23248 => conv_std_logic_vector(73, 8),
23249 => conv_std_logic_vector(73, 8),
23250 => conv_std_logic_vector(73, 8),
23251 => conv_std_logic_vector(74, 8),
23252 => conv_std_logic_vector(74, 8),
23253 => conv_std_logic_vector(74, 8),
23254 => conv_std_logic_vector(75, 8),
23255 => conv_std_logic_vector(75, 8),
23256 => conv_std_logic_vector(75, 8),
23257 => conv_std_logic_vector(76, 8),
23258 => conv_std_logic_vector(76, 8),
23259 => conv_std_logic_vector(76, 8),
23260 => conv_std_logic_vector(77, 8),
23261 => conv_std_logic_vector(77, 8),
23262 => conv_std_logic_vector(78, 8),
23263 => conv_std_logic_vector(78, 8),
23264 => conv_std_logic_vector(78, 8),
23265 => conv_std_logic_vector(79, 8),
23266 => conv_std_logic_vector(79, 8),
23267 => conv_std_logic_vector(79, 8),
23268 => conv_std_logic_vector(80, 8),
23269 => conv_std_logic_vector(80, 8),
23270 => conv_std_logic_vector(80, 8),
23271 => conv_std_logic_vector(81, 8),
23272 => conv_std_logic_vector(81, 8),
23273 => conv_std_logic_vector(81, 8),
23274 => conv_std_logic_vector(82, 8),
23275 => conv_std_logic_vector(82, 8),
23276 => conv_std_logic_vector(82, 8),
23277 => conv_std_logic_vector(83, 8),
23278 => conv_std_logic_vector(83, 8),
23279 => conv_std_logic_vector(84, 8),
23280 => conv_std_logic_vector(84, 8),
23281 => conv_std_logic_vector(84, 8),
23282 => conv_std_logic_vector(85, 8),
23283 => conv_std_logic_vector(85, 8),
23284 => conv_std_logic_vector(85, 8),
23285 => conv_std_logic_vector(86, 8),
23286 => conv_std_logic_vector(86, 8),
23287 => conv_std_logic_vector(86, 8),
23288 => conv_std_logic_vector(87, 8),
23289 => conv_std_logic_vector(87, 8),
23290 => conv_std_logic_vector(87, 8),
23291 => conv_std_logic_vector(88, 8),
23292 => conv_std_logic_vector(88, 8),
23293 => conv_std_logic_vector(88, 8),
23294 => conv_std_logic_vector(89, 8),
23295 => conv_std_logic_vector(89, 8),
23296 => conv_std_logic_vector(0, 8),
23297 => conv_std_logic_vector(0, 8),
23298 => conv_std_logic_vector(0, 8),
23299 => conv_std_logic_vector(1, 8),
23300 => conv_std_logic_vector(1, 8),
23301 => conv_std_logic_vector(1, 8),
23302 => conv_std_logic_vector(2, 8),
23303 => conv_std_logic_vector(2, 8),
23304 => conv_std_logic_vector(2, 8),
23305 => conv_std_logic_vector(3, 8),
23306 => conv_std_logic_vector(3, 8),
23307 => conv_std_logic_vector(3, 8),
23308 => conv_std_logic_vector(4, 8),
23309 => conv_std_logic_vector(4, 8),
23310 => conv_std_logic_vector(4, 8),
23311 => conv_std_logic_vector(5, 8),
23312 => conv_std_logic_vector(5, 8),
23313 => conv_std_logic_vector(6, 8),
23314 => conv_std_logic_vector(6, 8),
23315 => conv_std_logic_vector(6, 8),
23316 => conv_std_logic_vector(7, 8),
23317 => conv_std_logic_vector(7, 8),
23318 => conv_std_logic_vector(7, 8),
23319 => conv_std_logic_vector(8, 8),
23320 => conv_std_logic_vector(8, 8),
23321 => conv_std_logic_vector(8, 8),
23322 => conv_std_logic_vector(9, 8),
23323 => conv_std_logic_vector(9, 8),
23324 => conv_std_logic_vector(9, 8),
23325 => conv_std_logic_vector(10, 8),
23326 => conv_std_logic_vector(10, 8),
23327 => conv_std_logic_vector(11, 8),
23328 => conv_std_logic_vector(11, 8),
23329 => conv_std_logic_vector(11, 8),
23330 => conv_std_logic_vector(12, 8),
23331 => conv_std_logic_vector(12, 8),
23332 => conv_std_logic_vector(12, 8),
23333 => conv_std_logic_vector(13, 8),
23334 => conv_std_logic_vector(13, 8),
23335 => conv_std_logic_vector(13, 8),
23336 => conv_std_logic_vector(14, 8),
23337 => conv_std_logic_vector(14, 8),
23338 => conv_std_logic_vector(14, 8),
23339 => conv_std_logic_vector(15, 8),
23340 => conv_std_logic_vector(15, 8),
23341 => conv_std_logic_vector(15, 8),
23342 => conv_std_logic_vector(16, 8),
23343 => conv_std_logic_vector(16, 8),
23344 => conv_std_logic_vector(17, 8),
23345 => conv_std_logic_vector(17, 8),
23346 => conv_std_logic_vector(17, 8),
23347 => conv_std_logic_vector(18, 8),
23348 => conv_std_logic_vector(18, 8),
23349 => conv_std_logic_vector(18, 8),
23350 => conv_std_logic_vector(19, 8),
23351 => conv_std_logic_vector(19, 8),
23352 => conv_std_logic_vector(19, 8),
23353 => conv_std_logic_vector(20, 8),
23354 => conv_std_logic_vector(20, 8),
23355 => conv_std_logic_vector(20, 8),
23356 => conv_std_logic_vector(21, 8),
23357 => conv_std_logic_vector(21, 8),
23358 => conv_std_logic_vector(22, 8),
23359 => conv_std_logic_vector(22, 8),
23360 => conv_std_logic_vector(22, 8),
23361 => conv_std_logic_vector(23, 8),
23362 => conv_std_logic_vector(23, 8),
23363 => conv_std_logic_vector(23, 8),
23364 => conv_std_logic_vector(24, 8),
23365 => conv_std_logic_vector(24, 8),
23366 => conv_std_logic_vector(24, 8),
23367 => conv_std_logic_vector(25, 8),
23368 => conv_std_logic_vector(25, 8),
23369 => conv_std_logic_vector(25, 8),
23370 => conv_std_logic_vector(26, 8),
23371 => conv_std_logic_vector(26, 8),
23372 => conv_std_logic_vector(27, 8),
23373 => conv_std_logic_vector(27, 8),
23374 => conv_std_logic_vector(27, 8),
23375 => conv_std_logic_vector(28, 8),
23376 => conv_std_logic_vector(28, 8),
23377 => conv_std_logic_vector(28, 8),
23378 => conv_std_logic_vector(29, 8),
23379 => conv_std_logic_vector(29, 8),
23380 => conv_std_logic_vector(29, 8),
23381 => conv_std_logic_vector(30, 8),
23382 => conv_std_logic_vector(30, 8),
23383 => conv_std_logic_vector(30, 8),
23384 => conv_std_logic_vector(31, 8),
23385 => conv_std_logic_vector(31, 8),
23386 => conv_std_logic_vector(31, 8),
23387 => conv_std_logic_vector(32, 8),
23388 => conv_std_logic_vector(32, 8),
23389 => conv_std_logic_vector(33, 8),
23390 => conv_std_logic_vector(33, 8),
23391 => conv_std_logic_vector(33, 8),
23392 => conv_std_logic_vector(34, 8),
23393 => conv_std_logic_vector(34, 8),
23394 => conv_std_logic_vector(34, 8),
23395 => conv_std_logic_vector(35, 8),
23396 => conv_std_logic_vector(35, 8),
23397 => conv_std_logic_vector(35, 8),
23398 => conv_std_logic_vector(36, 8),
23399 => conv_std_logic_vector(36, 8),
23400 => conv_std_logic_vector(36, 8),
23401 => conv_std_logic_vector(37, 8),
23402 => conv_std_logic_vector(37, 8),
23403 => conv_std_logic_vector(38, 8),
23404 => conv_std_logic_vector(38, 8),
23405 => conv_std_logic_vector(38, 8),
23406 => conv_std_logic_vector(39, 8),
23407 => conv_std_logic_vector(39, 8),
23408 => conv_std_logic_vector(39, 8),
23409 => conv_std_logic_vector(40, 8),
23410 => conv_std_logic_vector(40, 8),
23411 => conv_std_logic_vector(40, 8),
23412 => conv_std_logic_vector(41, 8),
23413 => conv_std_logic_vector(41, 8),
23414 => conv_std_logic_vector(41, 8),
23415 => conv_std_logic_vector(42, 8),
23416 => conv_std_logic_vector(42, 8),
23417 => conv_std_logic_vector(43, 8),
23418 => conv_std_logic_vector(43, 8),
23419 => conv_std_logic_vector(43, 8),
23420 => conv_std_logic_vector(44, 8),
23421 => conv_std_logic_vector(44, 8),
23422 => conv_std_logic_vector(44, 8),
23423 => conv_std_logic_vector(45, 8),
23424 => conv_std_logic_vector(45, 8),
23425 => conv_std_logic_vector(45, 8),
23426 => conv_std_logic_vector(46, 8),
23427 => conv_std_logic_vector(46, 8),
23428 => conv_std_logic_vector(46, 8),
23429 => conv_std_logic_vector(47, 8),
23430 => conv_std_logic_vector(47, 8),
23431 => conv_std_logic_vector(47, 8),
23432 => conv_std_logic_vector(48, 8),
23433 => conv_std_logic_vector(48, 8),
23434 => conv_std_logic_vector(49, 8),
23435 => conv_std_logic_vector(49, 8),
23436 => conv_std_logic_vector(49, 8),
23437 => conv_std_logic_vector(50, 8),
23438 => conv_std_logic_vector(50, 8),
23439 => conv_std_logic_vector(50, 8),
23440 => conv_std_logic_vector(51, 8),
23441 => conv_std_logic_vector(51, 8),
23442 => conv_std_logic_vector(51, 8),
23443 => conv_std_logic_vector(52, 8),
23444 => conv_std_logic_vector(52, 8),
23445 => conv_std_logic_vector(52, 8),
23446 => conv_std_logic_vector(53, 8),
23447 => conv_std_logic_vector(53, 8),
23448 => conv_std_logic_vector(54, 8),
23449 => conv_std_logic_vector(54, 8),
23450 => conv_std_logic_vector(54, 8),
23451 => conv_std_logic_vector(55, 8),
23452 => conv_std_logic_vector(55, 8),
23453 => conv_std_logic_vector(55, 8),
23454 => conv_std_logic_vector(56, 8),
23455 => conv_std_logic_vector(56, 8),
23456 => conv_std_logic_vector(56, 8),
23457 => conv_std_logic_vector(57, 8),
23458 => conv_std_logic_vector(57, 8),
23459 => conv_std_logic_vector(57, 8),
23460 => conv_std_logic_vector(58, 8),
23461 => conv_std_logic_vector(58, 8),
23462 => conv_std_logic_vector(59, 8),
23463 => conv_std_logic_vector(59, 8),
23464 => conv_std_logic_vector(59, 8),
23465 => conv_std_logic_vector(60, 8),
23466 => conv_std_logic_vector(60, 8),
23467 => conv_std_logic_vector(60, 8),
23468 => conv_std_logic_vector(61, 8),
23469 => conv_std_logic_vector(61, 8),
23470 => conv_std_logic_vector(61, 8),
23471 => conv_std_logic_vector(62, 8),
23472 => conv_std_logic_vector(62, 8),
23473 => conv_std_logic_vector(62, 8),
23474 => conv_std_logic_vector(63, 8),
23475 => conv_std_logic_vector(63, 8),
23476 => conv_std_logic_vector(63, 8),
23477 => conv_std_logic_vector(64, 8),
23478 => conv_std_logic_vector(64, 8),
23479 => conv_std_logic_vector(65, 8),
23480 => conv_std_logic_vector(65, 8),
23481 => conv_std_logic_vector(65, 8),
23482 => conv_std_logic_vector(66, 8),
23483 => conv_std_logic_vector(66, 8),
23484 => conv_std_logic_vector(66, 8),
23485 => conv_std_logic_vector(67, 8),
23486 => conv_std_logic_vector(67, 8),
23487 => conv_std_logic_vector(67, 8),
23488 => conv_std_logic_vector(68, 8),
23489 => conv_std_logic_vector(68, 8),
23490 => conv_std_logic_vector(68, 8),
23491 => conv_std_logic_vector(69, 8),
23492 => conv_std_logic_vector(69, 8),
23493 => conv_std_logic_vector(70, 8),
23494 => conv_std_logic_vector(70, 8),
23495 => conv_std_logic_vector(70, 8),
23496 => conv_std_logic_vector(71, 8),
23497 => conv_std_logic_vector(71, 8),
23498 => conv_std_logic_vector(71, 8),
23499 => conv_std_logic_vector(72, 8),
23500 => conv_std_logic_vector(72, 8),
23501 => conv_std_logic_vector(72, 8),
23502 => conv_std_logic_vector(73, 8),
23503 => conv_std_logic_vector(73, 8),
23504 => conv_std_logic_vector(73, 8),
23505 => conv_std_logic_vector(74, 8),
23506 => conv_std_logic_vector(74, 8),
23507 => conv_std_logic_vector(75, 8),
23508 => conv_std_logic_vector(75, 8),
23509 => conv_std_logic_vector(75, 8),
23510 => conv_std_logic_vector(76, 8),
23511 => conv_std_logic_vector(76, 8),
23512 => conv_std_logic_vector(76, 8),
23513 => conv_std_logic_vector(77, 8),
23514 => conv_std_logic_vector(77, 8),
23515 => conv_std_logic_vector(77, 8),
23516 => conv_std_logic_vector(78, 8),
23517 => conv_std_logic_vector(78, 8),
23518 => conv_std_logic_vector(78, 8),
23519 => conv_std_logic_vector(79, 8),
23520 => conv_std_logic_vector(79, 8),
23521 => conv_std_logic_vector(79, 8),
23522 => conv_std_logic_vector(80, 8),
23523 => conv_std_logic_vector(80, 8),
23524 => conv_std_logic_vector(81, 8),
23525 => conv_std_logic_vector(81, 8),
23526 => conv_std_logic_vector(81, 8),
23527 => conv_std_logic_vector(82, 8),
23528 => conv_std_logic_vector(82, 8),
23529 => conv_std_logic_vector(82, 8),
23530 => conv_std_logic_vector(83, 8),
23531 => conv_std_logic_vector(83, 8),
23532 => conv_std_logic_vector(83, 8),
23533 => conv_std_logic_vector(84, 8),
23534 => conv_std_logic_vector(84, 8),
23535 => conv_std_logic_vector(84, 8),
23536 => conv_std_logic_vector(85, 8),
23537 => conv_std_logic_vector(85, 8),
23538 => conv_std_logic_vector(86, 8),
23539 => conv_std_logic_vector(86, 8),
23540 => conv_std_logic_vector(86, 8),
23541 => conv_std_logic_vector(87, 8),
23542 => conv_std_logic_vector(87, 8),
23543 => conv_std_logic_vector(87, 8),
23544 => conv_std_logic_vector(88, 8),
23545 => conv_std_logic_vector(88, 8),
23546 => conv_std_logic_vector(88, 8),
23547 => conv_std_logic_vector(89, 8),
23548 => conv_std_logic_vector(89, 8),
23549 => conv_std_logic_vector(89, 8),
23550 => conv_std_logic_vector(90, 8),
23551 => conv_std_logic_vector(90, 8),
23552 => conv_std_logic_vector(0, 8),
23553 => conv_std_logic_vector(0, 8),
23554 => conv_std_logic_vector(0, 8),
23555 => conv_std_logic_vector(1, 8),
23556 => conv_std_logic_vector(1, 8),
23557 => conv_std_logic_vector(1, 8),
23558 => conv_std_logic_vector(2, 8),
23559 => conv_std_logic_vector(2, 8),
23560 => conv_std_logic_vector(2, 8),
23561 => conv_std_logic_vector(3, 8),
23562 => conv_std_logic_vector(3, 8),
23563 => conv_std_logic_vector(3, 8),
23564 => conv_std_logic_vector(4, 8),
23565 => conv_std_logic_vector(4, 8),
23566 => conv_std_logic_vector(5, 8),
23567 => conv_std_logic_vector(5, 8),
23568 => conv_std_logic_vector(5, 8),
23569 => conv_std_logic_vector(6, 8),
23570 => conv_std_logic_vector(6, 8),
23571 => conv_std_logic_vector(6, 8),
23572 => conv_std_logic_vector(7, 8),
23573 => conv_std_logic_vector(7, 8),
23574 => conv_std_logic_vector(7, 8),
23575 => conv_std_logic_vector(8, 8),
23576 => conv_std_logic_vector(8, 8),
23577 => conv_std_logic_vector(8, 8),
23578 => conv_std_logic_vector(9, 8),
23579 => conv_std_logic_vector(9, 8),
23580 => conv_std_logic_vector(10, 8),
23581 => conv_std_logic_vector(10, 8),
23582 => conv_std_logic_vector(10, 8),
23583 => conv_std_logic_vector(11, 8),
23584 => conv_std_logic_vector(11, 8),
23585 => conv_std_logic_vector(11, 8),
23586 => conv_std_logic_vector(12, 8),
23587 => conv_std_logic_vector(12, 8),
23588 => conv_std_logic_vector(12, 8),
23589 => conv_std_logic_vector(13, 8),
23590 => conv_std_logic_vector(13, 8),
23591 => conv_std_logic_vector(14, 8),
23592 => conv_std_logic_vector(14, 8),
23593 => conv_std_logic_vector(14, 8),
23594 => conv_std_logic_vector(15, 8),
23595 => conv_std_logic_vector(15, 8),
23596 => conv_std_logic_vector(15, 8),
23597 => conv_std_logic_vector(16, 8),
23598 => conv_std_logic_vector(16, 8),
23599 => conv_std_logic_vector(16, 8),
23600 => conv_std_logic_vector(17, 8),
23601 => conv_std_logic_vector(17, 8),
23602 => conv_std_logic_vector(17, 8),
23603 => conv_std_logic_vector(18, 8),
23604 => conv_std_logic_vector(18, 8),
23605 => conv_std_logic_vector(19, 8),
23606 => conv_std_logic_vector(19, 8),
23607 => conv_std_logic_vector(19, 8),
23608 => conv_std_logic_vector(20, 8),
23609 => conv_std_logic_vector(20, 8),
23610 => conv_std_logic_vector(20, 8),
23611 => conv_std_logic_vector(21, 8),
23612 => conv_std_logic_vector(21, 8),
23613 => conv_std_logic_vector(21, 8),
23614 => conv_std_logic_vector(22, 8),
23615 => conv_std_logic_vector(22, 8),
23616 => conv_std_logic_vector(23, 8),
23617 => conv_std_logic_vector(23, 8),
23618 => conv_std_logic_vector(23, 8),
23619 => conv_std_logic_vector(24, 8),
23620 => conv_std_logic_vector(24, 8),
23621 => conv_std_logic_vector(24, 8),
23622 => conv_std_logic_vector(25, 8),
23623 => conv_std_logic_vector(25, 8),
23624 => conv_std_logic_vector(25, 8),
23625 => conv_std_logic_vector(26, 8),
23626 => conv_std_logic_vector(26, 8),
23627 => conv_std_logic_vector(26, 8),
23628 => conv_std_logic_vector(27, 8),
23629 => conv_std_logic_vector(27, 8),
23630 => conv_std_logic_vector(28, 8),
23631 => conv_std_logic_vector(28, 8),
23632 => conv_std_logic_vector(28, 8),
23633 => conv_std_logic_vector(29, 8),
23634 => conv_std_logic_vector(29, 8),
23635 => conv_std_logic_vector(29, 8),
23636 => conv_std_logic_vector(30, 8),
23637 => conv_std_logic_vector(30, 8),
23638 => conv_std_logic_vector(30, 8),
23639 => conv_std_logic_vector(31, 8),
23640 => conv_std_logic_vector(31, 8),
23641 => conv_std_logic_vector(31, 8),
23642 => conv_std_logic_vector(32, 8),
23643 => conv_std_logic_vector(32, 8),
23644 => conv_std_logic_vector(33, 8),
23645 => conv_std_logic_vector(33, 8),
23646 => conv_std_logic_vector(33, 8),
23647 => conv_std_logic_vector(34, 8),
23648 => conv_std_logic_vector(34, 8),
23649 => conv_std_logic_vector(34, 8),
23650 => conv_std_logic_vector(35, 8),
23651 => conv_std_logic_vector(35, 8),
23652 => conv_std_logic_vector(35, 8),
23653 => conv_std_logic_vector(36, 8),
23654 => conv_std_logic_vector(36, 8),
23655 => conv_std_logic_vector(37, 8),
23656 => conv_std_logic_vector(37, 8),
23657 => conv_std_logic_vector(37, 8),
23658 => conv_std_logic_vector(38, 8),
23659 => conv_std_logic_vector(38, 8),
23660 => conv_std_logic_vector(38, 8),
23661 => conv_std_logic_vector(39, 8),
23662 => conv_std_logic_vector(39, 8),
23663 => conv_std_logic_vector(39, 8),
23664 => conv_std_logic_vector(40, 8),
23665 => conv_std_logic_vector(40, 8),
23666 => conv_std_logic_vector(40, 8),
23667 => conv_std_logic_vector(41, 8),
23668 => conv_std_logic_vector(41, 8),
23669 => conv_std_logic_vector(42, 8),
23670 => conv_std_logic_vector(42, 8),
23671 => conv_std_logic_vector(42, 8),
23672 => conv_std_logic_vector(43, 8),
23673 => conv_std_logic_vector(43, 8),
23674 => conv_std_logic_vector(43, 8),
23675 => conv_std_logic_vector(44, 8),
23676 => conv_std_logic_vector(44, 8),
23677 => conv_std_logic_vector(44, 8),
23678 => conv_std_logic_vector(45, 8),
23679 => conv_std_logic_vector(45, 8),
23680 => conv_std_logic_vector(46, 8),
23681 => conv_std_logic_vector(46, 8),
23682 => conv_std_logic_vector(46, 8),
23683 => conv_std_logic_vector(47, 8),
23684 => conv_std_logic_vector(47, 8),
23685 => conv_std_logic_vector(47, 8),
23686 => conv_std_logic_vector(48, 8),
23687 => conv_std_logic_vector(48, 8),
23688 => conv_std_logic_vector(48, 8),
23689 => conv_std_logic_vector(49, 8),
23690 => conv_std_logic_vector(49, 8),
23691 => conv_std_logic_vector(49, 8),
23692 => conv_std_logic_vector(50, 8),
23693 => conv_std_logic_vector(50, 8),
23694 => conv_std_logic_vector(51, 8),
23695 => conv_std_logic_vector(51, 8),
23696 => conv_std_logic_vector(51, 8),
23697 => conv_std_logic_vector(52, 8),
23698 => conv_std_logic_vector(52, 8),
23699 => conv_std_logic_vector(52, 8),
23700 => conv_std_logic_vector(53, 8),
23701 => conv_std_logic_vector(53, 8),
23702 => conv_std_logic_vector(53, 8),
23703 => conv_std_logic_vector(54, 8),
23704 => conv_std_logic_vector(54, 8),
23705 => conv_std_logic_vector(54, 8),
23706 => conv_std_logic_vector(55, 8),
23707 => conv_std_logic_vector(55, 8),
23708 => conv_std_logic_vector(56, 8),
23709 => conv_std_logic_vector(56, 8),
23710 => conv_std_logic_vector(56, 8),
23711 => conv_std_logic_vector(57, 8),
23712 => conv_std_logic_vector(57, 8),
23713 => conv_std_logic_vector(57, 8),
23714 => conv_std_logic_vector(58, 8),
23715 => conv_std_logic_vector(58, 8),
23716 => conv_std_logic_vector(58, 8),
23717 => conv_std_logic_vector(59, 8),
23718 => conv_std_logic_vector(59, 8),
23719 => conv_std_logic_vector(60, 8),
23720 => conv_std_logic_vector(60, 8),
23721 => conv_std_logic_vector(60, 8),
23722 => conv_std_logic_vector(61, 8),
23723 => conv_std_logic_vector(61, 8),
23724 => conv_std_logic_vector(61, 8),
23725 => conv_std_logic_vector(62, 8),
23726 => conv_std_logic_vector(62, 8),
23727 => conv_std_logic_vector(62, 8),
23728 => conv_std_logic_vector(63, 8),
23729 => conv_std_logic_vector(63, 8),
23730 => conv_std_logic_vector(63, 8),
23731 => conv_std_logic_vector(64, 8),
23732 => conv_std_logic_vector(64, 8),
23733 => conv_std_logic_vector(65, 8),
23734 => conv_std_logic_vector(65, 8),
23735 => conv_std_logic_vector(65, 8),
23736 => conv_std_logic_vector(66, 8),
23737 => conv_std_logic_vector(66, 8),
23738 => conv_std_logic_vector(66, 8),
23739 => conv_std_logic_vector(67, 8),
23740 => conv_std_logic_vector(67, 8),
23741 => conv_std_logic_vector(67, 8),
23742 => conv_std_logic_vector(68, 8),
23743 => conv_std_logic_vector(68, 8),
23744 => conv_std_logic_vector(69, 8),
23745 => conv_std_logic_vector(69, 8),
23746 => conv_std_logic_vector(69, 8),
23747 => conv_std_logic_vector(70, 8),
23748 => conv_std_logic_vector(70, 8),
23749 => conv_std_logic_vector(70, 8),
23750 => conv_std_logic_vector(71, 8),
23751 => conv_std_logic_vector(71, 8),
23752 => conv_std_logic_vector(71, 8),
23753 => conv_std_logic_vector(72, 8),
23754 => conv_std_logic_vector(72, 8),
23755 => conv_std_logic_vector(72, 8),
23756 => conv_std_logic_vector(73, 8),
23757 => conv_std_logic_vector(73, 8),
23758 => conv_std_logic_vector(74, 8),
23759 => conv_std_logic_vector(74, 8),
23760 => conv_std_logic_vector(74, 8),
23761 => conv_std_logic_vector(75, 8),
23762 => conv_std_logic_vector(75, 8),
23763 => conv_std_logic_vector(75, 8),
23764 => conv_std_logic_vector(76, 8),
23765 => conv_std_logic_vector(76, 8),
23766 => conv_std_logic_vector(76, 8),
23767 => conv_std_logic_vector(77, 8),
23768 => conv_std_logic_vector(77, 8),
23769 => conv_std_logic_vector(77, 8),
23770 => conv_std_logic_vector(78, 8),
23771 => conv_std_logic_vector(78, 8),
23772 => conv_std_logic_vector(79, 8),
23773 => conv_std_logic_vector(79, 8),
23774 => conv_std_logic_vector(79, 8),
23775 => conv_std_logic_vector(80, 8),
23776 => conv_std_logic_vector(80, 8),
23777 => conv_std_logic_vector(80, 8),
23778 => conv_std_logic_vector(81, 8),
23779 => conv_std_logic_vector(81, 8),
23780 => conv_std_logic_vector(81, 8),
23781 => conv_std_logic_vector(82, 8),
23782 => conv_std_logic_vector(82, 8),
23783 => conv_std_logic_vector(83, 8),
23784 => conv_std_logic_vector(83, 8),
23785 => conv_std_logic_vector(83, 8),
23786 => conv_std_logic_vector(84, 8),
23787 => conv_std_logic_vector(84, 8),
23788 => conv_std_logic_vector(84, 8),
23789 => conv_std_logic_vector(85, 8),
23790 => conv_std_logic_vector(85, 8),
23791 => conv_std_logic_vector(85, 8),
23792 => conv_std_logic_vector(86, 8),
23793 => conv_std_logic_vector(86, 8),
23794 => conv_std_logic_vector(86, 8),
23795 => conv_std_logic_vector(87, 8),
23796 => conv_std_logic_vector(87, 8),
23797 => conv_std_logic_vector(88, 8),
23798 => conv_std_logic_vector(88, 8),
23799 => conv_std_logic_vector(88, 8),
23800 => conv_std_logic_vector(89, 8),
23801 => conv_std_logic_vector(89, 8),
23802 => conv_std_logic_vector(89, 8),
23803 => conv_std_logic_vector(90, 8),
23804 => conv_std_logic_vector(90, 8),
23805 => conv_std_logic_vector(90, 8),
23806 => conv_std_logic_vector(91, 8),
23807 => conv_std_logic_vector(91, 8),
23808 => conv_std_logic_vector(0, 8),
23809 => conv_std_logic_vector(0, 8),
23810 => conv_std_logic_vector(0, 8),
23811 => conv_std_logic_vector(1, 8),
23812 => conv_std_logic_vector(1, 8),
23813 => conv_std_logic_vector(1, 8),
23814 => conv_std_logic_vector(2, 8),
23815 => conv_std_logic_vector(2, 8),
23816 => conv_std_logic_vector(2, 8),
23817 => conv_std_logic_vector(3, 8),
23818 => conv_std_logic_vector(3, 8),
23819 => conv_std_logic_vector(3, 8),
23820 => conv_std_logic_vector(4, 8),
23821 => conv_std_logic_vector(4, 8),
23822 => conv_std_logic_vector(5, 8),
23823 => conv_std_logic_vector(5, 8),
23824 => conv_std_logic_vector(5, 8),
23825 => conv_std_logic_vector(6, 8),
23826 => conv_std_logic_vector(6, 8),
23827 => conv_std_logic_vector(6, 8),
23828 => conv_std_logic_vector(7, 8),
23829 => conv_std_logic_vector(7, 8),
23830 => conv_std_logic_vector(7, 8),
23831 => conv_std_logic_vector(8, 8),
23832 => conv_std_logic_vector(8, 8),
23833 => conv_std_logic_vector(9, 8),
23834 => conv_std_logic_vector(9, 8),
23835 => conv_std_logic_vector(9, 8),
23836 => conv_std_logic_vector(10, 8),
23837 => conv_std_logic_vector(10, 8),
23838 => conv_std_logic_vector(10, 8),
23839 => conv_std_logic_vector(11, 8),
23840 => conv_std_logic_vector(11, 8),
23841 => conv_std_logic_vector(11, 8),
23842 => conv_std_logic_vector(12, 8),
23843 => conv_std_logic_vector(12, 8),
23844 => conv_std_logic_vector(13, 8),
23845 => conv_std_logic_vector(13, 8),
23846 => conv_std_logic_vector(13, 8),
23847 => conv_std_logic_vector(14, 8),
23848 => conv_std_logic_vector(14, 8),
23849 => conv_std_logic_vector(14, 8),
23850 => conv_std_logic_vector(15, 8),
23851 => conv_std_logic_vector(15, 8),
23852 => conv_std_logic_vector(15, 8),
23853 => conv_std_logic_vector(16, 8),
23854 => conv_std_logic_vector(16, 8),
23855 => conv_std_logic_vector(17, 8),
23856 => conv_std_logic_vector(17, 8),
23857 => conv_std_logic_vector(17, 8),
23858 => conv_std_logic_vector(18, 8),
23859 => conv_std_logic_vector(18, 8),
23860 => conv_std_logic_vector(18, 8),
23861 => conv_std_logic_vector(19, 8),
23862 => conv_std_logic_vector(19, 8),
23863 => conv_std_logic_vector(19, 8),
23864 => conv_std_logic_vector(20, 8),
23865 => conv_std_logic_vector(20, 8),
23866 => conv_std_logic_vector(21, 8),
23867 => conv_std_logic_vector(21, 8),
23868 => conv_std_logic_vector(21, 8),
23869 => conv_std_logic_vector(22, 8),
23870 => conv_std_logic_vector(22, 8),
23871 => conv_std_logic_vector(22, 8),
23872 => conv_std_logic_vector(23, 8),
23873 => conv_std_logic_vector(23, 8),
23874 => conv_std_logic_vector(23, 8),
23875 => conv_std_logic_vector(24, 8),
23876 => conv_std_logic_vector(24, 8),
23877 => conv_std_logic_vector(25, 8),
23878 => conv_std_logic_vector(25, 8),
23879 => conv_std_logic_vector(25, 8),
23880 => conv_std_logic_vector(26, 8),
23881 => conv_std_logic_vector(26, 8),
23882 => conv_std_logic_vector(26, 8),
23883 => conv_std_logic_vector(27, 8),
23884 => conv_std_logic_vector(27, 8),
23885 => conv_std_logic_vector(27, 8),
23886 => conv_std_logic_vector(28, 8),
23887 => conv_std_logic_vector(28, 8),
23888 => conv_std_logic_vector(29, 8),
23889 => conv_std_logic_vector(29, 8),
23890 => conv_std_logic_vector(29, 8),
23891 => conv_std_logic_vector(30, 8),
23892 => conv_std_logic_vector(30, 8),
23893 => conv_std_logic_vector(30, 8),
23894 => conv_std_logic_vector(31, 8),
23895 => conv_std_logic_vector(31, 8),
23896 => conv_std_logic_vector(31, 8),
23897 => conv_std_logic_vector(32, 8),
23898 => conv_std_logic_vector(32, 8),
23899 => conv_std_logic_vector(33, 8),
23900 => conv_std_logic_vector(33, 8),
23901 => conv_std_logic_vector(33, 8),
23902 => conv_std_logic_vector(34, 8),
23903 => conv_std_logic_vector(34, 8),
23904 => conv_std_logic_vector(34, 8),
23905 => conv_std_logic_vector(35, 8),
23906 => conv_std_logic_vector(35, 8),
23907 => conv_std_logic_vector(35, 8),
23908 => conv_std_logic_vector(36, 8),
23909 => conv_std_logic_vector(36, 8),
23910 => conv_std_logic_vector(37, 8),
23911 => conv_std_logic_vector(37, 8),
23912 => conv_std_logic_vector(37, 8),
23913 => conv_std_logic_vector(38, 8),
23914 => conv_std_logic_vector(38, 8),
23915 => conv_std_logic_vector(38, 8),
23916 => conv_std_logic_vector(39, 8),
23917 => conv_std_logic_vector(39, 8),
23918 => conv_std_logic_vector(39, 8),
23919 => conv_std_logic_vector(40, 8),
23920 => conv_std_logic_vector(40, 8),
23921 => conv_std_logic_vector(41, 8),
23922 => conv_std_logic_vector(41, 8),
23923 => conv_std_logic_vector(41, 8),
23924 => conv_std_logic_vector(42, 8),
23925 => conv_std_logic_vector(42, 8),
23926 => conv_std_logic_vector(42, 8),
23927 => conv_std_logic_vector(43, 8),
23928 => conv_std_logic_vector(43, 8),
23929 => conv_std_logic_vector(43, 8),
23930 => conv_std_logic_vector(44, 8),
23931 => conv_std_logic_vector(44, 8),
23932 => conv_std_logic_vector(45, 8),
23933 => conv_std_logic_vector(45, 8),
23934 => conv_std_logic_vector(45, 8),
23935 => conv_std_logic_vector(46, 8),
23936 => conv_std_logic_vector(46, 8),
23937 => conv_std_logic_vector(46, 8),
23938 => conv_std_logic_vector(47, 8),
23939 => conv_std_logic_vector(47, 8),
23940 => conv_std_logic_vector(47, 8),
23941 => conv_std_logic_vector(48, 8),
23942 => conv_std_logic_vector(48, 8),
23943 => conv_std_logic_vector(49, 8),
23944 => conv_std_logic_vector(49, 8),
23945 => conv_std_logic_vector(49, 8),
23946 => conv_std_logic_vector(50, 8),
23947 => conv_std_logic_vector(50, 8),
23948 => conv_std_logic_vector(50, 8),
23949 => conv_std_logic_vector(51, 8),
23950 => conv_std_logic_vector(51, 8),
23951 => conv_std_logic_vector(51, 8),
23952 => conv_std_logic_vector(52, 8),
23953 => conv_std_logic_vector(52, 8),
23954 => conv_std_logic_vector(53, 8),
23955 => conv_std_logic_vector(53, 8),
23956 => conv_std_logic_vector(53, 8),
23957 => conv_std_logic_vector(54, 8),
23958 => conv_std_logic_vector(54, 8),
23959 => conv_std_logic_vector(54, 8),
23960 => conv_std_logic_vector(55, 8),
23961 => conv_std_logic_vector(55, 8),
23962 => conv_std_logic_vector(55, 8),
23963 => conv_std_logic_vector(56, 8),
23964 => conv_std_logic_vector(56, 8),
23965 => conv_std_logic_vector(57, 8),
23966 => conv_std_logic_vector(57, 8),
23967 => conv_std_logic_vector(57, 8),
23968 => conv_std_logic_vector(58, 8),
23969 => conv_std_logic_vector(58, 8),
23970 => conv_std_logic_vector(58, 8),
23971 => conv_std_logic_vector(59, 8),
23972 => conv_std_logic_vector(59, 8),
23973 => conv_std_logic_vector(59, 8),
23974 => conv_std_logic_vector(60, 8),
23975 => conv_std_logic_vector(60, 8),
23976 => conv_std_logic_vector(61, 8),
23977 => conv_std_logic_vector(61, 8),
23978 => conv_std_logic_vector(61, 8),
23979 => conv_std_logic_vector(62, 8),
23980 => conv_std_logic_vector(62, 8),
23981 => conv_std_logic_vector(62, 8),
23982 => conv_std_logic_vector(63, 8),
23983 => conv_std_logic_vector(63, 8),
23984 => conv_std_logic_vector(63, 8),
23985 => conv_std_logic_vector(64, 8),
23986 => conv_std_logic_vector(64, 8),
23987 => conv_std_logic_vector(65, 8),
23988 => conv_std_logic_vector(65, 8),
23989 => conv_std_logic_vector(65, 8),
23990 => conv_std_logic_vector(66, 8),
23991 => conv_std_logic_vector(66, 8),
23992 => conv_std_logic_vector(66, 8),
23993 => conv_std_logic_vector(67, 8),
23994 => conv_std_logic_vector(67, 8),
23995 => conv_std_logic_vector(67, 8),
23996 => conv_std_logic_vector(68, 8),
23997 => conv_std_logic_vector(68, 8),
23998 => conv_std_logic_vector(69, 8),
23999 => conv_std_logic_vector(69, 8),
24000 => conv_std_logic_vector(69, 8),
24001 => conv_std_logic_vector(70, 8),
24002 => conv_std_logic_vector(70, 8),
24003 => conv_std_logic_vector(70, 8),
24004 => conv_std_logic_vector(71, 8),
24005 => conv_std_logic_vector(71, 8),
24006 => conv_std_logic_vector(71, 8),
24007 => conv_std_logic_vector(72, 8),
24008 => conv_std_logic_vector(72, 8),
24009 => conv_std_logic_vector(73, 8),
24010 => conv_std_logic_vector(73, 8),
24011 => conv_std_logic_vector(73, 8),
24012 => conv_std_logic_vector(74, 8),
24013 => conv_std_logic_vector(74, 8),
24014 => conv_std_logic_vector(74, 8),
24015 => conv_std_logic_vector(75, 8),
24016 => conv_std_logic_vector(75, 8),
24017 => conv_std_logic_vector(75, 8),
24018 => conv_std_logic_vector(76, 8),
24019 => conv_std_logic_vector(76, 8),
24020 => conv_std_logic_vector(77, 8),
24021 => conv_std_logic_vector(77, 8),
24022 => conv_std_logic_vector(77, 8),
24023 => conv_std_logic_vector(78, 8),
24024 => conv_std_logic_vector(78, 8),
24025 => conv_std_logic_vector(78, 8),
24026 => conv_std_logic_vector(79, 8),
24027 => conv_std_logic_vector(79, 8),
24028 => conv_std_logic_vector(79, 8),
24029 => conv_std_logic_vector(80, 8),
24030 => conv_std_logic_vector(80, 8),
24031 => conv_std_logic_vector(81, 8),
24032 => conv_std_logic_vector(81, 8),
24033 => conv_std_logic_vector(81, 8),
24034 => conv_std_logic_vector(82, 8),
24035 => conv_std_logic_vector(82, 8),
24036 => conv_std_logic_vector(82, 8),
24037 => conv_std_logic_vector(83, 8),
24038 => conv_std_logic_vector(83, 8),
24039 => conv_std_logic_vector(83, 8),
24040 => conv_std_logic_vector(84, 8),
24041 => conv_std_logic_vector(84, 8),
24042 => conv_std_logic_vector(85, 8),
24043 => conv_std_logic_vector(85, 8),
24044 => conv_std_logic_vector(85, 8),
24045 => conv_std_logic_vector(86, 8),
24046 => conv_std_logic_vector(86, 8),
24047 => conv_std_logic_vector(86, 8),
24048 => conv_std_logic_vector(87, 8),
24049 => conv_std_logic_vector(87, 8),
24050 => conv_std_logic_vector(87, 8),
24051 => conv_std_logic_vector(88, 8),
24052 => conv_std_logic_vector(88, 8),
24053 => conv_std_logic_vector(89, 8),
24054 => conv_std_logic_vector(89, 8),
24055 => conv_std_logic_vector(89, 8),
24056 => conv_std_logic_vector(90, 8),
24057 => conv_std_logic_vector(90, 8),
24058 => conv_std_logic_vector(90, 8),
24059 => conv_std_logic_vector(91, 8),
24060 => conv_std_logic_vector(91, 8),
24061 => conv_std_logic_vector(91, 8),
24062 => conv_std_logic_vector(92, 8),
24063 => conv_std_logic_vector(92, 8),
24064 => conv_std_logic_vector(0, 8),
24065 => conv_std_logic_vector(0, 8),
24066 => conv_std_logic_vector(0, 8),
24067 => conv_std_logic_vector(1, 8),
24068 => conv_std_logic_vector(1, 8),
24069 => conv_std_logic_vector(1, 8),
24070 => conv_std_logic_vector(2, 8),
24071 => conv_std_logic_vector(2, 8),
24072 => conv_std_logic_vector(2, 8),
24073 => conv_std_logic_vector(3, 8),
24074 => conv_std_logic_vector(3, 8),
24075 => conv_std_logic_vector(4, 8),
24076 => conv_std_logic_vector(4, 8),
24077 => conv_std_logic_vector(4, 8),
24078 => conv_std_logic_vector(5, 8),
24079 => conv_std_logic_vector(5, 8),
24080 => conv_std_logic_vector(5, 8),
24081 => conv_std_logic_vector(6, 8),
24082 => conv_std_logic_vector(6, 8),
24083 => conv_std_logic_vector(6, 8),
24084 => conv_std_logic_vector(7, 8),
24085 => conv_std_logic_vector(7, 8),
24086 => conv_std_logic_vector(8, 8),
24087 => conv_std_logic_vector(8, 8),
24088 => conv_std_logic_vector(8, 8),
24089 => conv_std_logic_vector(9, 8),
24090 => conv_std_logic_vector(9, 8),
24091 => conv_std_logic_vector(9, 8),
24092 => conv_std_logic_vector(10, 8),
24093 => conv_std_logic_vector(10, 8),
24094 => conv_std_logic_vector(11, 8),
24095 => conv_std_logic_vector(11, 8),
24096 => conv_std_logic_vector(11, 8),
24097 => conv_std_logic_vector(12, 8),
24098 => conv_std_logic_vector(12, 8),
24099 => conv_std_logic_vector(12, 8),
24100 => conv_std_logic_vector(13, 8),
24101 => conv_std_logic_vector(13, 8),
24102 => conv_std_logic_vector(13, 8),
24103 => conv_std_logic_vector(14, 8),
24104 => conv_std_logic_vector(14, 8),
24105 => conv_std_logic_vector(15, 8),
24106 => conv_std_logic_vector(15, 8),
24107 => conv_std_logic_vector(15, 8),
24108 => conv_std_logic_vector(16, 8),
24109 => conv_std_logic_vector(16, 8),
24110 => conv_std_logic_vector(16, 8),
24111 => conv_std_logic_vector(17, 8),
24112 => conv_std_logic_vector(17, 8),
24113 => conv_std_logic_vector(17, 8),
24114 => conv_std_logic_vector(18, 8),
24115 => conv_std_logic_vector(18, 8),
24116 => conv_std_logic_vector(19, 8),
24117 => conv_std_logic_vector(19, 8),
24118 => conv_std_logic_vector(19, 8),
24119 => conv_std_logic_vector(20, 8),
24120 => conv_std_logic_vector(20, 8),
24121 => conv_std_logic_vector(20, 8),
24122 => conv_std_logic_vector(21, 8),
24123 => conv_std_logic_vector(21, 8),
24124 => conv_std_logic_vector(22, 8),
24125 => conv_std_logic_vector(22, 8),
24126 => conv_std_logic_vector(22, 8),
24127 => conv_std_logic_vector(23, 8),
24128 => conv_std_logic_vector(23, 8),
24129 => conv_std_logic_vector(23, 8),
24130 => conv_std_logic_vector(24, 8),
24131 => conv_std_logic_vector(24, 8),
24132 => conv_std_logic_vector(24, 8),
24133 => conv_std_logic_vector(25, 8),
24134 => conv_std_logic_vector(25, 8),
24135 => conv_std_logic_vector(26, 8),
24136 => conv_std_logic_vector(26, 8),
24137 => conv_std_logic_vector(26, 8),
24138 => conv_std_logic_vector(27, 8),
24139 => conv_std_logic_vector(27, 8),
24140 => conv_std_logic_vector(27, 8),
24141 => conv_std_logic_vector(28, 8),
24142 => conv_std_logic_vector(28, 8),
24143 => conv_std_logic_vector(29, 8),
24144 => conv_std_logic_vector(29, 8),
24145 => conv_std_logic_vector(29, 8),
24146 => conv_std_logic_vector(30, 8),
24147 => conv_std_logic_vector(30, 8),
24148 => conv_std_logic_vector(30, 8),
24149 => conv_std_logic_vector(31, 8),
24150 => conv_std_logic_vector(31, 8),
24151 => conv_std_logic_vector(31, 8),
24152 => conv_std_logic_vector(32, 8),
24153 => conv_std_logic_vector(32, 8),
24154 => conv_std_logic_vector(33, 8),
24155 => conv_std_logic_vector(33, 8),
24156 => conv_std_logic_vector(33, 8),
24157 => conv_std_logic_vector(34, 8),
24158 => conv_std_logic_vector(34, 8),
24159 => conv_std_logic_vector(34, 8),
24160 => conv_std_logic_vector(35, 8),
24161 => conv_std_logic_vector(35, 8),
24162 => conv_std_logic_vector(35, 8),
24163 => conv_std_logic_vector(36, 8),
24164 => conv_std_logic_vector(36, 8),
24165 => conv_std_logic_vector(37, 8),
24166 => conv_std_logic_vector(37, 8),
24167 => conv_std_logic_vector(37, 8),
24168 => conv_std_logic_vector(38, 8),
24169 => conv_std_logic_vector(38, 8),
24170 => conv_std_logic_vector(38, 8),
24171 => conv_std_logic_vector(39, 8),
24172 => conv_std_logic_vector(39, 8),
24173 => conv_std_logic_vector(40, 8),
24174 => conv_std_logic_vector(40, 8),
24175 => conv_std_logic_vector(40, 8),
24176 => conv_std_logic_vector(41, 8),
24177 => conv_std_logic_vector(41, 8),
24178 => conv_std_logic_vector(41, 8),
24179 => conv_std_logic_vector(42, 8),
24180 => conv_std_logic_vector(42, 8),
24181 => conv_std_logic_vector(42, 8),
24182 => conv_std_logic_vector(43, 8),
24183 => conv_std_logic_vector(43, 8),
24184 => conv_std_logic_vector(44, 8),
24185 => conv_std_logic_vector(44, 8),
24186 => conv_std_logic_vector(44, 8),
24187 => conv_std_logic_vector(45, 8),
24188 => conv_std_logic_vector(45, 8),
24189 => conv_std_logic_vector(45, 8),
24190 => conv_std_logic_vector(46, 8),
24191 => conv_std_logic_vector(46, 8),
24192 => conv_std_logic_vector(47, 8),
24193 => conv_std_logic_vector(47, 8),
24194 => conv_std_logic_vector(47, 8),
24195 => conv_std_logic_vector(48, 8),
24196 => conv_std_logic_vector(48, 8),
24197 => conv_std_logic_vector(48, 8),
24198 => conv_std_logic_vector(49, 8),
24199 => conv_std_logic_vector(49, 8),
24200 => conv_std_logic_vector(49, 8),
24201 => conv_std_logic_vector(50, 8),
24202 => conv_std_logic_vector(50, 8),
24203 => conv_std_logic_vector(51, 8),
24204 => conv_std_logic_vector(51, 8),
24205 => conv_std_logic_vector(51, 8),
24206 => conv_std_logic_vector(52, 8),
24207 => conv_std_logic_vector(52, 8),
24208 => conv_std_logic_vector(52, 8),
24209 => conv_std_logic_vector(53, 8),
24210 => conv_std_logic_vector(53, 8),
24211 => conv_std_logic_vector(53, 8),
24212 => conv_std_logic_vector(54, 8),
24213 => conv_std_logic_vector(54, 8),
24214 => conv_std_logic_vector(55, 8),
24215 => conv_std_logic_vector(55, 8),
24216 => conv_std_logic_vector(55, 8),
24217 => conv_std_logic_vector(56, 8),
24218 => conv_std_logic_vector(56, 8),
24219 => conv_std_logic_vector(56, 8),
24220 => conv_std_logic_vector(57, 8),
24221 => conv_std_logic_vector(57, 8),
24222 => conv_std_logic_vector(58, 8),
24223 => conv_std_logic_vector(58, 8),
24224 => conv_std_logic_vector(58, 8),
24225 => conv_std_logic_vector(59, 8),
24226 => conv_std_logic_vector(59, 8),
24227 => conv_std_logic_vector(59, 8),
24228 => conv_std_logic_vector(60, 8),
24229 => conv_std_logic_vector(60, 8),
24230 => conv_std_logic_vector(60, 8),
24231 => conv_std_logic_vector(61, 8),
24232 => conv_std_logic_vector(61, 8),
24233 => conv_std_logic_vector(62, 8),
24234 => conv_std_logic_vector(62, 8),
24235 => conv_std_logic_vector(62, 8),
24236 => conv_std_logic_vector(63, 8),
24237 => conv_std_logic_vector(63, 8),
24238 => conv_std_logic_vector(63, 8),
24239 => conv_std_logic_vector(64, 8),
24240 => conv_std_logic_vector(64, 8),
24241 => conv_std_logic_vector(64, 8),
24242 => conv_std_logic_vector(65, 8),
24243 => conv_std_logic_vector(65, 8),
24244 => conv_std_logic_vector(66, 8),
24245 => conv_std_logic_vector(66, 8),
24246 => conv_std_logic_vector(66, 8),
24247 => conv_std_logic_vector(67, 8),
24248 => conv_std_logic_vector(67, 8),
24249 => conv_std_logic_vector(67, 8),
24250 => conv_std_logic_vector(68, 8),
24251 => conv_std_logic_vector(68, 8),
24252 => conv_std_logic_vector(69, 8),
24253 => conv_std_logic_vector(69, 8),
24254 => conv_std_logic_vector(69, 8),
24255 => conv_std_logic_vector(70, 8),
24256 => conv_std_logic_vector(70, 8),
24257 => conv_std_logic_vector(70, 8),
24258 => conv_std_logic_vector(71, 8),
24259 => conv_std_logic_vector(71, 8),
24260 => conv_std_logic_vector(71, 8),
24261 => conv_std_logic_vector(72, 8),
24262 => conv_std_logic_vector(72, 8),
24263 => conv_std_logic_vector(73, 8),
24264 => conv_std_logic_vector(73, 8),
24265 => conv_std_logic_vector(73, 8),
24266 => conv_std_logic_vector(74, 8),
24267 => conv_std_logic_vector(74, 8),
24268 => conv_std_logic_vector(74, 8),
24269 => conv_std_logic_vector(75, 8),
24270 => conv_std_logic_vector(75, 8),
24271 => conv_std_logic_vector(76, 8),
24272 => conv_std_logic_vector(76, 8),
24273 => conv_std_logic_vector(76, 8),
24274 => conv_std_logic_vector(77, 8),
24275 => conv_std_logic_vector(77, 8),
24276 => conv_std_logic_vector(77, 8),
24277 => conv_std_logic_vector(78, 8),
24278 => conv_std_logic_vector(78, 8),
24279 => conv_std_logic_vector(78, 8),
24280 => conv_std_logic_vector(79, 8),
24281 => conv_std_logic_vector(79, 8),
24282 => conv_std_logic_vector(80, 8),
24283 => conv_std_logic_vector(80, 8),
24284 => conv_std_logic_vector(80, 8),
24285 => conv_std_logic_vector(81, 8),
24286 => conv_std_logic_vector(81, 8),
24287 => conv_std_logic_vector(81, 8),
24288 => conv_std_logic_vector(82, 8),
24289 => conv_std_logic_vector(82, 8),
24290 => conv_std_logic_vector(82, 8),
24291 => conv_std_logic_vector(83, 8),
24292 => conv_std_logic_vector(83, 8),
24293 => conv_std_logic_vector(84, 8),
24294 => conv_std_logic_vector(84, 8),
24295 => conv_std_logic_vector(84, 8),
24296 => conv_std_logic_vector(85, 8),
24297 => conv_std_logic_vector(85, 8),
24298 => conv_std_logic_vector(85, 8),
24299 => conv_std_logic_vector(86, 8),
24300 => conv_std_logic_vector(86, 8),
24301 => conv_std_logic_vector(87, 8),
24302 => conv_std_logic_vector(87, 8),
24303 => conv_std_logic_vector(87, 8),
24304 => conv_std_logic_vector(88, 8),
24305 => conv_std_logic_vector(88, 8),
24306 => conv_std_logic_vector(88, 8),
24307 => conv_std_logic_vector(89, 8),
24308 => conv_std_logic_vector(89, 8),
24309 => conv_std_logic_vector(89, 8),
24310 => conv_std_logic_vector(90, 8),
24311 => conv_std_logic_vector(90, 8),
24312 => conv_std_logic_vector(91, 8),
24313 => conv_std_logic_vector(91, 8),
24314 => conv_std_logic_vector(91, 8),
24315 => conv_std_logic_vector(92, 8),
24316 => conv_std_logic_vector(92, 8),
24317 => conv_std_logic_vector(92, 8),
24318 => conv_std_logic_vector(93, 8),
24319 => conv_std_logic_vector(93, 8),
24320 => conv_std_logic_vector(0, 8),
24321 => conv_std_logic_vector(0, 8),
24322 => conv_std_logic_vector(0, 8),
24323 => conv_std_logic_vector(1, 8),
24324 => conv_std_logic_vector(1, 8),
24325 => conv_std_logic_vector(1, 8),
24326 => conv_std_logic_vector(2, 8),
24327 => conv_std_logic_vector(2, 8),
24328 => conv_std_logic_vector(2, 8),
24329 => conv_std_logic_vector(3, 8),
24330 => conv_std_logic_vector(3, 8),
24331 => conv_std_logic_vector(4, 8),
24332 => conv_std_logic_vector(4, 8),
24333 => conv_std_logic_vector(4, 8),
24334 => conv_std_logic_vector(5, 8),
24335 => conv_std_logic_vector(5, 8),
24336 => conv_std_logic_vector(5, 8),
24337 => conv_std_logic_vector(6, 8),
24338 => conv_std_logic_vector(6, 8),
24339 => conv_std_logic_vector(7, 8),
24340 => conv_std_logic_vector(7, 8),
24341 => conv_std_logic_vector(7, 8),
24342 => conv_std_logic_vector(8, 8),
24343 => conv_std_logic_vector(8, 8),
24344 => conv_std_logic_vector(8, 8),
24345 => conv_std_logic_vector(9, 8),
24346 => conv_std_logic_vector(9, 8),
24347 => conv_std_logic_vector(10, 8),
24348 => conv_std_logic_vector(10, 8),
24349 => conv_std_logic_vector(10, 8),
24350 => conv_std_logic_vector(11, 8),
24351 => conv_std_logic_vector(11, 8),
24352 => conv_std_logic_vector(11, 8),
24353 => conv_std_logic_vector(12, 8),
24354 => conv_std_logic_vector(12, 8),
24355 => conv_std_logic_vector(12, 8),
24356 => conv_std_logic_vector(13, 8),
24357 => conv_std_logic_vector(13, 8),
24358 => conv_std_logic_vector(14, 8),
24359 => conv_std_logic_vector(14, 8),
24360 => conv_std_logic_vector(14, 8),
24361 => conv_std_logic_vector(15, 8),
24362 => conv_std_logic_vector(15, 8),
24363 => conv_std_logic_vector(15, 8),
24364 => conv_std_logic_vector(16, 8),
24365 => conv_std_logic_vector(16, 8),
24366 => conv_std_logic_vector(17, 8),
24367 => conv_std_logic_vector(17, 8),
24368 => conv_std_logic_vector(17, 8),
24369 => conv_std_logic_vector(18, 8),
24370 => conv_std_logic_vector(18, 8),
24371 => conv_std_logic_vector(18, 8),
24372 => conv_std_logic_vector(19, 8),
24373 => conv_std_logic_vector(19, 8),
24374 => conv_std_logic_vector(20, 8),
24375 => conv_std_logic_vector(20, 8),
24376 => conv_std_logic_vector(20, 8),
24377 => conv_std_logic_vector(21, 8),
24378 => conv_std_logic_vector(21, 8),
24379 => conv_std_logic_vector(21, 8),
24380 => conv_std_logic_vector(22, 8),
24381 => conv_std_logic_vector(22, 8),
24382 => conv_std_logic_vector(23, 8),
24383 => conv_std_logic_vector(23, 8),
24384 => conv_std_logic_vector(23, 8),
24385 => conv_std_logic_vector(24, 8),
24386 => conv_std_logic_vector(24, 8),
24387 => conv_std_logic_vector(24, 8),
24388 => conv_std_logic_vector(25, 8),
24389 => conv_std_logic_vector(25, 8),
24390 => conv_std_logic_vector(25, 8),
24391 => conv_std_logic_vector(26, 8),
24392 => conv_std_logic_vector(26, 8),
24393 => conv_std_logic_vector(27, 8),
24394 => conv_std_logic_vector(27, 8),
24395 => conv_std_logic_vector(27, 8),
24396 => conv_std_logic_vector(28, 8),
24397 => conv_std_logic_vector(28, 8),
24398 => conv_std_logic_vector(28, 8),
24399 => conv_std_logic_vector(29, 8),
24400 => conv_std_logic_vector(29, 8),
24401 => conv_std_logic_vector(30, 8),
24402 => conv_std_logic_vector(30, 8),
24403 => conv_std_logic_vector(30, 8),
24404 => conv_std_logic_vector(31, 8),
24405 => conv_std_logic_vector(31, 8),
24406 => conv_std_logic_vector(31, 8),
24407 => conv_std_logic_vector(32, 8),
24408 => conv_std_logic_vector(32, 8),
24409 => conv_std_logic_vector(33, 8),
24410 => conv_std_logic_vector(33, 8),
24411 => conv_std_logic_vector(33, 8),
24412 => conv_std_logic_vector(34, 8),
24413 => conv_std_logic_vector(34, 8),
24414 => conv_std_logic_vector(34, 8),
24415 => conv_std_logic_vector(35, 8),
24416 => conv_std_logic_vector(35, 8),
24417 => conv_std_logic_vector(35, 8),
24418 => conv_std_logic_vector(36, 8),
24419 => conv_std_logic_vector(36, 8),
24420 => conv_std_logic_vector(37, 8),
24421 => conv_std_logic_vector(37, 8),
24422 => conv_std_logic_vector(37, 8),
24423 => conv_std_logic_vector(38, 8),
24424 => conv_std_logic_vector(38, 8),
24425 => conv_std_logic_vector(38, 8),
24426 => conv_std_logic_vector(39, 8),
24427 => conv_std_logic_vector(39, 8),
24428 => conv_std_logic_vector(40, 8),
24429 => conv_std_logic_vector(40, 8),
24430 => conv_std_logic_vector(40, 8),
24431 => conv_std_logic_vector(41, 8),
24432 => conv_std_logic_vector(41, 8),
24433 => conv_std_logic_vector(41, 8),
24434 => conv_std_logic_vector(42, 8),
24435 => conv_std_logic_vector(42, 8),
24436 => conv_std_logic_vector(43, 8),
24437 => conv_std_logic_vector(43, 8),
24438 => conv_std_logic_vector(43, 8),
24439 => conv_std_logic_vector(44, 8),
24440 => conv_std_logic_vector(44, 8),
24441 => conv_std_logic_vector(44, 8),
24442 => conv_std_logic_vector(45, 8),
24443 => conv_std_logic_vector(45, 8),
24444 => conv_std_logic_vector(46, 8),
24445 => conv_std_logic_vector(46, 8),
24446 => conv_std_logic_vector(46, 8),
24447 => conv_std_logic_vector(47, 8),
24448 => conv_std_logic_vector(47, 8),
24449 => conv_std_logic_vector(47, 8),
24450 => conv_std_logic_vector(48, 8),
24451 => conv_std_logic_vector(48, 8),
24452 => conv_std_logic_vector(48, 8),
24453 => conv_std_logic_vector(49, 8),
24454 => conv_std_logic_vector(49, 8),
24455 => conv_std_logic_vector(50, 8),
24456 => conv_std_logic_vector(50, 8),
24457 => conv_std_logic_vector(50, 8),
24458 => conv_std_logic_vector(51, 8),
24459 => conv_std_logic_vector(51, 8),
24460 => conv_std_logic_vector(51, 8),
24461 => conv_std_logic_vector(52, 8),
24462 => conv_std_logic_vector(52, 8),
24463 => conv_std_logic_vector(53, 8),
24464 => conv_std_logic_vector(53, 8),
24465 => conv_std_logic_vector(53, 8),
24466 => conv_std_logic_vector(54, 8),
24467 => conv_std_logic_vector(54, 8),
24468 => conv_std_logic_vector(54, 8),
24469 => conv_std_logic_vector(55, 8),
24470 => conv_std_logic_vector(55, 8),
24471 => conv_std_logic_vector(56, 8),
24472 => conv_std_logic_vector(56, 8),
24473 => conv_std_logic_vector(56, 8),
24474 => conv_std_logic_vector(57, 8),
24475 => conv_std_logic_vector(57, 8),
24476 => conv_std_logic_vector(57, 8),
24477 => conv_std_logic_vector(58, 8),
24478 => conv_std_logic_vector(58, 8),
24479 => conv_std_logic_vector(59, 8),
24480 => conv_std_logic_vector(59, 8),
24481 => conv_std_logic_vector(59, 8),
24482 => conv_std_logic_vector(60, 8),
24483 => conv_std_logic_vector(60, 8),
24484 => conv_std_logic_vector(60, 8),
24485 => conv_std_logic_vector(61, 8),
24486 => conv_std_logic_vector(61, 8),
24487 => conv_std_logic_vector(61, 8),
24488 => conv_std_logic_vector(62, 8),
24489 => conv_std_logic_vector(62, 8),
24490 => conv_std_logic_vector(63, 8),
24491 => conv_std_logic_vector(63, 8),
24492 => conv_std_logic_vector(63, 8),
24493 => conv_std_logic_vector(64, 8),
24494 => conv_std_logic_vector(64, 8),
24495 => conv_std_logic_vector(64, 8),
24496 => conv_std_logic_vector(65, 8),
24497 => conv_std_logic_vector(65, 8),
24498 => conv_std_logic_vector(66, 8),
24499 => conv_std_logic_vector(66, 8),
24500 => conv_std_logic_vector(66, 8),
24501 => conv_std_logic_vector(67, 8),
24502 => conv_std_logic_vector(67, 8),
24503 => conv_std_logic_vector(67, 8),
24504 => conv_std_logic_vector(68, 8),
24505 => conv_std_logic_vector(68, 8),
24506 => conv_std_logic_vector(69, 8),
24507 => conv_std_logic_vector(69, 8),
24508 => conv_std_logic_vector(69, 8),
24509 => conv_std_logic_vector(70, 8),
24510 => conv_std_logic_vector(70, 8),
24511 => conv_std_logic_vector(70, 8),
24512 => conv_std_logic_vector(71, 8),
24513 => conv_std_logic_vector(71, 8),
24514 => conv_std_logic_vector(71, 8),
24515 => conv_std_logic_vector(72, 8),
24516 => conv_std_logic_vector(72, 8),
24517 => conv_std_logic_vector(73, 8),
24518 => conv_std_logic_vector(73, 8),
24519 => conv_std_logic_vector(73, 8),
24520 => conv_std_logic_vector(74, 8),
24521 => conv_std_logic_vector(74, 8),
24522 => conv_std_logic_vector(74, 8),
24523 => conv_std_logic_vector(75, 8),
24524 => conv_std_logic_vector(75, 8),
24525 => conv_std_logic_vector(76, 8),
24526 => conv_std_logic_vector(76, 8),
24527 => conv_std_logic_vector(76, 8),
24528 => conv_std_logic_vector(77, 8),
24529 => conv_std_logic_vector(77, 8),
24530 => conv_std_logic_vector(77, 8),
24531 => conv_std_logic_vector(78, 8),
24532 => conv_std_logic_vector(78, 8),
24533 => conv_std_logic_vector(79, 8),
24534 => conv_std_logic_vector(79, 8),
24535 => conv_std_logic_vector(79, 8),
24536 => conv_std_logic_vector(80, 8),
24537 => conv_std_logic_vector(80, 8),
24538 => conv_std_logic_vector(80, 8),
24539 => conv_std_logic_vector(81, 8),
24540 => conv_std_logic_vector(81, 8),
24541 => conv_std_logic_vector(82, 8),
24542 => conv_std_logic_vector(82, 8),
24543 => conv_std_logic_vector(82, 8),
24544 => conv_std_logic_vector(83, 8),
24545 => conv_std_logic_vector(83, 8),
24546 => conv_std_logic_vector(83, 8),
24547 => conv_std_logic_vector(84, 8),
24548 => conv_std_logic_vector(84, 8),
24549 => conv_std_logic_vector(84, 8),
24550 => conv_std_logic_vector(85, 8),
24551 => conv_std_logic_vector(85, 8),
24552 => conv_std_logic_vector(86, 8),
24553 => conv_std_logic_vector(86, 8),
24554 => conv_std_logic_vector(86, 8),
24555 => conv_std_logic_vector(87, 8),
24556 => conv_std_logic_vector(87, 8),
24557 => conv_std_logic_vector(87, 8),
24558 => conv_std_logic_vector(88, 8),
24559 => conv_std_logic_vector(88, 8),
24560 => conv_std_logic_vector(89, 8),
24561 => conv_std_logic_vector(89, 8),
24562 => conv_std_logic_vector(89, 8),
24563 => conv_std_logic_vector(90, 8),
24564 => conv_std_logic_vector(90, 8),
24565 => conv_std_logic_vector(90, 8),
24566 => conv_std_logic_vector(91, 8),
24567 => conv_std_logic_vector(91, 8),
24568 => conv_std_logic_vector(92, 8),
24569 => conv_std_logic_vector(92, 8),
24570 => conv_std_logic_vector(92, 8),
24571 => conv_std_logic_vector(93, 8),
24572 => conv_std_logic_vector(93, 8),
24573 => conv_std_logic_vector(93, 8),
24574 => conv_std_logic_vector(94, 8),
24575 => conv_std_logic_vector(94, 8),
24576 => conv_std_logic_vector(0, 8),
24577 => conv_std_logic_vector(0, 8),
24578 => conv_std_logic_vector(0, 8),
24579 => conv_std_logic_vector(1, 8),
24580 => conv_std_logic_vector(1, 8),
24581 => conv_std_logic_vector(1, 8),
24582 => conv_std_logic_vector(2, 8),
24583 => conv_std_logic_vector(2, 8),
24584 => conv_std_logic_vector(3, 8),
24585 => conv_std_logic_vector(3, 8),
24586 => conv_std_logic_vector(3, 8),
24587 => conv_std_logic_vector(4, 8),
24588 => conv_std_logic_vector(4, 8),
24589 => conv_std_logic_vector(4, 8),
24590 => conv_std_logic_vector(5, 8),
24591 => conv_std_logic_vector(5, 8),
24592 => conv_std_logic_vector(6, 8),
24593 => conv_std_logic_vector(6, 8),
24594 => conv_std_logic_vector(6, 8),
24595 => conv_std_logic_vector(7, 8),
24596 => conv_std_logic_vector(7, 8),
24597 => conv_std_logic_vector(7, 8),
24598 => conv_std_logic_vector(8, 8),
24599 => conv_std_logic_vector(8, 8),
24600 => conv_std_logic_vector(9, 8),
24601 => conv_std_logic_vector(9, 8),
24602 => conv_std_logic_vector(9, 8),
24603 => conv_std_logic_vector(10, 8),
24604 => conv_std_logic_vector(10, 8),
24605 => conv_std_logic_vector(10, 8),
24606 => conv_std_logic_vector(11, 8),
24607 => conv_std_logic_vector(11, 8),
24608 => conv_std_logic_vector(12, 8),
24609 => conv_std_logic_vector(12, 8),
24610 => conv_std_logic_vector(12, 8),
24611 => conv_std_logic_vector(13, 8),
24612 => conv_std_logic_vector(13, 8),
24613 => conv_std_logic_vector(13, 8),
24614 => conv_std_logic_vector(14, 8),
24615 => conv_std_logic_vector(14, 8),
24616 => conv_std_logic_vector(15, 8),
24617 => conv_std_logic_vector(15, 8),
24618 => conv_std_logic_vector(15, 8),
24619 => conv_std_logic_vector(16, 8),
24620 => conv_std_logic_vector(16, 8),
24621 => conv_std_logic_vector(16, 8),
24622 => conv_std_logic_vector(17, 8),
24623 => conv_std_logic_vector(17, 8),
24624 => conv_std_logic_vector(18, 8),
24625 => conv_std_logic_vector(18, 8),
24626 => conv_std_logic_vector(18, 8),
24627 => conv_std_logic_vector(19, 8),
24628 => conv_std_logic_vector(19, 8),
24629 => conv_std_logic_vector(19, 8),
24630 => conv_std_logic_vector(20, 8),
24631 => conv_std_logic_vector(20, 8),
24632 => conv_std_logic_vector(21, 8),
24633 => conv_std_logic_vector(21, 8),
24634 => conv_std_logic_vector(21, 8),
24635 => conv_std_logic_vector(22, 8),
24636 => conv_std_logic_vector(22, 8),
24637 => conv_std_logic_vector(22, 8),
24638 => conv_std_logic_vector(23, 8),
24639 => conv_std_logic_vector(23, 8),
24640 => conv_std_logic_vector(24, 8),
24641 => conv_std_logic_vector(24, 8),
24642 => conv_std_logic_vector(24, 8),
24643 => conv_std_logic_vector(25, 8),
24644 => conv_std_logic_vector(25, 8),
24645 => conv_std_logic_vector(25, 8),
24646 => conv_std_logic_vector(26, 8),
24647 => conv_std_logic_vector(26, 8),
24648 => conv_std_logic_vector(27, 8),
24649 => conv_std_logic_vector(27, 8),
24650 => conv_std_logic_vector(27, 8),
24651 => conv_std_logic_vector(28, 8),
24652 => conv_std_logic_vector(28, 8),
24653 => conv_std_logic_vector(28, 8),
24654 => conv_std_logic_vector(29, 8),
24655 => conv_std_logic_vector(29, 8),
24656 => conv_std_logic_vector(30, 8),
24657 => conv_std_logic_vector(30, 8),
24658 => conv_std_logic_vector(30, 8),
24659 => conv_std_logic_vector(31, 8),
24660 => conv_std_logic_vector(31, 8),
24661 => conv_std_logic_vector(31, 8),
24662 => conv_std_logic_vector(32, 8),
24663 => conv_std_logic_vector(32, 8),
24664 => conv_std_logic_vector(33, 8),
24665 => conv_std_logic_vector(33, 8),
24666 => conv_std_logic_vector(33, 8),
24667 => conv_std_logic_vector(34, 8),
24668 => conv_std_logic_vector(34, 8),
24669 => conv_std_logic_vector(34, 8),
24670 => conv_std_logic_vector(35, 8),
24671 => conv_std_logic_vector(35, 8),
24672 => conv_std_logic_vector(36, 8),
24673 => conv_std_logic_vector(36, 8),
24674 => conv_std_logic_vector(36, 8),
24675 => conv_std_logic_vector(37, 8),
24676 => conv_std_logic_vector(37, 8),
24677 => conv_std_logic_vector(37, 8),
24678 => conv_std_logic_vector(38, 8),
24679 => conv_std_logic_vector(38, 8),
24680 => conv_std_logic_vector(39, 8),
24681 => conv_std_logic_vector(39, 8),
24682 => conv_std_logic_vector(39, 8),
24683 => conv_std_logic_vector(40, 8),
24684 => conv_std_logic_vector(40, 8),
24685 => conv_std_logic_vector(40, 8),
24686 => conv_std_logic_vector(41, 8),
24687 => conv_std_logic_vector(41, 8),
24688 => conv_std_logic_vector(42, 8),
24689 => conv_std_logic_vector(42, 8),
24690 => conv_std_logic_vector(42, 8),
24691 => conv_std_logic_vector(43, 8),
24692 => conv_std_logic_vector(43, 8),
24693 => conv_std_logic_vector(43, 8),
24694 => conv_std_logic_vector(44, 8),
24695 => conv_std_logic_vector(44, 8),
24696 => conv_std_logic_vector(45, 8),
24697 => conv_std_logic_vector(45, 8),
24698 => conv_std_logic_vector(45, 8),
24699 => conv_std_logic_vector(46, 8),
24700 => conv_std_logic_vector(46, 8),
24701 => conv_std_logic_vector(46, 8),
24702 => conv_std_logic_vector(47, 8),
24703 => conv_std_logic_vector(47, 8),
24704 => conv_std_logic_vector(48, 8),
24705 => conv_std_logic_vector(48, 8),
24706 => conv_std_logic_vector(48, 8),
24707 => conv_std_logic_vector(49, 8),
24708 => conv_std_logic_vector(49, 8),
24709 => conv_std_logic_vector(49, 8),
24710 => conv_std_logic_vector(50, 8),
24711 => conv_std_logic_vector(50, 8),
24712 => conv_std_logic_vector(51, 8),
24713 => conv_std_logic_vector(51, 8),
24714 => conv_std_logic_vector(51, 8),
24715 => conv_std_logic_vector(52, 8),
24716 => conv_std_logic_vector(52, 8),
24717 => conv_std_logic_vector(52, 8),
24718 => conv_std_logic_vector(53, 8),
24719 => conv_std_logic_vector(53, 8),
24720 => conv_std_logic_vector(54, 8),
24721 => conv_std_logic_vector(54, 8),
24722 => conv_std_logic_vector(54, 8),
24723 => conv_std_logic_vector(55, 8),
24724 => conv_std_logic_vector(55, 8),
24725 => conv_std_logic_vector(55, 8),
24726 => conv_std_logic_vector(56, 8),
24727 => conv_std_logic_vector(56, 8),
24728 => conv_std_logic_vector(57, 8),
24729 => conv_std_logic_vector(57, 8),
24730 => conv_std_logic_vector(57, 8),
24731 => conv_std_logic_vector(58, 8),
24732 => conv_std_logic_vector(58, 8),
24733 => conv_std_logic_vector(58, 8),
24734 => conv_std_logic_vector(59, 8),
24735 => conv_std_logic_vector(59, 8),
24736 => conv_std_logic_vector(60, 8),
24737 => conv_std_logic_vector(60, 8),
24738 => conv_std_logic_vector(60, 8),
24739 => conv_std_logic_vector(61, 8),
24740 => conv_std_logic_vector(61, 8),
24741 => conv_std_logic_vector(61, 8),
24742 => conv_std_logic_vector(62, 8),
24743 => conv_std_logic_vector(62, 8),
24744 => conv_std_logic_vector(63, 8),
24745 => conv_std_logic_vector(63, 8),
24746 => conv_std_logic_vector(63, 8),
24747 => conv_std_logic_vector(64, 8),
24748 => conv_std_logic_vector(64, 8),
24749 => conv_std_logic_vector(64, 8),
24750 => conv_std_logic_vector(65, 8),
24751 => conv_std_logic_vector(65, 8),
24752 => conv_std_logic_vector(66, 8),
24753 => conv_std_logic_vector(66, 8),
24754 => conv_std_logic_vector(66, 8),
24755 => conv_std_logic_vector(67, 8),
24756 => conv_std_logic_vector(67, 8),
24757 => conv_std_logic_vector(67, 8),
24758 => conv_std_logic_vector(68, 8),
24759 => conv_std_logic_vector(68, 8),
24760 => conv_std_logic_vector(69, 8),
24761 => conv_std_logic_vector(69, 8),
24762 => conv_std_logic_vector(69, 8),
24763 => conv_std_logic_vector(70, 8),
24764 => conv_std_logic_vector(70, 8),
24765 => conv_std_logic_vector(70, 8),
24766 => conv_std_logic_vector(71, 8),
24767 => conv_std_logic_vector(71, 8),
24768 => conv_std_logic_vector(72, 8),
24769 => conv_std_logic_vector(72, 8),
24770 => conv_std_logic_vector(72, 8),
24771 => conv_std_logic_vector(73, 8),
24772 => conv_std_logic_vector(73, 8),
24773 => conv_std_logic_vector(73, 8),
24774 => conv_std_logic_vector(74, 8),
24775 => conv_std_logic_vector(74, 8),
24776 => conv_std_logic_vector(75, 8),
24777 => conv_std_logic_vector(75, 8),
24778 => conv_std_logic_vector(75, 8),
24779 => conv_std_logic_vector(76, 8),
24780 => conv_std_logic_vector(76, 8),
24781 => conv_std_logic_vector(76, 8),
24782 => conv_std_logic_vector(77, 8),
24783 => conv_std_logic_vector(77, 8),
24784 => conv_std_logic_vector(78, 8),
24785 => conv_std_logic_vector(78, 8),
24786 => conv_std_logic_vector(78, 8),
24787 => conv_std_logic_vector(79, 8),
24788 => conv_std_logic_vector(79, 8),
24789 => conv_std_logic_vector(79, 8),
24790 => conv_std_logic_vector(80, 8),
24791 => conv_std_logic_vector(80, 8),
24792 => conv_std_logic_vector(81, 8),
24793 => conv_std_logic_vector(81, 8),
24794 => conv_std_logic_vector(81, 8),
24795 => conv_std_logic_vector(82, 8),
24796 => conv_std_logic_vector(82, 8),
24797 => conv_std_logic_vector(82, 8),
24798 => conv_std_logic_vector(83, 8),
24799 => conv_std_logic_vector(83, 8),
24800 => conv_std_logic_vector(84, 8),
24801 => conv_std_logic_vector(84, 8),
24802 => conv_std_logic_vector(84, 8),
24803 => conv_std_logic_vector(85, 8),
24804 => conv_std_logic_vector(85, 8),
24805 => conv_std_logic_vector(85, 8),
24806 => conv_std_logic_vector(86, 8),
24807 => conv_std_logic_vector(86, 8),
24808 => conv_std_logic_vector(87, 8),
24809 => conv_std_logic_vector(87, 8),
24810 => conv_std_logic_vector(87, 8),
24811 => conv_std_logic_vector(88, 8),
24812 => conv_std_logic_vector(88, 8),
24813 => conv_std_logic_vector(88, 8),
24814 => conv_std_logic_vector(89, 8),
24815 => conv_std_logic_vector(89, 8),
24816 => conv_std_logic_vector(90, 8),
24817 => conv_std_logic_vector(90, 8),
24818 => conv_std_logic_vector(90, 8),
24819 => conv_std_logic_vector(91, 8),
24820 => conv_std_logic_vector(91, 8),
24821 => conv_std_logic_vector(91, 8),
24822 => conv_std_logic_vector(92, 8),
24823 => conv_std_logic_vector(92, 8),
24824 => conv_std_logic_vector(93, 8),
24825 => conv_std_logic_vector(93, 8),
24826 => conv_std_logic_vector(93, 8),
24827 => conv_std_logic_vector(94, 8),
24828 => conv_std_logic_vector(94, 8),
24829 => conv_std_logic_vector(94, 8),
24830 => conv_std_logic_vector(95, 8),
24831 => conv_std_logic_vector(95, 8),
24832 => conv_std_logic_vector(0, 8),
24833 => conv_std_logic_vector(0, 8),
24834 => conv_std_logic_vector(0, 8),
24835 => conv_std_logic_vector(1, 8),
24836 => conv_std_logic_vector(1, 8),
24837 => conv_std_logic_vector(1, 8),
24838 => conv_std_logic_vector(2, 8),
24839 => conv_std_logic_vector(2, 8),
24840 => conv_std_logic_vector(3, 8),
24841 => conv_std_logic_vector(3, 8),
24842 => conv_std_logic_vector(3, 8),
24843 => conv_std_logic_vector(4, 8),
24844 => conv_std_logic_vector(4, 8),
24845 => conv_std_logic_vector(4, 8),
24846 => conv_std_logic_vector(5, 8),
24847 => conv_std_logic_vector(5, 8),
24848 => conv_std_logic_vector(6, 8),
24849 => conv_std_logic_vector(6, 8),
24850 => conv_std_logic_vector(6, 8),
24851 => conv_std_logic_vector(7, 8),
24852 => conv_std_logic_vector(7, 8),
24853 => conv_std_logic_vector(7, 8),
24854 => conv_std_logic_vector(8, 8),
24855 => conv_std_logic_vector(8, 8),
24856 => conv_std_logic_vector(9, 8),
24857 => conv_std_logic_vector(9, 8),
24858 => conv_std_logic_vector(9, 8),
24859 => conv_std_logic_vector(10, 8),
24860 => conv_std_logic_vector(10, 8),
24861 => conv_std_logic_vector(10, 8),
24862 => conv_std_logic_vector(11, 8),
24863 => conv_std_logic_vector(11, 8),
24864 => conv_std_logic_vector(12, 8),
24865 => conv_std_logic_vector(12, 8),
24866 => conv_std_logic_vector(12, 8),
24867 => conv_std_logic_vector(13, 8),
24868 => conv_std_logic_vector(13, 8),
24869 => conv_std_logic_vector(14, 8),
24870 => conv_std_logic_vector(14, 8),
24871 => conv_std_logic_vector(14, 8),
24872 => conv_std_logic_vector(15, 8),
24873 => conv_std_logic_vector(15, 8),
24874 => conv_std_logic_vector(15, 8),
24875 => conv_std_logic_vector(16, 8),
24876 => conv_std_logic_vector(16, 8),
24877 => conv_std_logic_vector(17, 8),
24878 => conv_std_logic_vector(17, 8),
24879 => conv_std_logic_vector(17, 8),
24880 => conv_std_logic_vector(18, 8),
24881 => conv_std_logic_vector(18, 8),
24882 => conv_std_logic_vector(18, 8),
24883 => conv_std_logic_vector(19, 8),
24884 => conv_std_logic_vector(19, 8),
24885 => conv_std_logic_vector(20, 8),
24886 => conv_std_logic_vector(20, 8),
24887 => conv_std_logic_vector(20, 8),
24888 => conv_std_logic_vector(21, 8),
24889 => conv_std_logic_vector(21, 8),
24890 => conv_std_logic_vector(21, 8),
24891 => conv_std_logic_vector(22, 8),
24892 => conv_std_logic_vector(22, 8),
24893 => conv_std_logic_vector(23, 8),
24894 => conv_std_logic_vector(23, 8),
24895 => conv_std_logic_vector(23, 8),
24896 => conv_std_logic_vector(24, 8),
24897 => conv_std_logic_vector(24, 8),
24898 => conv_std_logic_vector(25, 8),
24899 => conv_std_logic_vector(25, 8),
24900 => conv_std_logic_vector(25, 8),
24901 => conv_std_logic_vector(26, 8),
24902 => conv_std_logic_vector(26, 8),
24903 => conv_std_logic_vector(26, 8),
24904 => conv_std_logic_vector(27, 8),
24905 => conv_std_logic_vector(27, 8),
24906 => conv_std_logic_vector(28, 8),
24907 => conv_std_logic_vector(28, 8),
24908 => conv_std_logic_vector(28, 8),
24909 => conv_std_logic_vector(29, 8),
24910 => conv_std_logic_vector(29, 8),
24911 => conv_std_logic_vector(29, 8),
24912 => conv_std_logic_vector(30, 8),
24913 => conv_std_logic_vector(30, 8),
24914 => conv_std_logic_vector(31, 8),
24915 => conv_std_logic_vector(31, 8),
24916 => conv_std_logic_vector(31, 8),
24917 => conv_std_logic_vector(32, 8),
24918 => conv_std_logic_vector(32, 8),
24919 => conv_std_logic_vector(32, 8),
24920 => conv_std_logic_vector(33, 8),
24921 => conv_std_logic_vector(33, 8),
24922 => conv_std_logic_vector(34, 8),
24923 => conv_std_logic_vector(34, 8),
24924 => conv_std_logic_vector(34, 8),
24925 => conv_std_logic_vector(35, 8),
24926 => conv_std_logic_vector(35, 8),
24927 => conv_std_logic_vector(35, 8),
24928 => conv_std_logic_vector(36, 8),
24929 => conv_std_logic_vector(36, 8),
24930 => conv_std_logic_vector(37, 8),
24931 => conv_std_logic_vector(37, 8),
24932 => conv_std_logic_vector(37, 8),
24933 => conv_std_logic_vector(38, 8),
24934 => conv_std_logic_vector(38, 8),
24935 => conv_std_logic_vector(39, 8),
24936 => conv_std_logic_vector(39, 8),
24937 => conv_std_logic_vector(39, 8),
24938 => conv_std_logic_vector(40, 8),
24939 => conv_std_logic_vector(40, 8),
24940 => conv_std_logic_vector(40, 8),
24941 => conv_std_logic_vector(41, 8),
24942 => conv_std_logic_vector(41, 8),
24943 => conv_std_logic_vector(42, 8),
24944 => conv_std_logic_vector(42, 8),
24945 => conv_std_logic_vector(42, 8),
24946 => conv_std_logic_vector(43, 8),
24947 => conv_std_logic_vector(43, 8),
24948 => conv_std_logic_vector(43, 8),
24949 => conv_std_logic_vector(44, 8),
24950 => conv_std_logic_vector(44, 8),
24951 => conv_std_logic_vector(45, 8),
24952 => conv_std_logic_vector(45, 8),
24953 => conv_std_logic_vector(45, 8),
24954 => conv_std_logic_vector(46, 8),
24955 => conv_std_logic_vector(46, 8),
24956 => conv_std_logic_vector(46, 8),
24957 => conv_std_logic_vector(47, 8),
24958 => conv_std_logic_vector(47, 8),
24959 => conv_std_logic_vector(48, 8),
24960 => conv_std_logic_vector(48, 8),
24961 => conv_std_logic_vector(48, 8),
24962 => conv_std_logic_vector(49, 8),
24963 => conv_std_logic_vector(49, 8),
24964 => conv_std_logic_vector(50, 8),
24965 => conv_std_logic_vector(50, 8),
24966 => conv_std_logic_vector(50, 8),
24967 => conv_std_logic_vector(51, 8),
24968 => conv_std_logic_vector(51, 8),
24969 => conv_std_logic_vector(51, 8),
24970 => conv_std_logic_vector(52, 8),
24971 => conv_std_logic_vector(52, 8),
24972 => conv_std_logic_vector(53, 8),
24973 => conv_std_logic_vector(53, 8),
24974 => conv_std_logic_vector(53, 8),
24975 => conv_std_logic_vector(54, 8),
24976 => conv_std_logic_vector(54, 8),
24977 => conv_std_logic_vector(54, 8),
24978 => conv_std_logic_vector(55, 8),
24979 => conv_std_logic_vector(55, 8),
24980 => conv_std_logic_vector(56, 8),
24981 => conv_std_logic_vector(56, 8),
24982 => conv_std_logic_vector(56, 8),
24983 => conv_std_logic_vector(57, 8),
24984 => conv_std_logic_vector(57, 8),
24985 => conv_std_logic_vector(57, 8),
24986 => conv_std_logic_vector(58, 8),
24987 => conv_std_logic_vector(58, 8),
24988 => conv_std_logic_vector(59, 8),
24989 => conv_std_logic_vector(59, 8),
24990 => conv_std_logic_vector(59, 8),
24991 => conv_std_logic_vector(60, 8),
24992 => conv_std_logic_vector(60, 8),
24993 => conv_std_logic_vector(61, 8),
24994 => conv_std_logic_vector(61, 8),
24995 => conv_std_logic_vector(61, 8),
24996 => conv_std_logic_vector(62, 8),
24997 => conv_std_logic_vector(62, 8),
24998 => conv_std_logic_vector(62, 8),
24999 => conv_std_logic_vector(63, 8),
25000 => conv_std_logic_vector(63, 8),
25001 => conv_std_logic_vector(64, 8),
25002 => conv_std_logic_vector(64, 8),
25003 => conv_std_logic_vector(64, 8),
25004 => conv_std_logic_vector(65, 8),
25005 => conv_std_logic_vector(65, 8),
25006 => conv_std_logic_vector(65, 8),
25007 => conv_std_logic_vector(66, 8),
25008 => conv_std_logic_vector(66, 8),
25009 => conv_std_logic_vector(67, 8),
25010 => conv_std_logic_vector(67, 8),
25011 => conv_std_logic_vector(67, 8),
25012 => conv_std_logic_vector(68, 8),
25013 => conv_std_logic_vector(68, 8),
25014 => conv_std_logic_vector(68, 8),
25015 => conv_std_logic_vector(69, 8),
25016 => conv_std_logic_vector(69, 8),
25017 => conv_std_logic_vector(70, 8),
25018 => conv_std_logic_vector(70, 8),
25019 => conv_std_logic_vector(70, 8),
25020 => conv_std_logic_vector(71, 8),
25021 => conv_std_logic_vector(71, 8),
25022 => conv_std_logic_vector(71, 8),
25023 => conv_std_logic_vector(72, 8),
25024 => conv_std_logic_vector(72, 8),
25025 => conv_std_logic_vector(73, 8),
25026 => conv_std_logic_vector(73, 8),
25027 => conv_std_logic_vector(73, 8),
25028 => conv_std_logic_vector(74, 8),
25029 => conv_std_logic_vector(74, 8),
25030 => conv_std_logic_vector(75, 8),
25031 => conv_std_logic_vector(75, 8),
25032 => conv_std_logic_vector(75, 8),
25033 => conv_std_logic_vector(76, 8),
25034 => conv_std_logic_vector(76, 8),
25035 => conv_std_logic_vector(76, 8),
25036 => conv_std_logic_vector(77, 8),
25037 => conv_std_logic_vector(77, 8),
25038 => conv_std_logic_vector(78, 8),
25039 => conv_std_logic_vector(78, 8),
25040 => conv_std_logic_vector(78, 8),
25041 => conv_std_logic_vector(79, 8),
25042 => conv_std_logic_vector(79, 8),
25043 => conv_std_logic_vector(79, 8),
25044 => conv_std_logic_vector(80, 8),
25045 => conv_std_logic_vector(80, 8),
25046 => conv_std_logic_vector(81, 8),
25047 => conv_std_logic_vector(81, 8),
25048 => conv_std_logic_vector(81, 8),
25049 => conv_std_logic_vector(82, 8),
25050 => conv_std_logic_vector(82, 8),
25051 => conv_std_logic_vector(82, 8),
25052 => conv_std_logic_vector(83, 8),
25053 => conv_std_logic_vector(83, 8),
25054 => conv_std_logic_vector(84, 8),
25055 => conv_std_logic_vector(84, 8),
25056 => conv_std_logic_vector(84, 8),
25057 => conv_std_logic_vector(85, 8),
25058 => conv_std_logic_vector(85, 8),
25059 => conv_std_logic_vector(86, 8),
25060 => conv_std_logic_vector(86, 8),
25061 => conv_std_logic_vector(86, 8),
25062 => conv_std_logic_vector(87, 8),
25063 => conv_std_logic_vector(87, 8),
25064 => conv_std_logic_vector(87, 8),
25065 => conv_std_logic_vector(88, 8),
25066 => conv_std_logic_vector(88, 8),
25067 => conv_std_logic_vector(89, 8),
25068 => conv_std_logic_vector(89, 8),
25069 => conv_std_logic_vector(89, 8),
25070 => conv_std_logic_vector(90, 8),
25071 => conv_std_logic_vector(90, 8),
25072 => conv_std_logic_vector(90, 8),
25073 => conv_std_logic_vector(91, 8),
25074 => conv_std_logic_vector(91, 8),
25075 => conv_std_logic_vector(92, 8),
25076 => conv_std_logic_vector(92, 8),
25077 => conv_std_logic_vector(92, 8),
25078 => conv_std_logic_vector(93, 8),
25079 => conv_std_logic_vector(93, 8),
25080 => conv_std_logic_vector(93, 8),
25081 => conv_std_logic_vector(94, 8),
25082 => conv_std_logic_vector(94, 8),
25083 => conv_std_logic_vector(95, 8),
25084 => conv_std_logic_vector(95, 8),
25085 => conv_std_logic_vector(95, 8),
25086 => conv_std_logic_vector(96, 8),
25087 => conv_std_logic_vector(96, 8),
25088 => conv_std_logic_vector(0, 8),
25089 => conv_std_logic_vector(0, 8),
25090 => conv_std_logic_vector(0, 8),
25091 => conv_std_logic_vector(1, 8),
25092 => conv_std_logic_vector(1, 8),
25093 => conv_std_logic_vector(1, 8),
25094 => conv_std_logic_vector(2, 8),
25095 => conv_std_logic_vector(2, 8),
25096 => conv_std_logic_vector(3, 8),
25097 => conv_std_logic_vector(3, 8),
25098 => conv_std_logic_vector(3, 8),
25099 => conv_std_logic_vector(4, 8),
25100 => conv_std_logic_vector(4, 8),
25101 => conv_std_logic_vector(4, 8),
25102 => conv_std_logic_vector(5, 8),
25103 => conv_std_logic_vector(5, 8),
25104 => conv_std_logic_vector(6, 8),
25105 => conv_std_logic_vector(6, 8),
25106 => conv_std_logic_vector(6, 8),
25107 => conv_std_logic_vector(7, 8),
25108 => conv_std_logic_vector(7, 8),
25109 => conv_std_logic_vector(8, 8),
25110 => conv_std_logic_vector(8, 8),
25111 => conv_std_logic_vector(8, 8),
25112 => conv_std_logic_vector(9, 8),
25113 => conv_std_logic_vector(9, 8),
25114 => conv_std_logic_vector(9, 8),
25115 => conv_std_logic_vector(10, 8),
25116 => conv_std_logic_vector(10, 8),
25117 => conv_std_logic_vector(11, 8),
25118 => conv_std_logic_vector(11, 8),
25119 => conv_std_logic_vector(11, 8),
25120 => conv_std_logic_vector(12, 8),
25121 => conv_std_logic_vector(12, 8),
25122 => conv_std_logic_vector(13, 8),
25123 => conv_std_logic_vector(13, 8),
25124 => conv_std_logic_vector(13, 8),
25125 => conv_std_logic_vector(14, 8),
25126 => conv_std_logic_vector(14, 8),
25127 => conv_std_logic_vector(14, 8),
25128 => conv_std_logic_vector(15, 8),
25129 => conv_std_logic_vector(15, 8),
25130 => conv_std_logic_vector(16, 8),
25131 => conv_std_logic_vector(16, 8),
25132 => conv_std_logic_vector(16, 8),
25133 => conv_std_logic_vector(17, 8),
25134 => conv_std_logic_vector(17, 8),
25135 => conv_std_logic_vector(17, 8),
25136 => conv_std_logic_vector(18, 8),
25137 => conv_std_logic_vector(18, 8),
25138 => conv_std_logic_vector(19, 8),
25139 => conv_std_logic_vector(19, 8),
25140 => conv_std_logic_vector(19, 8),
25141 => conv_std_logic_vector(20, 8),
25142 => conv_std_logic_vector(20, 8),
25143 => conv_std_logic_vector(21, 8),
25144 => conv_std_logic_vector(21, 8),
25145 => conv_std_logic_vector(21, 8),
25146 => conv_std_logic_vector(22, 8),
25147 => conv_std_logic_vector(22, 8),
25148 => conv_std_logic_vector(22, 8),
25149 => conv_std_logic_vector(23, 8),
25150 => conv_std_logic_vector(23, 8),
25151 => conv_std_logic_vector(24, 8),
25152 => conv_std_logic_vector(24, 8),
25153 => conv_std_logic_vector(24, 8),
25154 => conv_std_logic_vector(25, 8),
25155 => conv_std_logic_vector(25, 8),
25156 => conv_std_logic_vector(26, 8),
25157 => conv_std_logic_vector(26, 8),
25158 => conv_std_logic_vector(26, 8),
25159 => conv_std_logic_vector(27, 8),
25160 => conv_std_logic_vector(27, 8),
25161 => conv_std_logic_vector(27, 8),
25162 => conv_std_logic_vector(28, 8),
25163 => conv_std_logic_vector(28, 8),
25164 => conv_std_logic_vector(29, 8),
25165 => conv_std_logic_vector(29, 8),
25166 => conv_std_logic_vector(29, 8),
25167 => conv_std_logic_vector(30, 8),
25168 => conv_std_logic_vector(30, 8),
25169 => conv_std_logic_vector(31, 8),
25170 => conv_std_logic_vector(31, 8),
25171 => conv_std_logic_vector(31, 8),
25172 => conv_std_logic_vector(32, 8),
25173 => conv_std_logic_vector(32, 8),
25174 => conv_std_logic_vector(32, 8),
25175 => conv_std_logic_vector(33, 8),
25176 => conv_std_logic_vector(33, 8),
25177 => conv_std_logic_vector(34, 8),
25178 => conv_std_logic_vector(34, 8),
25179 => conv_std_logic_vector(34, 8),
25180 => conv_std_logic_vector(35, 8),
25181 => conv_std_logic_vector(35, 8),
25182 => conv_std_logic_vector(35, 8),
25183 => conv_std_logic_vector(36, 8),
25184 => conv_std_logic_vector(36, 8),
25185 => conv_std_logic_vector(37, 8),
25186 => conv_std_logic_vector(37, 8),
25187 => conv_std_logic_vector(37, 8),
25188 => conv_std_logic_vector(38, 8),
25189 => conv_std_logic_vector(38, 8),
25190 => conv_std_logic_vector(39, 8),
25191 => conv_std_logic_vector(39, 8),
25192 => conv_std_logic_vector(39, 8),
25193 => conv_std_logic_vector(40, 8),
25194 => conv_std_logic_vector(40, 8),
25195 => conv_std_logic_vector(40, 8),
25196 => conv_std_logic_vector(41, 8),
25197 => conv_std_logic_vector(41, 8),
25198 => conv_std_logic_vector(42, 8),
25199 => conv_std_logic_vector(42, 8),
25200 => conv_std_logic_vector(42, 8),
25201 => conv_std_logic_vector(43, 8),
25202 => conv_std_logic_vector(43, 8),
25203 => conv_std_logic_vector(44, 8),
25204 => conv_std_logic_vector(44, 8),
25205 => conv_std_logic_vector(44, 8),
25206 => conv_std_logic_vector(45, 8),
25207 => conv_std_logic_vector(45, 8),
25208 => conv_std_logic_vector(45, 8),
25209 => conv_std_logic_vector(46, 8),
25210 => conv_std_logic_vector(46, 8),
25211 => conv_std_logic_vector(47, 8),
25212 => conv_std_logic_vector(47, 8),
25213 => conv_std_logic_vector(47, 8),
25214 => conv_std_logic_vector(48, 8),
25215 => conv_std_logic_vector(48, 8),
25216 => conv_std_logic_vector(49, 8),
25217 => conv_std_logic_vector(49, 8),
25218 => conv_std_logic_vector(49, 8),
25219 => conv_std_logic_vector(50, 8),
25220 => conv_std_logic_vector(50, 8),
25221 => conv_std_logic_vector(50, 8),
25222 => conv_std_logic_vector(51, 8),
25223 => conv_std_logic_vector(51, 8),
25224 => conv_std_logic_vector(52, 8),
25225 => conv_std_logic_vector(52, 8),
25226 => conv_std_logic_vector(52, 8),
25227 => conv_std_logic_vector(53, 8),
25228 => conv_std_logic_vector(53, 8),
25229 => conv_std_logic_vector(53, 8),
25230 => conv_std_logic_vector(54, 8),
25231 => conv_std_logic_vector(54, 8),
25232 => conv_std_logic_vector(55, 8),
25233 => conv_std_logic_vector(55, 8),
25234 => conv_std_logic_vector(55, 8),
25235 => conv_std_logic_vector(56, 8),
25236 => conv_std_logic_vector(56, 8),
25237 => conv_std_logic_vector(57, 8),
25238 => conv_std_logic_vector(57, 8),
25239 => conv_std_logic_vector(57, 8),
25240 => conv_std_logic_vector(58, 8),
25241 => conv_std_logic_vector(58, 8),
25242 => conv_std_logic_vector(58, 8),
25243 => conv_std_logic_vector(59, 8),
25244 => conv_std_logic_vector(59, 8),
25245 => conv_std_logic_vector(60, 8),
25246 => conv_std_logic_vector(60, 8),
25247 => conv_std_logic_vector(60, 8),
25248 => conv_std_logic_vector(61, 8),
25249 => conv_std_logic_vector(61, 8),
25250 => conv_std_logic_vector(62, 8),
25251 => conv_std_logic_vector(62, 8),
25252 => conv_std_logic_vector(62, 8),
25253 => conv_std_logic_vector(63, 8),
25254 => conv_std_logic_vector(63, 8),
25255 => conv_std_logic_vector(63, 8),
25256 => conv_std_logic_vector(64, 8),
25257 => conv_std_logic_vector(64, 8),
25258 => conv_std_logic_vector(65, 8),
25259 => conv_std_logic_vector(65, 8),
25260 => conv_std_logic_vector(65, 8),
25261 => conv_std_logic_vector(66, 8),
25262 => conv_std_logic_vector(66, 8),
25263 => conv_std_logic_vector(66, 8),
25264 => conv_std_logic_vector(67, 8),
25265 => conv_std_logic_vector(67, 8),
25266 => conv_std_logic_vector(68, 8),
25267 => conv_std_logic_vector(68, 8),
25268 => conv_std_logic_vector(68, 8),
25269 => conv_std_logic_vector(69, 8),
25270 => conv_std_logic_vector(69, 8),
25271 => conv_std_logic_vector(70, 8),
25272 => conv_std_logic_vector(70, 8),
25273 => conv_std_logic_vector(70, 8),
25274 => conv_std_logic_vector(71, 8),
25275 => conv_std_logic_vector(71, 8),
25276 => conv_std_logic_vector(71, 8),
25277 => conv_std_logic_vector(72, 8),
25278 => conv_std_logic_vector(72, 8),
25279 => conv_std_logic_vector(73, 8),
25280 => conv_std_logic_vector(73, 8),
25281 => conv_std_logic_vector(73, 8),
25282 => conv_std_logic_vector(74, 8),
25283 => conv_std_logic_vector(74, 8),
25284 => conv_std_logic_vector(75, 8),
25285 => conv_std_logic_vector(75, 8),
25286 => conv_std_logic_vector(75, 8),
25287 => conv_std_logic_vector(76, 8),
25288 => conv_std_logic_vector(76, 8),
25289 => conv_std_logic_vector(76, 8),
25290 => conv_std_logic_vector(77, 8),
25291 => conv_std_logic_vector(77, 8),
25292 => conv_std_logic_vector(78, 8),
25293 => conv_std_logic_vector(78, 8),
25294 => conv_std_logic_vector(78, 8),
25295 => conv_std_logic_vector(79, 8),
25296 => conv_std_logic_vector(79, 8),
25297 => conv_std_logic_vector(80, 8),
25298 => conv_std_logic_vector(80, 8),
25299 => conv_std_logic_vector(80, 8),
25300 => conv_std_logic_vector(81, 8),
25301 => conv_std_logic_vector(81, 8),
25302 => conv_std_logic_vector(81, 8),
25303 => conv_std_logic_vector(82, 8),
25304 => conv_std_logic_vector(82, 8),
25305 => conv_std_logic_vector(83, 8),
25306 => conv_std_logic_vector(83, 8),
25307 => conv_std_logic_vector(83, 8),
25308 => conv_std_logic_vector(84, 8),
25309 => conv_std_logic_vector(84, 8),
25310 => conv_std_logic_vector(84, 8),
25311 => conv_std_logic_vector(85, 8),
25312 => conv_std_logic_vector(85, 8),
25313 => conv_std_logic_vector(86, 8),
25314 => conv_std_logic_vector(86, 8),
25315 => conv_std_logic_vector(86, 8),
25316 => conv_std_logic_vector(87, 8),
25317 => conv_std_logic_vector(87, 8),
25318 => conv_std_logic_vector(88, 8),
25319 => conv_std_logic_vector(88, 8),
25320 => conv_std_logic_vector(88, 8),
25321 => conv_std_logic_vector(89, 8),
25322 => conv_std_logic_vector(89, 8),
25323 => conv_std_logic_vector(89, 8),
25324 => conv_std_logic_vector(90, 8),
25325 => conv_std_logic_vector(90, 8),
25326 => conv_std_logic_vector(91, 8),
25327 => conv_std_logic_vector(91, 8),
25328 => conv_std_logic_vector(91, 8),
25329 => conv_std_logic_vector(92, 8),
25330 => conv_std_logic_vector(92, 8),
25331 => conv_std_logic_vector(93, 8),
25332 => conv_std_logic_vector(93, 8),
25333 => conv_std_logic_vector(93, 8),
25334 => conv_std_logic_vector(94, 8),
25335 => conv_std_logic_vector(94, 8),
25336 => conv_std_logic_vector(94, 8),
25337 => conv_std_logic_vector(95, 8),
25338 => conv_std_logic_vector(95, 8),
25339 => conv_std_logic_vector(96, 8),
25340 => conv_std_logic_vector(96, 8),
25341 => conv_std_logic_vector(96, 8),
25342 => conv_std_logic_vector(97, 8),
25343 => conv_std_logic_vector(97, 8),
25344 => conv_std_logic_vector(0, 8),
25345 => conv_std_logic_vector(0, 8),
25346 => conv_std_logic_vector(0, 8),
25347 => conv_std_logic_vector(1, 8),
25348 => conv_std_logic_vector(1, 8),
25349 => conv_std_logic_vector(1, 8),
25350 => conv_std_logic_vector(2, 8),
25351 => conv_std_logic_vector(2, 8),
25352 => conv_std_logic_vector(3, 8),
25353 => conv_std_logic_vector(3, 8),
25354 => conv_std_logic_vector(3, 8),
25355 => conv_std_logic_vector(4, 8),
25356 => conv_std_logic_vector(4, 8),
25357 => conv_std_logic_vector(5, 8),
25358 => conv_std_logic_vector(5, 8),
25359 => conv_std_logic_vector(5, 8),
25360 => conv_std_logic_vector(6, 8),
25361 => conv_std_logic_vector(6, 8),
25362 => conv_std_logic_vector(6, 8),
25363 => conv_std_logic_vector(7, 8),
25364 => conv_std_logic_vector(7, 8),
25365 => conv_std_logic_vector(8, 8),
25366 => conv_std_logic_vector(8, 8),
25367 => conv_std_logic_vector(8, 8),
25368 => conv_std_logic_vector(9, 8),
25369 => conv_std_logic_vector(9, 8),
25370 => conv_std_logic_vector(10, 8),
25371 => conv_std_logic_vector(10, 8),
25372 => conv_std_logic_vector(10, 8),
25373 => conv_std_logic_vector(11, 8),
25374 => conv_std_logic_vector(11, 8),
25375 => conv_std_logic_vector(11, 8),
25376 => conv_std_logic_vector(12, 8),
25377 => conv_std_logic_vector(12, 8),
25378 => conv_std_logic_vector(13, 8),
25379 => conv_std_logic_vector(13, 8),
25380 => conv_std_logic_vector(13, 8),
25381 => conv_std_logic_vector(14, 8),
25382 => conv_std_logic_vector(14, 8),
25383 => conv_std_logic_vector(15, 8),
25384 => conv_std_logic_vector(15, 8),
25385 => conv_std_logic_vector(15, 8),
25386 => conv_std_logic_vector(16, 8),
25387 => conv_std_logic_vector(16, 8),
25388 => conv_std_logic_vector(17, 8),
25389 => conv_std_logic_vector(17, 8),
25390 => conv_std_logic_vector(17, 8),
25391 => conv_std_logic_vector(18, 8),
25392 => conv_std_logic_vector(18, 8),
25393 => conv_std_logic_vector(18, 8),
25394 => conv_std_logic_vector(19, 8),
25395 => conv_std_logic_vector(19, 8),
25396 => conv_std_logic_vector(20, 8),
25397 => conv_std_logic_vector(20, 8),
25398 => conv_std_logic_vector(20, 8),
25399 => conv_std_logic_vector(21, 8),
25400 => conv_std_logic_vector(21, 8),
25401 => conv_std_logic_vector(22, 8),
25402 => conv_std_logic_vector(22, 8),
25403 => conv_std_logic_vector(22, 8),
25404 => conv_std_logic_vector(23, 8),
25405 => conv_std_logic_vector(23, 8),
25406 => conv_std_logic_vector(23, 8),
25407 => conv_std_logic_vector(24, 8),
25408 => conv_std_logic_vector(24, 8),
25409 => conv_std_logic_vector(25, 8),
25410 => conv_std_logic_vector(25, 8),
25411 => conv_std_logic_vector(25, 8),
25412 => conv_std_logic_vector(26, 8),
25413 => conv_std_logic_vector(26, 8),
25414 => conv_std_logic_vector(27, 8),
25415 => conv_std_logic_vector(27, 8),
25416 => conv_std_logic_vector(27, 8),
25417 => conv_std_logic_vector(28, 8),
25418 => conv_std_logic_vector(28, 8),
25419 => conv_std_logic_vector(29, 8),
25420 => conv_std_logic_vector(29, 8),
25421 => conv_std_logic_vector(29, 8),
25422 => conv_std_logic_vector(30, 8),
25423 => conv_std_logic_vector(30, 8),
25424 => conv_std_logic_vector(30, 8),
25425 => conv_std_logic_vector(31, 8),
25426 => conv_std_logic_vector(31, 8),
25427 => conv_std_logic_vector(32, 8),
25428 => conv_std_logic_vector(32, 8),
25429 => conv_std_logic_vector(32, 8),
25430 => conv_std_logic_vector(33, 8),
25431 => conv_std_logic_vector(33, 8),
25432 => conv_std_logic_vector(34, 8),
25433 => conv_std_logic_vector(34, 8),
25434 => conv_std_logic_vector(34, 8),
25435 => conv_std_logic_vector(35, 8),
25436 => conv_std_logic_vector(35, 8),
25437 => conv_std_logic_vector(35, 8),
25438 => conv_std_logic_vector(36, 8),
25439 => conv_std_logic_vector(36, 8),
25440 => conv_std_logic_vector(37, 8),
25441 => conv_std_logic_vector(37, 8),
25442 => conv_std_logic_vector(37, 8),
25443 => conv_std_logic_vector(38, 8),
25444 => conv_std_logic_vector(38, 8),
25445 => conv_std_logic_vector(39, 8),
25446 => conv_std_logic_vector(39, 8),
25447 => conv_std_logic_vector(39, 8),
25448 => conv_std_logic_vector(40, 8),
25449 => conv_std_logic_vector(40, 8),
25450 => conv_std_logic_vector(40, 8),
25451 => conv_std_logic_vector(41, 8),
25452 => conv_std_logic_vector(41, 8),
25453 => conv_std_logic_vector(42, 8),
25454 => conv_std_logic_vector(42, 8),
25455 => conv_std_logic_vector(42, 8),
25456 => conv_std_logic_vector(43, 8),
25457 => conv_std_logic_vector(43, 8),
25458 => conv_std_logic_vector(44, 8),
25459 => conv_std_logic_vector(44, 8),
25460 => conv_std_logic_vector(44, 8),
25461 => conv_std_logic_vector(45, 8),
25462 => conv_std_logic_vector(45, 8),
25463 => conv_std_logic_vector(46, 8),
25464 => conv_std_logic_vector(46, 8),
25465 => conv_std_logic_vector(46, 8),
25466 => conv_std_logic_vector(47, 8),
25467 => conv_std_logic_vector(47, 8),
25468 => conv_std_logic_vector(47, 8),
25469 => conv_std_logic_vector(48, 8),
25470 => conv_std_logic_vector(48, 8),
25471 => conv_std_logic_vector(49, 8),
25472 => conv_std_logic_vector(49, 8),
25473 => conv_std_logic_vector(49, 8),
25474 => conv_std_logic_vector(50, 8),
25475 => conv_std_logic_vector(50, 8),
25476 => conv_std_logic_vector(51, 8),
25477 => conv_std_logic_vector(51, 8),
25478 => conv_std_logic_vector(51, 8),
25479 => conv_std_logic_vector(52, 8),
25480 => conv_std_logic_vector(52, 8),
25481 => conv_std_logic_vector(52, 8),
25482 => conv_std_logic_vector(53, 8),
25483 => conv_std_logic_vector(53, 8),
25484 => conv_std_logic_vector(54, 8),
25485 => conv_std_logic_vector(54, 8),
25486 => conv_std_logic_vector(54, 8),
25487 => conv_std_logic_vector(55, 8),
25488 => conv_std_logic_vector(55, 8),
25489 => conv_std_logic_vector(56, 8),
25490 => conv_std_logic_vector(56, 8),
25491 => conv_std_logic_vector(56, 8),
25492 => conv_std_logic_vector(57, 8),
25493 => conv_std_logic_vector(57, 8),
25494 => conv_std_logic_vector(58, 8),
25495 => conv_std_logic_vector(58, 8),
25496 => conv_std_logic_vector(58, 8),
25497 => conv_std_logic_vector(59, 8),
25498 => conv_std_logic_vector(59, 8),
25499 => conv_std_logic_vector(59, 8),
25500 => conv_std_logic_vector(60, 8),
25501 => conv_std_logic_vector(60, 8),
25502 => conv_std_logic_vector(61, 8),
25503 => conv_std_logic_vector(61, 8),
25504 => conv_std_logic_vector(61, 8),
25505 => conv_std_logic_vector(62, 8),
25506 => conv_std_logic_vector(62, 8),
25507 => conv_std_logic_vector(63, 8),
25508 => conv_std_logic_vector(63, 8),
25509 => conv_std_logic_vector(63, 8),
25510 => conv_std_logic_vector(64, 8),
25511 => conv_std_logic_vector(64, 8),
25512 => conv_std_logic_vector(64, 8),
25513 => conv_std_logic_vector(65, 8),
25514 => conv_std_logic_vector(65, 8),
25515 => conv_std_logic_vector(66, 8),
25516 => conv_std_logic_vector(66, 8),
25517 => conv_std_logic_vector(66, 8),
25518 => conv_std_logic_vector(67, 8),
25519 => conv_std_logic_vector(67, 8),
25520 => conv_std_logic_vector(68, 8),
25521 => conv_std_logic_vector(68, 8),
25522 => conv_std_logic_vector(68, 8),
25523 => conv_std_logic_vector(69, 8),
25524 => conv_std_logic_vector(69, 8),
25525 => conv_std_logic_vector(69, 8),
25526 => conv_std_logic_vector(70, 8),
25527 => conv_std_logic_vector(70, 8),
25528 => conv_std_logic_vector(71, 8),
25529 => conv_std_logic_vector(71, 8),
25530 => conv_std_logic_vector(71, 8),
25531 => conv_std_logic_vector(72, 8),
25532 => conv_std_logic_vector(72, 8),
25533 => conv_std_logic_vector(73, 8),
25534 => conv_std_logic_vector(73, 8),
25535 => conv_std_logic_vector(73, 8),
25536 => conv_std_logic_vector(74, 8),
25537 => conv_std_logic_vector(74, 8),
25538 => conv_std_logic_vector(75, 8),
25539 => conv_std_logic_vector(75, 8),
25540 => conv_std_logic_vector(75, 8),
25541 => conv_std_logic_vector(76, 8),
25542 => conv_std_logic_vector(76, 8),
25543 => conv_std_logic_vector(76, 8),
25544 => conv_std_logic_vector(77, 8),
25545 => conv_std_logic_vector(77, 8),
25546 => conv_std_logic_vector(78, 8),
25547 => conv_std_logic_vector(78, 8),
25548 => conv_std_logic_vector(78, 8),
25549 => conv_std_logic_vector(79, 8),
25550 => conv_std_logic_vector(79, 8),
25551 => conv_std_logic_vector(80, 8),
25552 => conv_std_logic_vector(80, 8),
25553 => conv_std_logic_vector(80, 8),
25554 => conv_std_logic_vector(81, 8),
25555 => conv_std_logic_vector(81, 8),
25556 => conv_std_logic_vector(81, 8),
25557 => conv_std_logic_vector(82, 8),
25558 => conv_std_logic_vector(82, 8),
25559 => conv_std_logic_vector(83, 8),
25560 => conv_std_logic_vector(83, 8),
25561 => conv_std_logic_vector(83, 8),
25562 => conv_std_logic_vector(84, 8),
25563 => conv_std_logic_vector(84, 8),
25564 => conv_std_logic_vector(85, 8),
25565 => conv_std_logic_vector(85, 8),
25566 => conv_std_logic_vector(85, 8),
25567 => conv_std_logic_vector(86, 8),
25568 => conv_std_logic_vector(86, 8),
25569 => conv_std_logic_vector(87, 8),
25570 => conv_std_logic_vector(87, 8),
25571 => conv_std_logic_vector(87, 8),
25572 => conv_std_logic_vector(88, 8),
25573 => conv_std_logic_vector(88, 8),
25574 => conv_std_logic_vector(88, 8),
25575 => conv_std_logic_vector(89, 8),
25576 => conv_std_logic_vector(89, 8),
25577 => conv_std_logic_vector(90, 8),
25578 => conv_std_logic_vector(90, 8),
25579 => conv_std_logic_vector(90, 8),
25580 => conv_std_logic_vector(91, 8),
25581 => conv_std_logic_vector(91, 8),
25582 => conv_std_logic_vector(92, 8),
25583 => conv_std_logic_vector(92, 8),
25584 => conv_std_logic_vector(92, 8),
25585 => conv_std_logic_vector(93, 8),
25586 => conv_std_logic_vector(93, 8),
25587 => conv_std_logic_vector(93, 8),
25588 => conv_std_logic_vector(94, 8),
25589 => conv_std_logic_vector(94, 8),
25590 => conv_std_logic_vector(95, 8),
25591 => conv_std_logic_vector(95, 8),
25592 => conv_std_logic_vector(95, 8),
25593 => conv_std_logic_vector(96, 8),
25594 => conv_std_logic_vector(96, 8),
25595 => conv_std_logic_vector(97, 8),
25596 => conv_std_logic_vector(97, 8),
25597 => conv_std_logic_vector(97, 8),
25598 => conv_std_logic_vector(98, 8),
25599 => conv_std_logic_vector(98, 8),
25600 => conv_std_logic_vector(0, 8),
25601 => conv_std_logic_vector(0, 8),
25602 => conv_std_logic_vector(0, 8),
25603 => conv_std_logic_vector(1, 8),
25604 => conv_std_logic_vector(1, 8),
25605 => conv_std_logic_vector(1, 8),
25606 => conv_std_logic_vector(2, 8),
25607 => conv_std_logic_vector(2, 8),
25608 => conv_std_logic_vector(3, 8),
25609 => conv_std_logic_vector(3, 8),
25610 => conv_std_logic_vector(3, 8),
25611 => conv_std_logic_vector(4, 8),
25612 => conv_std_logic_vector(4, 8),
25613 => conv_std_logic_vector(5, 8),
25614 => conv_std_logic_vector(5, 8),
25615 => conv_std_logic_vector(5, 8),
25616 => conv_std_logic_vector(6, 8),
25617 => conv_std_logic_vector(6, 8),
25618 => conv_std_logic_vector(7, 8),
25619 => conv_std_logic_vector(7, 8),
25620 => conv_std_logic_vector(7, 8),
25621 => conv_std_logic_vector(8, 8),
25622 => conv_std_logic_vector(8, 8),
25623 => conv_std_logic_vector(8, 8),
25624 => conv_std_logic_vector(9, 8),
25625 => conv_std_logic_vector(9, 8),
25626 => conv_std_logic_vector(10, 8),
25627 => conv_std_logic_vector(10, 8),
25628 => conv_std_logic_vector(10, 8),
25629 => conv_std_logic_vector(11, 8),
25630 => conv_std_logic_vector(11, 8),
25631 => conv_std_logic_vector(12, 8),
25632 => conv_std_logic_vector(12, 8),
25633 => conv_std_logic_vector(12, 8),
25634 => conv_std_logic_vector(13, 8),
25635 => conv_std_logic_vector(13, 8),
25636 => conv_std_logic_vector(14, 8),
25637 => conv_std_logic_vector(14, 8),
25638 => conv_std_logic_vector(14, 8),
25639 => conv_std_logic_vector(15, 8),
25640 => conv_std_logic_vector(15, 8),
25641 => conv_std_logic_vector(16, 8),
25642 => conv_std_logic_vector(16, 8),
25643 => conv_std_logic_vector(16, 8),
25644 => conv_std_logic_vector(17, 8),
25645 => conv_std_logic_vector(17, 8),
25646 => conv_std_logic_vector(17, 8),
25647 => conv_std_logic_vector(18, 8),
25648 => conv_std_logic_vector(18, 8),
25649 => conv_std_logic_vector(19, 8),
25650 => conv_std_logic_vector(19, 8),
25651 => conv_std_logic_vector(19, 8),
25652 => conv_std_logic_vector(20, 8),
25653 => conv_std_logic_vector(20, 8),
25654 => conv_std_logic_vector(21, 8),
25655 => conv_std_logic_vector(21, 8),
25656 => conv_std_logic_vector(21, 8),
25657 => conv_std_logic_vector(22, 8),
25658 => conv_std_logic_vector(22, 8),
25659 => conv_std_logic_vector(23, 8),
25660 => conv_std_logic_vector(23, 8),
25661 => conv_std_logic_vector(23, 8),
25662 => conv_std_logic_vector(24, 8),
25663 => conv_std_logic_vector(24, 8),
25664 => conv_std_logic_vector(25, 8),
25665 => conv_std_logic_vector(25, 8),
25666 => conv_std_logic_vector(25, 8),
25667 => conv_std_logic_vector(26, 8),
25668 => conv_std_logic_vector(26, 8),
25669 => conv_std_logic_vector(26, 8),
25670 => conv_std_logic_vector(27, 8),
25671 => conv_std_logic_vector(27, 8),
25672 => conv_std_logic_vector(28, 8),
25673 => conv_std_logic_vector(28, 8),
25674 => conv_std_logic_vector(28, 8),
25675 => conv_std_logic_vector(29, 8),
25676 => conv_std_logic_vector(29, 8),
25677 => conv_std_logic_vector(30, 8),
25678 => conv_std_logic_vector(30, 8),
25679 => conv_std_logic_vector(30, 8),
25680 => conv_std_logic_vector(31, 8),
25681 => conv_std_logic_vector(31, 8),
25682 => conv_std_logic_vector(32, 8),
25683 => conv_std_logic_vector(32, 8),
25684 => conv_std_logic_vector(32, 8),
25685 => conv_std_logic_vector(33, 8),
25686 => conv_std_logic_vector(33, 8),
25687 => conv_std_logic_vector(33, 8),
25688 => conv_std_logic_vector(34, 8),
25689 => conv_std_logic_vector(34, 8),
25690 => conv_std_logic_vector(35, 8),
25691 => conv_std_logic_vector(35, 8),
25692 => conv_std_logic_vector(35, 8),
25693 => conv_std_logic_vector(36, 8),
25694 => conv_std_logic_vector(36, 8),
25695 => conv_std_logic_vector(37, 8),
25696 => conv_std_logic_vector(37, 8),
25697 => conv_std_logic_vector(37, 8),
25698 => conv_std_logic_vector(38, 8),
25699 => conv_std_logic_vector(38, 8),
25700 => conv_std_logic_vector(39, 8),
25701 => conv_std_logic_vector(39, 8),
25702 => conv_std_logic_vector(39, 8),
25703 => conv_std_logic_vector(40, 8),
25704 => conv_std_logic_vector(40, 8),
25705 => conv_std_logic_vector(41, 8),
25706 => conv_std_logic_vector(41, 8),
25707 => conv_std_logic_vector(41, 8),
25708 => conv_std_logic_vector(42, 8),
25709 => conv_std_logic_vector(42, 8),
25710 => conv_std_logic_vector(42, 8),
25711 => conv_std_logic_vector(43, 8),
25712 => conv_std_logic_vector(43, 8),
25713 => conv_std_logic_vector(44, 8),
25714 => conv_std_logic_vector(44, 8),
25715 => conv_std_logic_vector(44, 8),
25716 => conv_std_logic_vector(45, 8),
25717 => conv_std_logic_vector(45, 8),
25718 => conv_std_logic_vector(46, 8),
25719 => conv_std_logic_vector(46, 8),
25720 => conv_std_logic_vector(46, 8),
25721 => conv_std_logic_vector(47, 8),
25722 => conv_std_logic_vector(47, 8),
25723 => conv_std_logic_vector(48, 8),
25724 => conv_std_logic_vector(48, 8),
25725 => conv_std_logic_vector(48, 8),
25726 => conv_std_logic_vector(49, 8),
25727 => conv_std_logic_vector(49, 8),
25728 => conv_std_logic_vector(50, 8),
25729 => conv_std_logic_vector(50, 8),
25730 => conv_std_logic_vector(50, 8),
25731 => conv_std_logic_vector(51, 8),
25732 => conv_std_logic_vector(51, 8),
25733 => conv_std_logic_vector(51, 8),
25734 => conv_std_logic_vector(52, 8),
25735 => conv_std_logic_vector(52, 8),
25736 => conv_std_logic_vector(53, 8),
25737 => conv_std_logic_vector(53, 8),
25738 => conv_std_logic_vector(53, 8),
25739 => conv_std_logic_vector(54, 8),
25740 => conv_std_logic_vector(54, 8),
25741 => conv_std_logic_vector(55, 8),
25742 => conv_std_logic_vector(55, 8),
25743 => conv_std_logic_vector(55, 8),
25744 => conv_std_logic_vector(56, 8),
25745 => conv_std_logic_vector(56, 8),
25746 => conv_std_logic_vector(57, 8),
25747 => conv_std_logic_vector(57, 8),
25748 => conv_std_logic_vector(57, 8),
25749 => conv_std_logic_vector(58, 8),
25750 => conv_std_logic_vector(58, 8),
25751 => conv_std_logic_vector(58, 8),
25752 => conv_std_logic_vector(59, 8),
25753 => conv_std_logic_vector(59, 8),
25754 => conv_std_logic_vector(60, 8),
25755 => conv_std_logic_vector(60, 8),
25756 => conv_std_logic_vector(60, 8),
25757 => conv_std_logic_vector(61, 8),
25758 => conv_std_logic_vector(61, 8),
25759 => conv_std_logic_vector(62, 8),
25760 => conv_std_logic_vector(62, 8),
25761 => conv_std_logic_vector(62, 8),
25762 => conv_std_logic_vector(63, 8),
25763 => conv_std_logic_vector(63, 8),
25764 => conv_std_logic_vector(64, 8),
25765 => conv_std_logic_vector(64, 8),
25766 => conv_std_logic_vector(64, 8),
25767 => conv_std_logic_vector(65, 8),
25768 => conv_std_logic_vector(65, 8),
25769 => conv_std_logic_vector(66, 8),
25770 => conv_std_logic_vector(66, 8),
25771 => conv_std_logic_vector(66, 8),
25772 => conv_std_logic_vector(67, 8),
25773 => conv_std_logic_vector(67, 8),
25774 => conv_std_logic_vector(67, 8),
25775 => conv_std_logic_vector(68, 8),
25776 => conv_std_logic_vector(68, 8),
25777 => conv_std_logic_vector(69, 8),
25778 => conv_std_logic_vector(69, 8),
25779 => conv_std_logic_vector(69, 8),
25780 => conv_std_logic_vector(70, 8),
25781 => conv_std_logic_vector(70, 8),
25782 => conv_std_logic_vector(71, 8),
25783 => conv_std_logic_vector(71, 8),
25784 => conv_std_logic_vector(71, 8),
25785 => conv_std_logic_vector(72, 8),
25786 => conv_std_logic_vector(72, 8),
25787 => conv_std_logic_vector(73, 8),
25788 => conv_std_logic_vector(73, 8),
25789 => conv_std_logic_vector(73, 8),
25790 => conv_std_logic_vector(74, 8),
25791 => conv_std_logic_vector(74, 8),
25792 => conv_std_logic_vector(75, 8),
25793 => conv_std_logic_vector(75, 8),
25794 => conv_std_logic_vector(75, 8),
25795 => conv_std_logic_vector(76, 8),
25796 => conv_std_logic_vector(76, 8),
25797 => conv_std_logic_vector(76, 8),
25798 => conv_std_logic_vector(77, 8),
25799 => conv_std_logic_vector(77, 8),
25800 => conv_std_logic_vector(78, 8),
25801 => conv_std_logic_vector(78, 8),
25802 => conv_std_logic_vector(78, 8),
25803 => conv_std_logic_vector(79, 8),
25804 => conv_std_logic_vector(79, 8),
25805 => conv_std_logic_vector(80, 8),
25806 => conv_std_logic_vector(80, 8),
25807 => conv_std_logic_vector(80, 8),
25808 => conv_std_logic_vector(81, 8),
25809 => conv_std_logic_vector(81, 8),
25810 => conv_std_logic_vector(82, 8),
25811 => conv_std_logic_vector(82, 8),
25812 => conv_std_logic_vector(82, 8),
25813 => conv_std_logic_vector(83, 8),
25814 => conv_std_logic_vector(83, 8),
25815 => conv_std_logic_vector(83, 8),
25816 => conv_std_logic_vector(84, 8),
25817 => conv_std_logic_vector(84, 8),
25818 => conv_std_logic_vector(85, 8),
25819 => conv_std_logic_vector(85, 8),
25820 => conv_std_logic_vector(85, 8),
25821 => conv_std_logic_vector(86, 8),
25822 => conv_std_logic_vector(86, 8),
25823 => conv_std_logic_vector(87, 8),
25824 => conv_std_logic_vector(87, 8),
25825 => conv_std_logic_vector(87, 8),
25826 => conv_std_logic_vector(88, 8),
25827 => conv_std_logic_vector(88, 8),
25828 => conv_std_logic_vector(89, 8),
25829 => conv_std_logic_vector(89, 8),
25830 => conv_std_logic_vector(89, 8),
25831 => conv_std_logic_vector(90, 8),
25832 => conv_std_logic_vector(90, 8),
25833 => conv_std_logic_vector(91, 8),
25834 => conv_std_logic_vector(91, 8),
25835 => conv_std_logic_vector(91, 8),
25836 => conv_std_logic_vector(92, 8),
25837 => conv_std_logic_vector(92, 8),
25838 => conv_std_logic_vector(92, 8),
25839 => conv_std_logic_vector(93, 8),
25840 => conv_std_logic_vector(93, 8),
25841 => conv_std_logic_vector(94, 8),
25842 => conv_std_logic_vector(94, 8),
25843 => conv_std_logic_vector(94, 8),
25844 => conv_std_logic_vector(95, 8),
25845 => conv_std_logic_vector(95, 8),
25846 => conv_std_logic_vector(96, 8),
25847 => conv_std_logic_vector(96, 8),
25848 => conv_std_logic_vector(96, 8),
25849 => conv_std_logic_vector(97, 8),
25850 => conv_std_logic_vector(97, 8),
25851 => conv_std_logic_vector(98, 8),
25852 => conv_std_logic_vector(98, 8),
25853 => conv_std_logic_vector(98, 8),
25854 => conv_std_logic_vector(99, 8),
25855 => conv_std_logic_vector(99, 8),
25856 => conv_std_logic_vector(0, 8),
25857 => conv_std_logic_vector(0, 8),
25858 => conv_std_logic_vector(0, 8),
25859 => conv_std_logic_vector(1, 8),
25860 => conv_std_logic_vector(1, 8),
25861 => conv_std_logic_vector(1, 8),
25862 => conv_std_logic_vector(2, 8),
25863 => conv_std_logic_vector(2, 8),
25864 => conv_std_logic_vector(3, 8),
25865 => conv_std_logic_vector(3, 8),
25866 => conv_std_logic_vector(3, 8),
25867 => conv_std_logic_vector(4, 8),
25868 => conv_std_logic_vector(4, 8),
25869 => conv_std_logic_vector(5, 8),
25870 => conv_std_logic_vector(5, 8),
25871 => conv_std_logic_vector(5, 8),
25872 => conv_std_logic_vector(6, 8),
25873 => conv_std_logic_vector(6, 8),
25874 => conv_std_logic_vector(7, 8),
25875 => conv_std_logic_vector(7, 8),
25876 => conv_std_logic_vector(7, 8),
25877 => conv_std_logic_vector(8, 8),
25878 => conv_std_logic_vector(8, 8),
25879 => conv_std_logic_vector(9, 8),
25880 => conv_std_logic_vector(9, 8),
25881 => conv_std_logic_vector(9, 8),
25882 => conv_std_logic_vector(10, 8),
25883 => conv_std_logic_vector(10, 8),
25884 => conv_std_logic_vector(11, 8),
25885 => conv_std_logic_vector(11, 8),
25886 => conv_std_logic_vector(11, 8),
25887 => conv_std_logic_vector(12, 8),
25888 => conv_std_logic_vector(12, 8),
25889 => conv_std_logic_vector(13, 8),
25890 => conv_std_logic_vector(13, 8),
25891 => conv_std_logic_vector(13, 8),
25892 => conv_std_logic_vector(14, 8),
25893 => conv_std_logic_vector(14, 8),
25894 => conv_std_logic_vector(14, 8),
25895 => conv_std_logic_vector(15, 8),
25896 => conv_std_logic_vector(15, 8),
25897 => conv_std_logic_vector(16, 8),
25898 => conv_std_logic_vector(16, 8),
25899 => conv_std_logic_vector(16, 8),
25900 => conv_std_logic_vector(17, 8),
25901 => conv_std_logic_vector(17, 8),
25902 => conv_std_logic_vector(18, 8),
25903 => conv_std_logic_vector(18, 8),
25904 => conv_std_logic_vector(18, 8),
25905 => conv_std_logic_vector(19, 8),
25906 => conv_std_logic_vector(19, 8),
25907 => conv_std_logic_vector(20, 8),
25908 => conv_std_logic_vector(20, 8),
25909 => conv_std_logic_vector(20, 8),
25910 => conv_std_logic_vector(21, 8),
25911 => conv_std_logic_vector(21, 8),
25912 => conv_std_logic_vector(22, 8),
25913 => conv_std_logic_vector(22, 8),
25914 => conv_std_logic_vector(22, 8),
25915 => conv_std_logic_vector(23, 8),
25916 => conv_std_logic_vector(23, 8),
25917 => conv_std_logic_vector(24, 8),
25918 => conv_std_logic_vector(24, 8),
25919 => conv_std_logic_vector(24, 8),
25920 => conv_std_logic_vector(25, 8),
25921 => conv_std_logic_vector(25, 8),
25922 => conv_std_logic_vector(26, 8),
25923 => conv_std_logic_vector(26, 8),
25924 => conv_std_logic_vector(26, 8),
25925 => conv_std_logic_vector(27, 8),
25926 => conv_std_logic_vector(27, 8),
25927 => conv_std_logic_vector(28, 8),
25928 => conv_std_logic_vector(28, 8),
25929 => conv_std_logic_vector(28, 8),
25930 => conv_std_logic_vector(29, 8),
25931 => conv_std_logic_vector(29, 8),
25932 => conv_std_logic_vector(29, 8),
25933 => conv_std_logic_vector(30, 8),
25934 => conv_std_logic_vector(30, 8),
25935 => conv_std_logic_vector(31, 8),
25936 => conv_std_logic_vector(31, 8),
25937 => conv_std_logic_vector(31, 8),
25938 => conv_std_logic_vector(32, 8),
25939 => conv_std_logic_vector(32, 8),
25940 => conv_std_logic_vector(33, 8),
25941 => conv_std_logic_vector(33, 8),
25942 => conv_std_logic_vector(33, 8),
25943 => conv_std_logic_vector(34, 8),
25944 => conv_std_logic_vector(34, 8),
25945 => conv_std_logic_vector(35, 8),
25946 => conv_std_logic_vector(35, 8),
25947 => conv_std_logic_vector(35, 8),
25948 => conv_std_logic_vector(36, 8),
25949 => conv_std_logic_vector(36, 8),
25950 => conv_std_logic_vector(37, 8),
25951 => conv_std_logic_vector(37, 8),
25952 => conv_std_logic_vector(37, 8),
25953 => conv_std_logic_vector(38, 8),
25954 => conv_std_logic_vector(38, 8),
25955 => conv_std_logic_vector(39, 8),
25956 => conv_std_logic_vector(39, 8),
25957 => conv_std_logic_vector(39, 8),
25958 => conv_std_logic_vector(40, 8),
25959 => conv_std_logic_vector(40, 8),
25960 => conv_std_logic_vector(41, 8),
25961 => conv_std_logic_vector(41, 8),
25962 => conv_std_logic_vector(41, 8),
25963 => conv_std_logic_vector(42, 8),
25964 => conv_std_logic_vector(42, 8),
25965 => conv_std_logic_vector(43, 8),
25966 => conv_std_logic_vector(43, 8),
25967 => conv_std_logic_vector(43, 8),
25968 => conv_std_logic_vector(44, 8),
25969 => conv_std_logic_vector(44, 8),
25970 => conv_std_logic_vector(44, 8),
25971 => conv_std_logic_vector(45, 8),
25972 => conv_std_logic_vector(45, 8),
25973 => conv_std_logic_vector(46, 8),
25974 => conv_std_logic_vector(46, 8),
25975 => conv_std_logic_vector(46, 8),
25976 => conv_std_logic_vector(47, 8),
25977 => conv_std_logic_vector(47, 8),
25978 => conv_std_logic_vector(48, 8),
25979 => conv_std_logic_vector(48, 8),
25980 => conv_std_logic_vector(48, 8),
25981 => conv_std_logic_vector(49, 8),
25982 => conv_std_logic_vector(49, 8),
25983 => conv_std_logic_vector(50, 8),
25984 => conv_std_logic_vector(50, 8),
25985 => conv_std_logic_vector(50, 8),
25986 => conv_std_logic_vector(51, 8),
25987 => conv_std_logic_vector(51, 8),
25988 => conv_std_logic_vector(52, 8),
25989 => conv_std_logic_vector(52, 8),
25990 => conv_std_logic_vector(52, 8),
25991 => conv_std_logic_vector(53, 8),
25992 => conv_std_logic_vector(53, 8),
25993 => conv_std_logic_vector(54, 8),
25994 => conv_std_logic_vector(54, 8),
25995 => conv_std_logic_vector(54, 8),
25996 => conv_std_logic_vector(55, 8),
25997 => conv_std_logic_vector(55, 8),
25998 => conv_std_logic_vector(56, 8),
25999 => conv_std_logic_vector(56, 8),
26000 => conv_std_logic_vector(56, 8),
26001 => conv_std_logic_vector(57, 8),
26002 => conv_std_logic_vector(57, 8),
26003 => conv_std_logic_vector(57, 8),
26004 => conv_std_logic_vector(58, 8),
26005 => conv_std_logic_vector(58, 8),
26006 => conv_std_logic_vector(59, 8),
26007 => conv_std_logic_vector(59, 8),
26008 => conv_std_logic_vector(59, 8),
26009 => conv_std_logic_vector(60, 8),
26010 => conv_std_logic_vector(60, 8),
26011 => conv_std_logic_vector(61, 8),
26012 => conv_std_logic_vector(61, 8),
26013 => conv_std_logic_vector(61, 8),
26014 => conv_std_logic_vector(62, 8),
26015 => conv_std_logic_vector(62, 8),
26016 => conv_std_logic_vector(63, 8),
26017 => conv_std_logic_vector(63, 8),
26018 => conv_std_logic_vector(63, 8),
26019 => conv_std_logic_vector(64, 8),
26020 => conv_std_logic_vector(64, 8),
26021 => conv_std_logic_vector(65, 8),
26022 => conv_std_logic_vector(65, 8),
26023 => conv_std_logic_vector(65, 8),
26024 => conv_std_logic_vector(66, 8),
26025 => conv_std_logic_vector(66, 8),
26026 => conv_std_logic_vector(67, 8),
26027 => conv_std_logic_vector(67, 8),
26028 => conv_std_logic_vector(67, 8),
26029 => conv_std_logic_vector(68, 8),
26030 => conv_std_logic_vector(68, 8),
26031 => conv_std_logic_vector(69, 8),
26032 => conv_std_logic_vector(69, 8),
26033 => conv_std_logic_vector(69, 8),
26034 => conv_std_logic_vector(70, 8),
26035 => conv_std_logic_vector(70, 8),
26036 => conv_std_logic_vector(71, 8),
26037 => conv_std_logic_vector(71, 8),
26038 => conv_std_logic_vector(71, 8),
26039 => conv_std_logic_vector(72, 8),
26040 => conv_std_logic_vector(72, 8),
26041 => conv_std_logic_vector(72, 8),
26042 => conv_std_logic_vector(73, 8),
26043 => conv_std_logic_vector(73, 8),
26044 => conv_std_logic_vector(74, 8),
26045 => conv_std_logic_vector(74, 8),
26046 => conv_std_logic_vector(74, 8),
26047 => conv_std_logic_vector(75, 8),
26048 => conv_std_logic_vector(75, 8),
26049 => conv_std_logic_vector(76, 8),
26050 => conv_std_logic_vector(76, 8),
26051 => conv_std_logic_vector(76, 8),
26052 => conv_std_logic_vector(77, 8),
26053 => conv_std_logic_vector(77, 8),
26054 => conv_std_logic_vector(78, 8),
26055 => conv_std_logic_vector(78, 8),
26056 => conv_std_logic_vector(78, 8),
26057 => conv_std_logic_vector(79, 8),
26058 => conv_std_logic_vector(79, 8),
26059 => conv_std_logic_vector(80, 8),
26060 => conv_std_logic_vector(80, 8),
26061 => conv_std_logic_vector(80, 8),
26062 => conv_std_logic_vector(81, 8),
26063 => conv_std_logic_vector(81, 8),
26064 => conv_std_logic_vector(82, 8),
26065 => conv_std_logic_vector(82, 8),
26066 => conv_std_logic_vector(82, 8),
26067 => conv_std_logic_vector(83, 8),
26068 => conv_std_logic_vector(83, 8),
26069 => conv_std_logic_vector(84, 8),
26070 => conv_std_logic_vector(84, 8),
26071 => conv_std_logic_vector(84, 8),
26072 => conv_std_logic_vector(85, 8),
26073 => conv_std_logic_vector(85, 8),
26074 => conv_std_logic_vector(86, 8),
26075 => conv_std_logic_vector(86, 8),
26076 => conv_std_logic_vector(86, 8),
26077 => conv_std_logic_vector(87, 8),
26078 => conv_std_logic_vector(87, 8),
26079 => conv_std_logic_vector(87, 8),
26080 => conv_std_logic_vector(88, 8),
26081 => conv_std_logic_vector(88, 8),
26082 => conv_std_logic_vector(89, 8),
26083 => conv_std_logic_vector(89, 8),
26084 => conv_std_logic_vector(89, 8),
26085 => conv_std_logic_vector(90, 8),
26086 => conv_std_logic_vector(90, 8),
26087 => conv_std_logic_vector(91, 8),
26088 => conv_std_logic_vector(91, 8),
26089 => conv_std_logic_vector(91, 8),
26090 => conv_std_logic_vector(92, 8),
26091 => conv_std_logic_vector(92, 8),
26092 => conv_std_logic_vector(93, 8),
26093 => conv_std_logic_vector(93, 8),
26094 => conv_std_logic_vector(93, 8),
26095 => conv_std_logic_vector(94, 8),
26096 => conv_std_logic_vector(94, 8),
26097 => conv_std_logic_vector(95, 8),
26098 => conv_std_logic_vector(95, 8),
26099 => conv_std_logic_vector(95, 8),
26100 => conv_std_logic_vector(96, 8),
26101 => conv_std_logic_vector(96, 8),
26102 => conv_std_logic_vector(97, 8),
26103 => conv_std_logic_vector(97, 8),
26104 => conv_std_logic_vector(97, 8),
26105 => conv_std_logic_vector(98, 8),
26106 => conv_std_logic_vector(98, 8),
26107 => conv_std_logic_vector(99, 8),
26108 => conv_std_logic_vector(99, 8),
26109 => conv_std_logic_vector(99, 8),
26110 => conv_std_logic_vector(100, 8),
26111 => conv_std_logic_vector(100, 8),
26112 => conv_std_logic_vector(0, 8),
26113 => conv_std_logic_vector(0, 8),
26114 => conv_std_logic_vector(0, 8),
26115 => conv_std_logic_vector(1, 8),
26116 => conv_std_logic_vector(1, 8),
26117 => conv_std_logic_vector(1, 8),
26118 => conv_std_logic_vector(2, 8),
26119 => conv_std_logic_vector(2, 8),
26120 => conv_std_logic_vector(3, 8),
26121 => conv_std_logic_vector(3, 8),
26122 => conv_std_logic_vector(3, 8),
26123 => conv_std_logic_vector(4, 8),
26124 => conv_std_logic_vector(4, 8),
26125 => conv_std_logic_vector(5, 8),
26126 => conv_std_logic_vector(5, 8),
26127 => conv_std_logic_vector(5, 8),
26128 => conv_std_logic_vector(6, 8),
26129 => conv_std_logic_vector(6, 8),
26130 => conv_std_logic_vector(7, 8),
26131 => conv_std_logic_vector(7, 8),
26132 => conv_std_logic_vector(7, 8),
26133 => conv_std_logic_vector(8, 8),
26134 => conv_std_logic_vector(8, 8),
26135 => conv_std_logic_vector(9, 8),
26136 => conv_std_logic_vector(9, 8),
26137 => conv_std_logic_vector(9, 8),
26138 => conv_std_logic_vector(10, 8),
26139 => conv_std_logic_vector(10, 8),
26140 => conv_std_logic_vector(11, 8),
26141 => conv_std_logic_vector(11, 8),
26142 => conv_std_logic_vector(11, 8),
26143 => conv_std_logic_vector(12, 8),
26144 => conv_std_logic_vector(12, 8),
26145 => conv_std_logic_vector(13, 8),
26146 => conv_std_logic_vector(13, 8),
26147 => conv_std_logic_vector(13, 8),
26148 => conv_std_logic_vector(14, 8),
26149 => conv_std_logic_vector(14, 8),
26150 => conv_std_logic_vector(15, 8),
26151 => conv_std_logic_vector(15, 8),
26152 => conv_std_logic_vector(15, 8),
26153 => conv_std_logic_vector(16, 8),
26154 => conv_std_logic_vector(16, 8),
26155 => conv_std_logic_vector(17, 8),
26156 => conv_std_logic_vector(17, 8),
26157 => conv_std_logic_vector(17, 8),
26158 => conv_std_logic_vector(18, 8),
26159 => conv_std_logic_vector(18, 8),
26160 => conv_std_logic_vector(19, 8),
26161 => conv_std_logic_vector(19, 8),
26162 => conv_std_logic_vector(19, 8),
26163 => conv_std_logic_vector(20, 8),
26164 => conv_std_logic_vector(20, 8),
26165 => conv_std_logic_vector(21, 8),
26166 => conv_std_logic_vector(21, 8),
26167 => conv_std_logic_vector(21, 8),
26168 => conv_std_logic_vector(22, 8),
26169 => conv_std_logic_vector(22, 8),
26170 => conv_std_logic_vector(23, 8),
26171 => conv_std_logic_vector(23, 8),
26172 => conv_std_logic_vector(23, 8),
26173 => conv_std_logic_vector(24, 8),
26174 => conv_std_logic_vector(24, 8),
26175 => conv_std_logic_vector(25, 8),
26176 => conv_std_logic_vector(25, 8),
26177 => conv_std_logic_vector(25, 8),
26178 => conv_std_logic_vector(26, 8),
26179 => conv_std_logic_vector(26, 8),
26180 => conv_std_logic_vector(27, 8),
26181 => conv_std_logic_vector(27, 8),
26182 => conv_std_logic_vector(27, 8),
26183 => conv_std_logic_vector(28, 8),
26184 => conv_std_logic_vector(28, 8),
26185 => conv_std_logic_vector(29, 8),
26186 => conv_std_logic_vector(29, 8),
26187 => conv_std_logic_vector(29, 8),
26188 => conv_std_logic_vector(30, 8),
26189 => conv_std_logic_vector(30, 8),
26190 => conv_std_logic_vector(31, 8),
26191 => conv_std_logic_vector(31, 8),
26192 => conv_std_logic_vector(31, 8),
26193 => conv_std_logic_vector(32, 8),
26194 => conv_std_logic_vector(32, 8),
26195 => conv_std_logic_vector(33, 8),
26196 => conv_std_logic_vector(33, 8),
26197 => conv_std_logic_vector(33, 8),
26198 => conv_std_logic_vector(34, 8),
26199 => conv_std_logic_vector(34, 8),
26200 => conv_std_logic_vector(35, 8),
26201 => conv_std_logic_vector(35, 8),
26202 => conv_std_logic_vector(35, 8),
26203 => conv_std_logic_vector(36, 8),
26204 => conv_std_logic_vector(36, 8),
26205 => conv_std_logic_vector(37, 8),
26206 => conv_std_logic_vector(37, 8),
26207 => conv_std_logic_vector(37, 8),
26208 => conv_std_logic_vector(38, 8),
26209 => conv_std_logic_vector(38, 8),
26210 => conv_std_logic_vector(39, 8),
26211 => conv_std_logic_vector(39, 8),
26212 => conv_std_logic_vector(39, 8),
26213 => conv_std_logic_vector(40, 8),
26214 => conv_std_logic_vector(40, 8),
26215 => conv_std_logic_vector(41, 8),
26216 => conv_std_logic_vector(41, 8),
26217 => conv_std_logic_vector(41, 8),
26218 => conv_std_logic_vector(42, 8),
26219 => conv_std_logic_vector(42, 8),
26220 => conv_std_logic_vector(43, 8),
26221 => conv_std_logic_vector(43, 8),
26222 => conv_std_logic_vector(43, 8),
26223 => conv_std_logic_vector(44, 8),
26224 => conv_std_logic_vector(44, 8),
26225 => conv_std_logic_vector(45, 8),
26226 => conv_std_logic_vector(45, 8),
26227 => conv_std_logic_vector(45, 8),
26228 => conv_std_logic_vector(46, 8),
26229 => conv_std_logic_vector(46, 8),
26230 => conv_std_logic_vector(47, 8),
26231 => conv_std_logic_vector(47, 8),
26232 => conv_std_logic_vector(47, 8),
26233 => conv_std_logic_vector(48, 8),
26234 => conv_std_logic_vector(48, 8),
26235 => conv_std_logic_vector(49, 8),
26236 => conv_std_logic_vector(49, 8),
26237 => conv_std_logic_vector(49, 8),
26238 => conv_std_logic_vector(50, 8),
26239 => conv_std_logic_vector(50, 8),
26240 => conv_std_logic_vector(51, 8),
26241 => conv_std_logic_vector(51, 8),
26242 => conv_std_logic_vector(51, 8),
26243 => conv_std_logic_vector(52, 8),
26244 => conv_std_logic_vector(52, 8),
26245 => conv_std_logic_vector(52, 8),
26246 => conv_std_logic_vector(53, 8),
26247 => conv_std_logic_vector(53, 8),
26248 => conv_std_logic_vector(54, 8),
26249 => conv_std_logic_vector(54, 8),
26250 => conv_std_logic_vector(54, 8),
26251 => conv_std_logic_vector(55, 8),
26252 => conv_std_logic_vector(55, 8),
26253 => conv_std_logic_vector(56, 8),
26254 => conv_std_logic_vector(56, 8),
26255 => conv_std_logic_vector(56, 8),
26256 => conv_std_logic_vector(57, 8),
26257 => conv_std_logic_vector(57, 8),
26258 => conv_std_logic_vector(58, 8),
26259 => conv_std_logic_vector(58, 8),
26260 => conv_std_logic_vector(58, 8),
26261 => conv_std_logic_vector(59, 8),
26262 => conv_std_logic_vector(59, 8),
26263 => conv_std_logic_vector(60, 8),
26264 => conv_std_logic_vector(60, 8),
26265 => conv_std_logic_vector(60, 8),
26266 => conv_std_logic_vector(61, 8),
26267 => conv_std_logic_vector(61, 8),
26268 => conv_std_logic_vector(62, 8),
26269 => conv_std_logic_vector(62, 8),
26270 => conv_std_logic_vector(62, 8),
26271 => conv_std_logic_vector(63, 8),
26272 => conv_std_logic_vector(63, 8),
26273 => conv_std_logic_vector(64, 8),
26274 => conv_std_logic_vector(64, 8),
26275 => conv_std_logic_vector(64, 8),
26276 => conv_std_logic_vector(65, 8),
26277 => conv_std_logic_vector(65, 8),
26278 => conv_std_logic_vector(66, 8),
26279 => conv_std_logic_vector(66, 8),
26280 => conv_std_logic_vector(66, 8),
26281 => conv_std_logic_vector(67, 8),
26282 => conv_std_logic_vector(67, 8),
26283 => conv_std_logic_vector(68, 8),
26284 => conv_std_logic_vector(68, 8),
26285 => conv_std_logic_vector(68, 8),
26286 => conv_std_logic_vector(69, 8),
26287 => conv_std_logic_vector(69, 8),
26288 => conv_std_logic_vector(70, 8),
26289 => conv_std_logic_vector(70, 8),
26290 => conv_std_logic_vector(70, 8),
26291 => conv_std_logic_vector(71, 8),
26292 => conv_std_logic_vector(71, 8),
26293 => conv_std_logic_vector(72, 8),
26294 => conv_std_logic_vector(72, 8),
26295 => conv_std_logic_vector(72, 8),
26296 => conv_std_logic_vector(73, 8),
26297 => conv_std_logic_vector(73, 8),
26298 => conv_std_logic_vector(74, 8),
26299 => conv_std_logic_vector(74, 8),
26300 => conv_std_logic_vector(74, 8),
26301 => conv_std_logic_vector(75, 8),
26302 => conv_std_logic_vector(75, 8),
26303 => conv_std_logic_vector(76, 8),
26304 => conv_std_logic_vector(76, 8),
26305 => conv_std_logic_vector(76, 8),
26306 => conv_std_logic_vector(77, 8),
26307 => conv_std_logic_vector(77, 8),
26308 => conv_std_logic_vector(78, 8),
26309 => conv_std_logic_vector(78, 8),
26310 => conv_std_logic_vector(78, 8),
26311 => conv_std_logic_vector(79, 8),
26312 => conv_std_logic_vector(79, 8),
26313 => conv_std_logic_vector(80, 8),
26314 => conv_std_logic_vector(80, 8),
26315 => conv_std_logic_vector(80, 8),
26316 => conv_std_logic_vector(81, 8),
26317 => conv_std_logic_vector(81, 8),
26318 => conv_std_logic_vector(82, 8),
26319 => conv_std_logic_vector(82, 8),
26320 => conv_std_logic_vector(82, 8),
26321 => conv_std_logic_vector(83, 8),
26322 => conv_std_logic_vector(83, 8),
26323 => conv_std_logic_vector(84, 8),
26324 => conv_std_logic_vector(84, 8),
26325 => conv_std_logic_vector(84, 8),
26326 => conv_std_logic_vector(85, 8),
26327 => conv_std_logic_vector(85, 8),
26328 => conv_std_logic_vector(86, 8),
26329 => conv_std_logic_vector(86, 8),
26330 => conv_std_logic_vector(86, 8),
26331 => conv_std_logic_vector(87, 8),
26332 => conv_std_logic_vector(87, 8),
26333 => conv_std_logic_vector(88, 8),
26334 => conv_std_logic_vector(88, 8),
26335 => conv_std_logic_vector(88, 8),
26336 => conv_std_logic_vector(89, 8),
26337 => conv_std_logic_vector(89, 8),
26338 => conv_std_logic_vector(90, 8),
26339 => conv_std_logic_vector(90, 8),
26340 => conv_std_logic_vector(90, 8),
26341 => conv_std_logic_vector(91, 8),
26342 => conv_std_logic_vector(91, 8),
26343 => conv_std_logic_vector(92, 8),
26344 => conv_std_logic_vector(92, 8),
26345 => conv_std_logic_vector(92, 8),
26346 => conv_std_logic_vector(93, 8),
26347 => conv_std_logic_vector(93, 8),
26348 => conv_std_logic_vector(94, 8),
26349 => conv_std_logic_vector(94, 8),
26350 => conv_std_logic_vector(94, 8),
26351 => conv_std_logic_vector(95, 8),
26352 => conv_std_logic_vector(95, 8),
26353 => conv_std_logic_vector(96, 8),
26354 => conv_std_logic_vector(96, 8),
26355 => conv_std_logic_vector(96, 8),
26356 => conv_std_logic_vector(97, 8),
26357 => conv_std_logic_vector(97, 8),
26358 => conv_std_logic_vector(98, 8),
26359 => conv_std_logic_vector(98, 8),
26360 => conv_std_logic_vector(98, 8),
26361 => conv_std_logic_vector(99, 8),
26362 => conv_std_logic_vector(99, 8),
26363 => conv_std_logic_vector(100, 8),
26364 => conv_std_logic_vector(100, 8),
26365 => conv_std_logic_vector(100, 8),
26366 => conv_std_logic_vector(101, 8),
26367 => conv_std_logic_vector(101, 8),
26368 => conv_std_logic_vector(0, 8),
26369 => conv_std_logic_vector(0, 8),
26370 => conv_std_logic_vector(0, 8),
26371 => conv_std_logic_vector(1, 8),
26372 => conv_std_logic_vector(1, 8),
26373 => conv_std_logic_vector(2, 8),
26374 => conv_std_logic_vector(2, 8),
26375 => conv_std_logic_vector(2, 8),
26376 => conv_std_logic_vector(3, 8),
26377 => conv_std_logic_vector(3, 8),
26378 => conv_std_logic_vector(4, 8),
26379 => conv_std_logic_vector(4, 8),
26380 => conv_std_logic_vector(4, 8),
26381 => conv_std_logic_vector(5, 8),
26382 => conv_std_logic_vector(5, 8),
26383 => conv_std_logic_vector(6, 8),
26384 => conv_std_logic_vector(6, 8),
26385 => conv_std_logic_vector(6, 8),
26386 => conv_std_logic_vector(7, 8),
26387 => conv_std_logic_vector(7, 8),
26388 => conv_std_logic_vector(8, 8),
26389 => conv_std_logic_vector(8, 8),
26390 => conv_std_logic_vector(8, 8),
26391 => conv_std_logic_vector(9, 8),
26392 => conv_std_logic_vector(9, 8),
26393 => conv_std_logic_vector(10, 8),
26394 => conv_std_logic_vector(10, 8),
26395 => conv_std_logic_vector(10, 8),
26396 => conv_std_logic_vector(11, 8),
26397 => conv_std_logic_vector(11, 8),
26398 => conv_std_logic_vector(12, 8),
26399 => conv_std_logic_vector(12, 8),
26400 => conv_std_logic_vector(12, 8),
26401 => conv_std_logic_vector(13, 8),
26402 => conv_std_logic_vector(13, 8),
26403 => conv_std_logic_vector(14, 8),
26404 => conv_std_logic_vector(14, 8),
26405 => conv_std_logic_vector(14, 8),
26406 => conv_std_logic_vector(15, 8),
26407 => conv_std_logic_vector(15, 8),
26408 => conv_std_logic_vector(16, 8),
26409 => conv_std_logic_vector(16, 8),
26410 => conv_std_logic_vector(16, 8),
26411 => conv_std_logic_vector(17, 8),
26412 => conv_std_logic_vector(17, 8),
26413 => conv_std_logic_vector(18, 8),
26414 => conv_std_logic_vector(18, 8),
26415 => conv_std_logic_vector(18, 8),
26416 => conv_std_logic_vector(19, 8),
26417 => conv_std_logic_vector(19, 8),
26418 => conv_std_logic_vector(20, 8),
26419 => conv_std_logic_vector(20, 8),
26420 => conv_std_logic_vector(20, 8),
26421 => conv_std_logic_vector(21, 8),
26422 => conv_std_logic_vector(21, 8),
26423 => conv_std_logic_vector(22, 8),
26424 => conv_std_logic_vector(22, 8),
26425 => conv_std_logic_vector(22, 8),
26426 => conv_std_logic_vector(23, 8),
26427 => conv_std_logic_vector(23, 8),
26428 => conv_std_logic_vector(24, 8),
26429 => conv_std_logic_vector(24, 8),
26430 => conv_std_logic_vector(24, 8),
26431 => conv_std_logic_vector(25, 8),
26432 => conv_std_logic_vector(25, 8),
26433 => conv_std_logic_vector(26, 8),
26434 => conv_std_logic_vector(26, 8),
26435 => conv_std_logic_vector(26, 8),
26436 => conv_std_logic_vector(27, 8),
26437 => conv_std_logic_vector(27, 8),
26438 => conv_std_logic_vector(28, 8),
26439 => conv_std_logic_vector(28, 8),
26440 => conv_std_logic_vector(28, 8),
26441 => conv_std_logic_vector(29, 8),
26442 => conv_std_logic_vector(29, 8),
26443 => conv_std_logic_vector(30, 8),
26444 => conv_std_logic_vector(30, 8),
26445 => conv_std_logic_vector(30, 8),
26446 => conv_std_logic_vector(31, 8),
26447 => conv_std_logic_vector(31, 8),
26448 => conv_std_logic_vector(32, 8),
26449 => conv_std_logic_vector(32, 8),
26450 => conv_std_logic_vector(32, 8),
26451 => conv_std_logic_vector(33, 8),
26452 => conv_std_logic_vector(33, 8),
26453 => conv_std_logic_vector(34, 8),
26454 => conv_std_logic_vector(34, 8),
26455 => conv_std_logic_vector(35, 8),
26456 => conv_std_logic_vector(35, 8),
26457 => conv_std_logic_vector(35, 8),
26458 => conv_std_logic_vector(36, 8),
26459 => conv_std_logic_vector(36, 8),
26460 => conv_std_logic_vector(37, 8),
26461 => conv_std_logic_vector(37, 8),
26462 => conv_std_logic_vector(37, 8),
26463 => conv_std_logic_vector(38, 8),
26464 => conv_std_logic_vector(38, 8),
26465 => conv_std_logic_vector(39, 8),
26466 => conv_std_logic_vector(39, 8),
26467 => conv_std_logic_vector(39, 8),
26468 => conv_std_logic_vector(40, 8),
26469 => conv_std_logic_vector(40, 8),
26470 => conv_std_logic_vector(41, 8),
26471 => conv_std_logic_vector(41, 8),
26472 => conv_std_logic_vector(41, 8),
26473 => conv_std_logic_vector(42, 8),
26474 => conv_std_logic_vector(42, 8),
26475 => conv_std_logic_vector(43, 8),
26476 => conv_std_logic_vector(43, 8),
26477 => conv_std_logic_vector(43, 8),
26478 => conv_std_logic_vector(44, 8),
26479 => conv_std_logic_vector(44, 8),
26480 => conv_std_logic_vector(45, 8),
26481 => conv_std_logic_vector(45, 8),
26482 => conv_std_logic_vector(45, 8),
26483 => conv_std_logic_vector(46, 8),
26484 => conv_std_logic_vector(46, 8),
26485 => conv_std_logic_vector(47, 8),
26486 => conv_std_logic_vector(47, 8),
26487 => conv_std_logic_vector(47, 8),
26488 => conv_std_logic_vector(48, 8),
26489 => conv_std_logic_vector(48, 8),
26490 => conv_std_logic_vector(49, 8),
26491 => conv_std_logic_vector(49, 8),
26492 => conv_std_logic_vector(49, 8),
26493 => conv_std_logic_vector(50, 8),
26494 => conv_std_logic_vector(50, 8),
26495 => conv_std_logic_vector(51, 8),
26496 => conv_std_logic_vector(51, 8),
26497 => conv_std_logic_vector(51, 8),
26498 => conv_std_logic_vector(52, 8),
26499 => conv_std_logic_vector(52, 8),
26500 => conv_std_logic_vector(53, 8),
26501 => conv_std_logic_vector(53, 8),
26502 => conv_std_logic_vector(53, 8),
26503 => conv_std_logic_vector(54, 8),
26504 => conv_std_logic_vector(54, 8),
26505 => conv_std_logic_vector(55, 8),
26506 => conv_std_logic_vector(55, 8),
26507 => conv_std_logic_vector(55, 8),
26508 => conv_std_logic_vector(56, 8),
26509 => conv_std_logic_vector(56, 8),
26510 => conv_std_logic_vector(57, 8),
26511 => conv_std_logic_vector(57, 8),
26512 => conv_std_logic_vector(57, 8),
26513 => conv_std_logic_vector(58, 8),
26514 => conv_std_logic_vector(58, 8),
26515 => conv_std_logic_vector(59, 8),
26516 => conv_std_logic_vector(59, 8),
26517 => conv_std_logic_vector(59, 8),
26518 => conv_std_logic_vector(60, 8),
26519 => conv_std_logic_vector(60, 8),
26520 => conv_std_logic_vector(61, 8),
26521 => conv_std_logic_vector(61, 8),
26522 => conv_std_logic_vector(61, 8),
26523 => conv_std_logic_vector(62, 8),
26524 => conv_std_logic_vector(62, 8),
26525 => conv_std_logic_vector(63, 8),
26526 => conv_std_logic_vector(63, 8),
26527 => conv_std_logic_vector(63, 8),
26528 => conv_std_logic_vector(64, 8),
26529 => conv_std_logic_vector(64, 8),
26530 => conv_std_logic_vector(65, 8),
26531 => conv_std_logic_vector(65, 8),
26532 => conv_std_logic_vector(65, 8),
26533 => conv_std_logic_vector(66, 8),
26534 => conv_std_logic_vector(66, 8),
26535 => conv_std_logic_vector(67, 8),
26536 => conv_std_logic_vector(67, 8),
26537 => conv_std_logic_vector(67, 8),
26538 => conv_std_logic_vector(68, 8),
26539 => conv_std_logic_vector(68, 8),
26540 => conv_std_logic_vector(69, 8),
26541 => conv_std_logic_vector(69, 8),
26542 => conv_std_logic_vector(70, 8),
26543 => conv_std_logic_vector(70, 8),
26544 => conv_std_logic_vector(70, 8),
26545 => conv_std_logic_vector(71, 8),
26546 => conv_std_logic_vector(71, 8),
26547 => conv_std_logic_vector(72, 8),
26548 => conv_std_logic_vector(72, 8),
26549 => conv_std_logic_vector(72, 8),
26550 => conv_std_logic_vector(73, 8),
26551 => conv_std_logic_vector(73, 8),
26552 => conv_std_logic_vector(74, 8),
26553 => conv_std_logic_vector(74, 8),
26554 => conv_std_logic_vector(74, 8),
26555 => conv_std_logic_vector(75, 8),
26556 => conv_std_logic_vector(75, 8),
26557 => conv_std_logic_vector(76, 8),
26558 => conv_std_logic_vector(76, 8),
26559 => conv_std_logic_vector(76, 8),
26560 => conv_std_logic_vector(77, 8),
26561 => conv_std_logic_vector(77, 8),
26562 => conv_std_logic_vector(78, 8),
26563 => conv_std_logic_vector(78, 8),
26564 => conv_std_logic_vector(78, 8),
26565 => conv_std_logic_vector(79, 8),
26566 => conv_std_logic_vector(79, 8),
26567 => conv_std_logic_vector(80, 8),
26568 => conv_std_logic_vector(80, 8),
26569 => conv_std_logic_vector(80, 8),
26570 => conv_std_logic_vector(81, 8),
26571 => conv_std_logic_vector(81, 8),
26572 => conv_std_logic_vector(82, 8),
26573 => conv_std_logic_vector(82, 8),
26574 => conv_std_logic_vector(82, 8),
26575 => conv_std_logic_vector(83, 8),
26576 => conv_std_logic_vector(83, 8),
26577 => conv_std_logic_vector(84, 8),
26578 => conv_std_logic_vector(84, 8),
26579 => conv_std_logic_vector(84, 8),
26580 => conv_std_logic_vector(85, 8),
26581 => conv_std_logic_vector(85, 8),
26582 => conv_std_logic_vector(86, 8),
26583 => conv_std_logic_vector(86, 8),
26584 => conv_std_logic_vector(86, 8),
26585 => conv_std_logic_vector(87, 8),
26586 => conv_std_logic_vector(87, 8),
26587 => conv_std_logic_vector(88, 8),
26588 => conv_std_logic_vector(88, 8),
26589 => conv_std_logic_vector(88, 8),
26590 => conv_std_logic_vector(89, 8),
26591 => conv_std_logic_vector(89, 8),
26592 => conv_std_logic_vector(90, 8),
26593 => conv_std_logic_vector(90, 8),
26594 => conv_std_logic_vector(90, 8),
26595 => conv_std_logic_vector(91, 8),
26596 => conv_std_logic_vector(91, 8),
26597 => conv_std_logic_vector(92, 8),
26598 => conv_std_logic_vector(92, 8),
26599 => conv_std_logic_vector(92, 8),
26600 => conv_std_logic_vector(93, 8),
26601 => conv_std_logic_vector(93, 8),
26602 => conv_std_logic_vector(94, 8),
26603 => conv_std_logic_vector(94, 8),
26604 => conv_std_logic_vector(94, 8),
26605 => conv_std_logic_vector(95, 8),
26606 => conv_std_logic_vector(95, 8),
26607 => conv_std_logic_vector(96, 8),
26608 => conv_std_logic_vector(96, 8),
26609 => conv_std_logic_vector(96, 8),
26610 => conv_std_logic_vector(97, 8),
26611 => conv_std_logic_vector(97, 8),
26612 => conv_std_logic_vector(98, 8),
26613 => conv_std_logic_vector(98, 8),
26614 => conv_std_logic_vector(98, 8),
26615 => conv_std_logic_vector(99, 8),
26616 => conv_std_logic_vector(99, 8),
26617 => conv_std_logic_vector(100, 8),
26618 => conv_std_logic_vector(100, 8),
26619 => conv_std_logic_vector(100, 8),
26620 => conv_std_logic_vector(101, 8),
26621 => conv_std_logic_vector(101, 8),
26622 => conv_std_logic_vector(102, 8),
26623 => conv_std_logic_vector(102, 8),
26624 => conv_std_logic_vector(0, 8),
26625 => conv_std_logic_vector(0, 8),
26626 => conv_std_logic_vector(0, 8),
26627 => conv_std_logic_vector(1, 8),
26628 => conv_std_logic_vector(1, 8),
26629 => conv_std_logic_vector(2, 8),
26630 => conv_std_logic_vector(2, 8),
26631 => conv_std_logic_vector(2, 8),
26632 => conv_std_logic_vector(3, 8),
26633 => conv_std_logic_vector(3, 8),
26634 => conv_std_logic_vector(4, 8),
26635 => conv_std_logic_vector(4, 8),
26636 => conv_std_logic_vector(4, 8),
26637 => conv_std_logic_vector(5, 8),
26638 => conv_std_logic_vector(5, 8),
26639 => conv_std_logic_vector(6, 8),
26640 => conv_std_logic_vector(6, 8),
26641 => conv_std_logic_vector(6, 8),
26642 => conv_std_logic_vector(7, 8),
26643 => conv_std_logic_vector(7, 8),
26644 => conv_std_logic_vector(8, 8),
26645 => conv_std_logic_vector(8, 8),
26646 => conv_std_logic_vector(8, 8),
26647 => conv_std_logic_vector(9, 8),
26648 => conv_std_logic_vector(9, 8),
26649 => conv_std_logic_vector(10, 8),
26650 => conv_std_logic_vector(10, 8),
26651 => conv_std_logic_vector(10, 8),
26652 => conv_std_logic_vector(11, 8),
26653 => conv_std_logic_vector(11, 8),
26654 => conv_std_logic_vector(12, 8),
26655 => conv_std_logic_vector(12, 8),
26656 => conv_std_logic_vector(13, 8),
26657 => conv_std_logic_vector(13, 8),
26658 => conv_std_logic_vector(13, 8),
26659 => conv_std_logic_vector(14, 8),
26660 => conv_std_logic_vector(14, 8),
26661 => conv_std_logic_vector(15, 8),
26662 => conv_std_logic_vector(15, 8),
26663 => conv_std_logic_vector(15, 8),
26664 => conv_std_logic_vector(16, 8),
26665 => conv_std_logic_vector(16, 8),
26666 => conv_std_logic_vector(17, 8),
26667 => conv_std_logic_vector(17, 8),
26668 => conv_std_logic_vector(17, 8),
26669 => conv_std_logic_vector(18, 8),
26670 => conv_std_logic_vector(18, 8),
26671 => conv_std_logic_vector(19, 8),
26672 => conv_std_logic_vector(19, 8),
26673 => conv_std_logic_vector(19, 8),
26674 => conv_std_logic_vector(20, 8),
26675 => conv_std_logic_vector(20, 8),
26676 => conv_std_logic_vector(21, 8),
26677 => conv_std_logic_vector(21, 8),
26678 => conv_std_logic_vector(21, 8),
26679 => conv_std_logic_vector(22, 8),
26680 => conv_std_logic_vector(22, 8),
26681 => conv_std_logic_vector(23, 8),
26682 => conv_std_logic_vector(23, 8),
26683 => conv_std_logic_vector(23, 8),
26684 => conv_std_logic_vector(24, 8),
26685 => conv_std_logic_vector(24, 8),
26686 => conv_std_logic_vector(25, 8),
26687 => conv_std_logic_vector(25, 8),
26688 => conv_std_logic_vector(26, 8),
26689 => conv_std_logic_vector(26, 8),
26690 => conv_std_logic_vector(26, 8),
26691 => conv_std_logic_vector(27, 8),
26692 => conv_std_logic_vector(27, 8),
26693 => conv_std_logic_vector(28, 8),
26694 => conv_std_logic_vector(28, 8),
26695 => conv_std_logic_vector(28, 8),
26696 => conv_std_logic_vector(29, 8),
26697 => conv_std_logic_vector(29, 8),
26698 => conv_std_logic_vector(30, 8),
26699 => conv_std_logic_vector(30, 8),
26700 => conv_std_logic_vector(30, 8),
26701 => conv_std_logic_vector(31, 8),
26702 => conv_std_logic_vector(31, 8),
26703 => conv_std_logic_vector(32, 8),
26704 => conv_std_logic_vector(32, 8),
26705 => conv_std_logic_vector(32, 8),
26706 => conv_std_logic_vector(33, 8),
26707 => conv_std_logic_vector(33, 8),
26708 => conv_std_logic_vector(34, 8),
26709 => conv_std_logic_vector(34, 8),
26710 => conv_std_logic_vector(34, 8),
26711 => conv_std_logic_vector(35, 8),
26712 => conv_std_logic_vector(35, 8),
26713 => conv_std_logic_vector(36, 8),
26714 => conv_std_logic_vector(36, 8),
26715 => conv_std_logic_vector(36, 8),
26716 => conv_std_logic_vector(37, 8),
26717 => conv_std_logic_vector(37, 8),
26718 => conv_std_logic_vector(38, 8),
26719 => conv_std_logic_vector(38, 8),
26720 => conv_std_logic_vector(39, 8),
26721 => conv_std_logic_vector(39, 8),
26722 => conv_std_logic_vector(39, 8),
26723 => conv_std_logic_vector(40, 8),
26724 => conv_std_logic_vector(40, 8),
26725 => conv_std_logic_vector(41, 8),
26726 => conv_std_logic_vector(41, 8),
26727 => conv_std_logic_vector(41, 8),
26728 => conv_std_logic_vector(42, 8),
26729 => conv_std_logic_vector(42, 8),
26730 => conv_std_logic_vector(43, 8),
26731 => conv_std_logic_vector(43, 8),
26732 => conv_std_logic_vector(43, 8),
26733 => conv_std_logic_vector(44, 8),
26734 => conv_std_logic_vector(44, 8),
26735 => conv_std_logic_vector(45, 8),
26736 => conv_std_logic_vector(45, 8),
26737 => conv_std_logic_vector(45, 8),
26738 => conv_std_logic_vector(46, 8),
26739 => conv_std_logic_vector(46, 8),
26740 => conv_std_logic_vector(47, 8),
26741 => conv_std_logic_vector(47, 8),
26742 => conv_std_logic_vector(47, 8),
26743 => conv_std_logic_vector(48, 8),
26744 => conv_std_logic_vector(48, 8),
26745 => conv_std_logic_vector(49, 8),
26746 => conv_std_logic_vector(49, 8),
26747 => conv_std_logic_vector(49, 8),
26748 => conv_std_logic_vector(50, 8),
26749 => conv_std_logic_vector(50, 8),
26750 => conv_std_logic_vector(51, 8),
26751 => conv_std_logic_vector(51, 8),
26752 => conv_std_logic_vector(52, 8),
26753 => conv_std_logic_vector(52, 8),
26754 => conv_std_logic_vector(52, 8),
26755 => conv_std_logic_vector(53, 8),
26756 => conv_std_logic_vector(53, 8),
26757 => conv_std_logic_vector(54, 8),
26758 => conv_std_logic_vector(54, 8),
26759 => conv_std_logic_vector(54, 8),
26760 => conv_std_logic_vector(55, 8),
26761 => conv_std_logic_vector(55, 8),
26762 => conv_std_logic_vector(56, 8),
26763 => conv_std_logic_vector(56, 8),
26764 => conv_std_logic_vector(56, 8),
26765 => conv_std_logic_vector(57, 8),
26766 => conv_std_logic_vector(57, 8),
26767 => conv_std_logic_vector(58, 8),
26768 => conv_std_logic_vector(58, 8),
26769 => conv_std_logic_vector(58, 8),
26770 => conv_std_logic_vector(59, 8),
26771 => conv_std_logic_vector(59, 8),
26772 => conv_std_logic_vector(60, 8),
26773 => conv_std_logic_vector(60, 8),
26774 => conv_std_logic_vector(60, 8),
26775 => conv_std_logic_vector(61, 8),
26776 => conv_std_logic_vector(61, 8),
26777 => conv_std_logic_vector(62, 8),
26778 => conv_std_logic_vector(62, 8),
26779 => conv_std_logic_vector(62, 8),
26780 => conv_std_logic_vector(63, 8),
26781 => conv_std_logic_vector(63, 8),
26782 => conv_std_logic_vector(64, 8),
26783 => conv_std_logic_vector(64, 8),
26784 => conv_std_logic_vector(65, 8),
26785 => conv_std_logic_vector(65, 8),
26786 => conv_std_logic_vector(65, 8),
26787 => conv_std_logic_vector(66, 8),
26788 => conv_std_logic_vector(66, 8),
26789 => conv_std_logic_vector(67, 8),
26790 => conv_std_logic_vector(67, 8),
26791 => conv_std_logic_vector(67, 8),
26792 => conv_std_logic_vector(68, 8),
26793 => conv_std_logic_vector(68, 8),
26794 => conv_std_logic_vector(69, 8),
26795 => conv_std_logic_vector(69, 8),
26796 => conv_std_logic_vector(69, 8),
26797 => conv_std_logic_vector(70, 8),
26798 => conv_std_logic_vector(70, 8),
26799 => conv_std_logic_vector(71, 8),
26800 => conv_std_logic_vector(71, 8),
26801 => conv_std_logic_vector(71, 8),
26802 => conv_std_logic_vector(72, 8),
26803 => conv_std_logic_vector(72, 8),
26804 => conv_std_logic_vector(73, 8),
26805 => conv_std_logic_vector(73, 8),
26806 => conv_std_logic_vector(73, 8),
26807 => conv_std_logic_vector(74, 8),
26808 => conv_std_logic_vector(74, 8),
26809 => conv_std_logic_vector(75, 8),
26810 => conv_std_logic_vector(75, 8),
26811 => conv_std_logic_vector(75, 8),
26812 => conv_std_logic_vector(76, 8),
26813 => conv_std_logic_vector(76, 8),
26814 => conv_std_logic_vector(77, 8),
26815 => conv_std_logic_vector(77, 8),
26816 => conv_std_logic_vector(78, 8),
26817 => conv_std_logic_vector(78, 8),
26818 => conv_std_logic_vector(78, 8),
26819 => conv_std_logic_vector(79, 8),
26820 => conv_std_logic_vector(79, 8),
26821 => conv_std_logic_vector(80, 8),
26822 => conv_std_logic_vector(80, 8),
26823 => conv_std_logic_vector(80, 8),
26824 => conv_std_logic_vector(81, 8),
26825 => conv_std_logic_vector(81, 8),
26826 => conv_std_logic_vector(82, 8),
26827 => conv_std_logic_vector(82, 8),
26828 => conv_std_logic_vector(82, 8),
26829 => conv_std_logic_vector(83, 8),
26830 => conv_std_logic_vector(83, 8),
26831 => conv_std_logic_vector(84, 8),
26832 => conv_std_logic_vector(84, 8),
26833 => conv_std_logic_vector(84, 8),
26834 => conv_std_logic_vector(85, 8),
26835 => conv_std_logic_vector(85, 8),
26836 => conv_std_logic_vector(86, 8),
26837 => conv_std_logic_vector(86, 8),
26838 => conv_std_logic_vector(86, 8),
26839 => conv_std_logic_vector(87, 8),
26840 => conv_std_logic_vector(87, 8),
26841 => conv_std_logic_vector(88, 8),
26842 => conv_std_logic_vector(88, 8),
26843 => conv_std_logic_vector(88, 8),
26844 => conv_std_logic_vector(89, 8),
26845 => conv_std_logic_vector(89, 8),
26846 => conv_std_logic_vector(90, 8),
26847 => conv_std_logic_vector(90, 8),
26848 => conv_std_logic_vector(91, 8),
26849 => conv_std_logic_vector(91, 8),
26850 => conv_std_logic_vector(91, 8),
26851 => conv_std_logic_vector(92, 8),
26852 => conv_std_logic_vector(92, 8),
26853 => conv_std_logic_vector(93, 8),
26854 => conv_std_logic_vector(93, 8),
26855 => conv_std_logic_vector(93, 8),
26856 => conv_std_logic_vector(94, 8),
26857 => conv_std_logic_vector(94, 8),
26858 => conv_std_logic_vector(95, 8),
26859 => conv_std_logic_vector(95, 8),
26860 => conv_std_logic_vector(95, 8),
26861 => conv_std_logic_vector(96, 8),
26862 => conv_std_logic_vector(96, 8),
26863 => conv_std_logic_vector(97, 8),
26864 => conv_std_logic_vector(97, 8),
26865 => conv_std_logic_vector(97, 8),
26866 => conv_std_logic_vector(98, 8),
26867 => conv_std_logic_vector(98, 8),
26868 => conv_std_logic_vector(99, 8),
26869 => conv_std_logic_vector(99, 8),
26870 => conv_std_logic_vector(99, 8),
26871 => conv_std_logic_vector(100, 8),
26872 => conv_std_logic_vector(100, 8),
26873 => conv_std_logic_vector(101, 8),
26874 => conv_std_logic_vector(101, 8),
26875 => conv_std_logic_vector(101, 8),
26876 => conv_std_logic_vector(102, 8),
26877 => conv_std_logic_vector(102, 8),
26878 => conv_std_logic_vector(103, 8),
26879 => conv_std_logic_vector(103, 8),
26880 => conv_std_logic_vector(0, 8),
26881 => conv_std_logic_vector(0, 8),
26882 => conv_std_logic_vector(0, 8),
26883 => conv_std_logic_vector(1, 8),
26884 => conv_std_logic_vector(1, 8),
26885 => conv_std_logic_vector(2, 8),
26886 => conv_std_logic_vector(2, 8),
26887 => conv_std_logic_vector(2, 8),
26888 => conv_std_logic_vector(3, 8),
26889 => conv_std_logic_vector(3, 8),
26890 => conv_std_logic_vector(4, 8),
26891 => conv_std_logic_vector(4, 8),
26892 => conv_std_logic_vector(4, 8),
26893 => conv_std_logic_vector(5, 8),
26894 => conv_std_logic_vector(5, 8),
26895 => conv_std_logic_vector(6, 8),
26896 => conv_std_logic_vector(6, 8),
26897 => conv_std_logic_vector(6, 8),
26898 => conv_std_logic_vector(7, 8),
26899 => conv_std_logic_vector(7, 8),
26900 => conv_std_logic_vector(8, 8),
26901 => conv_std_logic_vector(8, 8),
26902 => conv_std_logic_vector(9, 8),
26903 => conv_std_logic_vector(9, 8),
26904 => conv_std_logic_vector(9, 8),
26905 => conv_std_logic_vector(10, 8),
26906 => conv_std_logic_vector(10, 8),
26907 => conv_std_logic_vector(11, 8),
26908 => conv_std_logic_vector(11, 8),
26909 => conv_std_logic_vector(11, 8),
26910 => conv_std_logic_vector(12, 8),
26911 => conv_std_logic_vector(12, 8),
26912 => conv_std_logic_vector(13, 8),
26913 => conv_std_logic_vector(13, 8),
26914 => conv_std_logic_vector(13, 8),
26915 => conv_std_logic_vector(14, 8),
26916 => conv_std_logic_vector(14, 8),
26917 => conv_std_logic_vector(15, 8),
26918 => conv_std_logic_vector(15, 8),
26919 => conv_std_logic_vector(15, 8),
26920 => conv_std_logic_vector(16, 8),
26921 => conv_std_logic_vector(16, 8),
26922 => conv_std_logic_vector(17, 8),
26923 => conv_std_logic_vector(17, 8),
26924 => conv_std_logic_vector(18, 8),
26925 => conv_std_logic_vector(18, 8),
26926 => conv_std_logic_vector(18, 8),
26927 => conv_std_logic_vector(19, 8),
26928 => conv_std_logic_vector(19, 8),
26929 => conv_std_logic_vector(20, 8),
26930 => conv_std_logic_vector(20, 8),
26931 => conv_std_logic_vector(20, 8),
26932 => conv_std_logic_vector(21, 8),
26933 => conv_std_logic_vector(21, 8),
26934 => conv_std_logic_vector(22, 8),
26935 => conv_std_logic_vector(22, 8),
26936 => conv_std_logic_vector(22, 8),
26937 => conv_std_logic_vector(23, 8),
26938 => conv_std_logic_vector(23, 8),
26939 => conv_std_logic_vector(24, 8),
26940 => conv_std_logic_vector(24, 8),
26941 => conv_std_logic_vector(25, 8),
26942 => conv_std_logic_vector(25, 8),
26943 => conv_std_logic_vector(25, 8),
26944 => conv_std_logic_vector(26, 8),
26945 => conv_std_logic_vector(26, 8),
26946 => conv_std_logic_vector(27, 8),
26947 => conv_std_logic_vector(27, 8),
26948 => conv_std_logic_vector(27, 8),
26949 => conv_std_logic_vector(28, 8),
26950 => conv_std_logic_vector(28, 8),
26951 => conv_std_logic_vector(29, 8),
26952 => conv_std_logic_vector(29, 8),
26953 => conv_std_logic_vector(29, 8),
26954 => conv_std_logic_vector(30, 8),
26955 => conv_std_logic_vector(30, 8),
26956 => conv_std_logic_vector(31, 8),
26957 => conv_std_logic_vector(31, 8),
26958 => conv_std_logic_vector(31, 8),
26959 => conv_std_logic_vector(32, 8),
26960 => conv_std_logic_vector(32, 8),
26961 => conv_std_logic_vector(33, 8),
26962 => conv_std_logic_vector(33, 8),
26963 => conv_std_logic_vector(34, 8),
26964 => conv_std_logic_vector(34, 8),
26965 => conv_std_logic_vector(34, 8),
26966 => conv_std_logic_vector(35, 8),
26967 => conv_std_logic_vector(35, 8),
26968 => conv_std_logic_vector(36, 8),
26969 => conv_std_logic_vector(36, 8),
26970 => conv_std_logic_vector(36, 8),
26971 => conv_std_logic_vector(37, 8),
26972 => conv_std_logic_vector(37, 8),
26973 => conv_std_logic_vector(38, 8),
26974 => conv_std_logic_vector(38, 8),
26975 => conv_std_logic_vector(38, 8),
26976 => conv_std_logic_vector(39, 8),
26977 => conv_std_logic_vector(39, 8),
26978 => conv_std_logic_vector(40, 8),
26979 => conv_std_logic_vector(40, 8),
26980 => conv_std_logic_vector(41, 8),
26981 => conv_std_logic_vector(41, 8),
26982 => conv_std_logic_vector(41, 8),
26983 => conv_std_logic_vector(42, 8),
26984 => conv_std_logic_vector(42, 8),
26985 => conv_std_logic_vector(43, 8),
26986 => conv_std_logic_vector(43, 8),
26987 => conv_std_logic_vector(43, 8),
26988 => conv_std_logic_vector(44, 8),
26989 => conv_std_logic_vector(44, 8),
26990 => conv_std_logic_vector(45, 8),
26991 => conv_std_logic_vector(45, 8),
26992 => conv_std_logic_vector(45, 8),
26993 => conv_std_logic_vector(46, 8),
26994 => conv_std_logic_vector(46, 8),
26995 => conv_std_logic_vector(47, 8),
26996 => conv_std_logic_vector(47, 8),
26997 => conv_std_logic_vector(47, 8),
26998 => conv_std_logic_vector(48, 8),
26999 => conv_std_logic_vector(48, 8),
27000 => conv_std_logic_vector(49, 8),
27001 => conv_std_logic_vector(49, 8),
27002 => conv_std_logic_vector(50, 8),
27003 => conv_std_logic_vector(50, 8),
27004 => conv_std_logic_vector(50, 8),
27005 => conv_std_logic_vector(51, 8),
27006 => conv_std_logic_vector(51, 8),
27007 => conv_std_logic_vector(52, 8),
27008 => conv_std_logic_vector(52, 8),
27009 => conv_std_logic_vector(52, 8),
27010 => conv_std_logic_vector(53, 8),
27011 => conv_std_logic_vector(53, 8),
27012 => conv_std_logic_vector(54, 8),
27013 => conv_std_logic_vector(54, 8),
27014 => conv_std_logic_vector(54, 8),
27015 => conv_std_logic_vector(55, 8),
27016 => conv_std_logic_vector(55, 8),
27017 => conv_std_logic_vector(56, 8),
27018 => conv_std_logic_vector(56, 8),
27019 => conv_std_logic_vector(57, 8),
27020 => conv_std_logic_vector(57, 8),
27021 => conv_std_logic_vector(57, 8),
27022 => conv_std_logic_vector(58, 8),
27023 => conv_std_logic_vector(58, 8),
27024 => conv_std_logic_vector(59, 8),
27025 => conv_std_logic_vector(59, 8),
27026 => conv_std_logic_vector(59, 8),
27027 => conv_std_logic_vector(60, 8),
27028 => conv_std_logic_vector(60, 8),
27029 => conv_std_logic_vector(61, 8),
27030 => conv_std_logic_vector(61, 8),
27031 => conv_std_logic_vector(61, 8),
27032 => conv_std_logic_vector(62, 8),
27033 => conv_std_logic_vector(62, 8),
27034 => conv_std_logic_vector(63, 8),
27035 => conv_std_logic_vector(63, 8),
27036 => conv_std_logic_vector(63, 8),
27037 => conv_std_logic_vector(64, 8),
27038 => conv_std_logic_vector(64, 8),
27039 => conv_std_logic_vector(65, 8),
27040 => conv_std_logic_vector(65, 8),
27041 => conv_std_logic_vector(66, 8),
27042 => conv_std_logic_vector(66, 8),
27043 => conv_std_logic_vector(66, 8),
27044 => conv_std_logic_vector(67, 8),
27045 => conv_std_logic_vector(67, 8),
27046 => conv_std_logic_vector(68, 8),
27047 => conv_std_logic_vector(68, 8),
27048 => conv_std_logic_vector(68, 8),
27049 => conv_std_logic_vector(69, 8),
27050 => conv_std_logic_vector(69, 8),
27051 => conv_std_logic_vector(70, 8),
27052 => conv_std_logic_vector(70, 8),
27053 => conv_std_logic_vector(70, 8),
27054 => conv_std_logic_vector(71, 8),
27055 => conv_std_logic_vector(71, 8),
27056 => conv_std_logic_vector(72, 8),
27057 => conv_std_logic_vector(72, 8),
27058 => conv_std_logic_vector(73, 8),
27059 => conv_std_logic_vector(73, 8),
27060 => conv_std_logic_vector(73, 8),
27061 => conv_std_logic_vector(74, 8),
27062 => conv_std_logic_vector(74, 8),
27063 => conv_std_logic_vector(75, 8),
27064 => conv_std_logic_vector(75, 8),
27065 => conv_std_logic_vector(75, 8),
27066 => conv_std_logic_vector(76, 8),
27067 => conv_std_logic_vector(76, 8),
27068 => conv_std_logic_vector(77, 8),
27069 => conv_std_logic_vector(77, 8),
27070 => conv_std_logic_vector(77, 8),
27071 => conv_std_logic_vector(78, 8),
27072 => conv_std_logic_vector(78, 8),
27073 => conv_std_logic_vector(79, 8),
27074 => conv_std_logic_vector(79, 8),
27075 => conv_std_logic_vector(79, 8),
27076 => conv_std_logic_vector(80, 8),
27077 => conv_std_logic_vector(80, 8),
27078 => conv_std_logic_vector(81, 8),
27079 => conv_std_logic_vector(81, 8),
27080 => conv_std_logic_vector(82, 8),
27081 => conv_std_logic_vector(82, 8),
27082 => conv_std_logic_vector(82, 8),
27083 => conv_std_logic_vector(83, 8),
27084 => conv_std_logic_vector(83, 8),
27085 => conv_std_logic_vector(84, 8),
27086 => conv_std_logic_vector(84, 8),
27087 => conv_std_logic_vector(84, 8),
27088 => conv_std_logic_vector(85, 8),
27089 => conv_std_logic_vector(85, 8),
27090 => conv_std_logic_vector(86, 8),
27091 => conv_std_logic_vector(86, 8),
27092 => conv_std_logic_vector(86, 8),
27093 => conv_std_logic_vector(87, 8),
27094 => conv_std_logic_vector(87, 8),
27095 => conv_std_logic_vector(88, 8),
27096 => conv_std_logic_vector(88, 8),
27097 => conv_std_logic_vector(89, 8),
27098 => conv_std_logic_vector(89, 8),
27099 => conv_std_logic_vector(89, 8),
27100 => conv_std_logic_vector(90, 8),
27101 => conv_std_logic_vector(90, 8),
27102 => conv_std_logic_vector(91, 8),
27103 => conv_std_logic_vector(91, 8),
27104 => conv_std_logic_vector(91, 8),
27105 => conv_std_logic_vector(92, 8),
27106 => conv_std_logic_vector(92, 8),
27107 => conv_std_logic_vector(93, 8),
27108 => conv_std_logic_vector(93, 8),
27109 => conv_std_logic_vector(93, 8),
27110 => conv_std_logic_vector(94, 8),
27111 => conv_std_logic_vector(94, 8),
27112 => conv_std_logic_vector(95, 8),
27113 => conv_std_logic_vector(95, 8),
27114 => conv_std_logic_vector(95, 8),
27115 => conv_std_logic_vector(96, 8),
27116 => conv_std_logic_vector(96, 8),
27117 => conv_std_logic_vector(97, 8),
27118 => conv_std_logic_vector(97, 8),
27119 => conv_std_logic_vector(98, 8),
27120 => conv_std_logic_vector(98, 8),
27121 => conv_std_logic_vector(98, 8),
27122 => conv_std_logic_vector(99, 8),
27123 => conv_std_logic_vector(99, 8),
27124 => conv_std_logic_vector(100, 8),
27125 => conv_std_logic_vector(100, 8),
27126 => conv_std_logic_vector(100, 8),
27127 => conv_std_logic_vector(101, 8),
27128 => conv_std_logic_vector(101, 8),
27129 => conv_std_logic_vector(102, 8),
27130 => conv_std_logic_vector(102, 8),
27131 => conv_std_logic_vector(102, 8),
27132 => conv_std_logic_vector(103, 8),
27133 => conv_std_logic_vector(103, 8),
27134 => conv_std_logic_vector(104, 8),
27135 => conv_std_logic_vector(104, 8),
27136 => conv_std_logic_vector(0, 8),
27137 => conv_std_logic_vector(0, 8),
27138 => conv_std_logic_vector(0, 8),
27139 => conv_std_logic_vector(1, 8),
27140 => conv_std_logic_vector(1, 8),
27141 => conv_std_logic_vector(2, 8),
27142 => conv_std_logic_vector(2, 8),
27143 => conv_std_logic_vector(2, 8),
27144 => conv_std_logic_vector(3, 8),
27145 => conv_std_logic_vector(3, 8),
27146 => conv_std_logic_vector(4, 8),
27147 => conv_std_logic_vector(4, 8),
27148 => conv_std_logic_vector(4, 8),
27149 => conv_std_logic_vector(5, 8),
27150 => conv_std_logic_vector(5, 8),
27151 => conv_std_logic_vector(6, 8),
27152 => conv_std_logic_vector(6, 8),
27153 => conv_std_logic_vector(7, 8),
27154 => conv_std_logic_vector(7, 8),
27155 => conv_std_logic_vector(7, 8),
27156 => conv_std_logic_vector(8, 8),
27157 => conv_std_logic_vector(8, 8),
27158 => conv_std_logic_vector(9, 8),
27159 => conv_std_logic_vector(9, 8),
27160 => conv_std_logic_vector(9, 8),
27161 => conv_std_logic_vector(10, 8),
27162 => conv_std_logic_vector(10, 8),
27163 => conv_std_logic_vector(11, 8),
27164 => conv_std_logic_vector(11, 8),
27165 => conv_std_logic_vector(12, 8),
27166 => conv_std_logic_vector(12, 8),
27167 => conv_std_logic_vector(12, 8),
27168 => conv_std_logic_vector(13, 8),
27169 => conv_std_logic_vector(13, 8),
27170 => conv_std_logic_vector(14, 8),
27171 => conv_std_logic_vector(14, 8),
27172 => conv_std_logic_vector(14, 8),
27173 => conv_std_logic_vector(15, 8),
27174 => conv_std_logic_vector(15, 8),
27175 => conv_std_logic_vector(16, 8),
27176 => conv_std_logic_vector(16, 8),
27177 => conv_std_logic_vector(16, 8),
27178 => conv_std_logic_vector(17, 8),
27179 => conv_std_logic_vector(17, 8),
27180 => conv_std_logic_vector(18, 8),
27181 => conv_std_logic_vector(18, 8),
27182 => conv_std_logic_vector(19, 8),
27183 => conv_std_logic_vector(19, 8),
27184 => conv_std_logic_vector(19, 8),
27185 => conv_std_logic_vector(20, 8),
27186 => conv_std_logic_vector(20, 8),
27187 => conv_std_logic_vector(21, 8),
27188 => conv_std_logic_vector(21, 8),
27189 => conv_std_logic_vector(21, 8),
27190 => conv_std_logic_vector(22, 8),
27191 => conv_std_logic_vector(22, 8),
27192 => conv_std_logic_vector(23, 8),
27193 => conv_std_logic_vector(23, 8),
27194 => conv_std_logic_vector(24, 8),
27195 => conv_std_logic_vector(24, 8),
27196 => conv_std_logic_vector(24, 8),
27197 => conv_std_logic_vector(25, 8),
27198 => conv_std_logic_vector(25, 8),
27199 => conv_std_logic_vector(26, 8),
27200 => conv_std_logic_vector(26, 8),
27201 => conv_std_logic_vector(26, 8),
27202 => conv_std_logic_vector(27, 8),
27203 => conv_std_logic_vector(27, 8),
27204 => conv_std_logic_vector(28, 8),
27205 => conv_std_logic_vector(28, 8),
27206 => conv_std_logic_vector(28, 8),
27207 => conv_std_logic_vector(29, 8),
27208 => conv_std_logic_vector(29, 8),
27209 => conv_std_logic_vector(30, 8),
27210 => conv_std_logic_vector(30, 8),
27211 => conv_std_logic_vector(31, 8),
27212 => conv_std_logic_vector(31, 8),
27213 => conv_std_logic_vector(31, 8),
27214 => conv_std_logic_vector(32, 8),
27215 => conv_std_logic_vector(32, 8),
27216 => conv_std_logic_vector(33, 8),
27217 => conv_std_logic_vector(33, 8),
27218 => conv_std_logic_vector(33, 8),
27219 => conv_std_logic_vector(34, 8),
27220 => conv_std_logic_vector(34, 8),
27221 => conv_std_logic_vector(35, 8),
27222 => conv_std_logic_vector(35, 8),
27223 => conv_std_logic_vector(36, 8),
27224 => conv_std_logic_vector(36, 8),
27225 => conv_std_logic_vector(36, 8),
27226 => conv_std_logic_vector(37, 8),
27227 => conv_std_logic_vector(37, 8),
27228 => conv_std_logic_vector(38, 8),
27229 => conv_std_logic_vector(38, 8),
27230 => conv_std_logic_vector(38, 8),
27231 => conv_std_logic_vector(39, 8),
27232 => conv_std_logic_vector(39, 8),
27233 => conv_std_logic_vector(40, 8),
27234 => conv_std_logic_vector(40, 8),
27235 => conv_std_logic_vector(40, 8),
27236 => conv_std_logic_vector(41, 8),
27237 => conv_std_logic_vector(41, 8),
27238 => conv_std_logic_vector(42, 8),
27239 => conv_std_logic_vector(42, 8),
27240 => conv_std_logic_vector(43, 8),
27241 => conv_std_logic_vector(43, 8),
27242 => conv_std_logic_vector(43, 8),
27243 => conv_std_logic_vector(44, 8),
27244 => conv_std_logic_vector(44, 8),
27245 => conv_std_logic_vector(45, 8),
27246 => conv_std_logic_vector(45, 8),
27247 => conv_std_logic_vector(45, 8),
27248 => conv_std_logic_vector(46, 8),
27249 => conv_std_logic_vector(46, 8),
27250 => conv_std_logic_vector(47, 8),
27251 => conv_std_logic_vector(47, 8),
27252 => conv_std_logic_vector(48, 8),
27253 => conv_std_logic_vector(48, 8),
27254 => conv_std_logic_vector(48, 8),
27255 => conv_std_logic_vector(49, 8),
27256 => conv_std_logic_vector(49, 8),
27257 => conv_std_logic_vector(50, 8),
27258 => conv_std_logic_vector(50, 8),
27259 => conv_std_logic_vector(50, 8),
27260 => conv_std_logic_vector(51, 8),
27261 => conv_std_logic_vector(51, 8),
27262 => conv_std_logic_vector(52, 8),
27263 => conv_std_logic_vector(52, 8),
27264 => conv_std_logic_vector(53, 8),
27265 => conv_std_logic_vector(53, 8),
27266 => conv_std_logic_vector(53, 8),
27267 => conv_std_logic_vector(54, 8),
27268 => conv_std_logic_vector(54, 8),
27269 => conv_std_logic_vector(55, 8),
27270 => conv_std_logic_vector(55, 8),
27271 => conv_std_logic_vector(55, 8),
27272 => conv_std_logic_vector(56, 8),
27273 => conv_std_logic_vector(56, 8),
27274 => conv_std_logic_vector(57, 8),
27275 => conv_std_logic_vector(57, 8),
27276 => conv_std_logic_vector(57, 8),
27277 => conv_std_logic_vector(58, 8),
27278 => conv_std_logic_vector(58, 8),
27279 => conv_std_logic_vector(59, 8),
27280 => conv_std_logic_vector(59, 8),
27281 => conv_std_logic_vector(60, 8),
27282 => conv_std_logic_vector(60, 8),
27283 => conv_std_logic_vector(60, 8),
27284 => conv_std_logic_vector(61, 8),
27285 => conv_std_logic_vector(61, 8),
27286 => conv_std_logic_vector(62, 8),
27287 => conv_std_logic_vector(62, 8),
27288 => conv_std_logic_vector(62, 8),
27289 => conv_std_logic_vector(63, 8),
27290 => conv_std_logic_vector(63, 8),
27291 => conv_std_logic_vector(64, 8),
27292 => conv_std_logic_vector(64, 8),
27293 => conv_std_logic_vector(65, 8),
27294 => conv_std_logic_vector(65, 8),
27295 => conv_std_logic_vector(65, 8),
27296 => conv_std_logic_vector(66, 8),
27297 => conv_std_logic_vector(66, 8),
27298 => conv_std_logic_vector(67, 8),
27299 => conv_std_logic_vector(67, 8),
27300 => conv_std_logic_vector(67, 8),
27301 => conv_std_logic_vector(68, 8),
27302 => conv_std_logic_vector(68, 8),
27303 => conv_std_logic_vector(69, 8),
27304 => conv_std_logic_vector(69, 8),
27305 => conv_std_logic_vector(69, 8),
27306 => conv_std_logic_vector(70, 8),
27307 => conv_std_logic_vector(70, 8),
27308 => conv_std_logic_vector(71, 8),
27309 => conv_std_logic_vector(71, 8),
27310 => conv_std_logic_vector(72, 8),
27311 => conv_std_logic_vector(72, 8),
27312 => conv_std_logic_vector(72, 8),
27313 => conv_std_logic_vector(73, 8),
27314 => conv_std_logic_vector(73, 8),
27315 => conv_std_logic_vector(74, 8),
27316 => conv_std_logic_vector(74, 8),
27317 => conv_std_logic_vector(74, 8),
27318 => conv_std_logic_vector(75, 8),
27319 => conv_std_logic_vector(75, 8),
27320 => conv_std_logic_vector(76, 8),
27321 => conv_std_logic_vector(76, 8),
27322 => conv_std_logic_vector(77, 8),
27323 => conv_std_logic_vector(77, 8),
27324 => conv_std_logic_vector(77, 8),
27325 => conv_std_logic_vector(78, 8),
27326 => conv_std_logic_vector(78, 8),
27327 => conv_std_logic_vector(79, 8),
27328 => conv_std_logic_vector(79, 8),
27329 => conv_std_logic_vector(79, 8),
27330 => conv_std_logic_vector(80, 8),
27331 => conv_std_logic_vector(80, 8),
27332 => conv_std_logic_vector(81, 8),
27333 => conv_std_logic_vector(81, 8),
27334 => conv_std_logic_vector(81, 8),
27335 => conv_std_logic_vector(82, 8),
27336 => conv_std_logic_vector(82, 8),
27337 => conv_std_logic_vector(83, 8),
27338 => conv_std_logic_vector(83, 8),
27339 => conv_std_logic_vector(84, 8),
27340 => conv_std_logic_vector(84, 8),
27341 => conv_std_logic_vector(84, 8),
27342 => conv_std_logic_vector(85, 8),
27343 => conv_std_logic_vector(85, 8),
27344 => conv_std_logic_vector(86, 8),
27345 => conv_std_logic_vector(86, 8),
27346 => conv_std_logic_vector(86, 8),
27347 => conv_std_logic_vector(87, 8),
27348 => conv_std_logic_vector(87, 8),
27349 => conv_std_logic_vector(88, 8),
27350 => conv_std_logic_vector(88, 8),
27351 => conv_std_logic_vector(89, 8),
27352 => conv_std_logic_vector(89, 8),
27353 => conv_std_logic_vector(89, 8),
27354 => conv_std_logic_vector(90, 8),
27355 => conv_std_logic_vector(90, 8),
27356 => conv_std_logic_vector(91, 8),
27357 => conv_std_logic_vector(91, 8),
27358 => conv_std_logic_vector(91, 8),
27359 => conv_std_logic_vector(92, 8),
27360 => conv_std_logic_vector(92, 8),
27361 => conv_std_logic_vector(93, 8),
27362 => conv_std_logic_vector(93, 8),
27363 => conv_std_logic_vector(93, 8),
27364 => conv_std_logic_vector(94, 8),
27365 => conv_std_logic_vector(94, 8),
27366 => conv_std_logic_vector(95, 8),
27367 => conv_std_logic_vector(95, 8),
27368 => conv_std_logic_vector(96, 8),
27369 => conv_std_logic_vector(96, 8),
27370 => conv_std_logic_vector(96, 8),
27371 => conv_std_logic_vector(97, 8),
27372 => conv_std_logic_vector(97, 8),
27373 => conv_std_logic_vector(98, 8),
27374 => conv_std_logic_vector(98, 8),
27375 => conv_std_logic_vector(98, 8),
27376 => conv_std_logic_vector(99, 8),
27377 => conv_std_logic_vector(99, 8),
27378 => conv_std_logic_vector(100, 8),
27379 => conv_std_logic_vector(100, 8),
27380 => conv_std_logic_vector(101, 8),
27381 => conv_std_logic_vector(101, 8),
27382 => conv_std_logic_vector(101, 8),
27383 => conv_std_logic_vector(102, 8),
27384 => conv_std_logic_vector(102, 8),
27385 => conv_std_logic_vector(103, 8),
27386 => conv_std_logic_vector(103, 8),
27387 => conv_std_logic_vector(103, 8),
27388 => conv_std_logic_vector(104, 8),
27389 => conv_std_logic_vector(104, 8),
27390 => conv_std_logic_vector(105, 8),
27391 => conv_std_logic_vector(105, 8),
27392 => conv_std_logic_vector(0, 8),
27393 => conv_std_logic_vector(0, 8),
27394 => conv_std_logic_vector(0, 8),
27395 => conv_std_logic_vector(1, 8),
27396 => conv_std_logic_vector(1, 8),
27397 => conv_std_logic_vector(2, 8),
27398 => conv_std_logic_vector(2, 8),
27399 => conv_std_logic_vector(2, 8),
27400 => conv_std_logic_vector(3, 8),
27401 => conv_std_logic_vector(3, 8),
27402 => conv_std_logic_vector(4, 8),
27403 => conv_std_logic_vector(4, 8),
27404 => conv_std_logic_vector(5, 8),
27405 => conv_std_logic_vector(5, 8),
27406 => conv_std_logic_vector(5, 8),
27407 => conv_std_logic_vector(6, 8),
27408 => conv_std_logic_vector(6, 8),
27409 => conv_std_logic_vector(7, 8),
27410 => conv_std_logic_vector(7, 8),
27411 => conv_std_logic_vector(7, 8),
27412 => conv_std_logic_vector(8, 8),
27413 => conv_std_logic_vector(8, 8),
27414 => conv_std_logic_vector(9, 8),
27415 => conv_std_logic_vector(9, 8),
27416 => conv_std_logic_vector(10, 8),
27417 => conv_std_logic_vector(10, 8),
27418 => conv_std_logic_vector(10, 8),
27419 => conv_std_logic_vector(11, 8),
27420 => conv_std_logic_vector(11, 8),
27421 => conv_std_logic_vector(12, 8),
27422 => conv_std_logic_vector(12, 8),
27423 => conv_std_logic_vector(12, 8),
27424 => conv_std_logic_vector(13, 8),
27425 => conv_std_logic_vector(13, 8),
27426 => conv_std_logic_vector(14, 8),
27427 => conv_std_logic_vector(14, 8),
27428 => conv_std_logic_vector(15, 8),
27429 => conv_std_logic_vector(15, 8),
27430 => conv_std_logic_vector(15, 8),
27431 => conv_std_logic_vector(16, 8),
27432 => conv_std_logic_vector(16, 8),
27433 => conv_std_logic_vector(17, 8),
27434 => conv_std_logic_vector(17, 8),
27435 => conv_std_logic_vector(17, 8),
27436 => conv_std_logic_vector(18, 8),
27437 => conv_std_logic_vector(18, 8),
27438 => conv_std_logic_vector(19, 8),
27439 => conv_std_logic_vector(19, 8),
27440 => conv_std_logic_vector(20, 8),
27441 => conv_std_logic_vector(20, 8),
27442 => conv_std_logic_vector(20, 8),
27443 => conv_std_logic_vector(21, 8),
27444 => conv_std_logic_vector(21, 8),
27445 => conv_std_logic_vector(22, 8),
27446 => conv_std_logic_vector(22, 8),
27447 => conv_std_logic_vector(22, 8),
27448 => conv_std_logic_vector(23, 8),
27449 => conv_std_logic_vector(23, 8),
27450 => conv_std_logic_vector(24, 8),
27451 => conv_std_logic_vector(24, 8),
27452 => conv_std_logic_vector(25, 8),
27453 => conv_std_logic_vector(25, 8),
27454 => conv_std_logic_vector(25, 8),
27455 => conv_std_logic_vector(26, 8),
27456 => conv_std_logic_vector(26, 8),
27457 => conv_std_logic_vector(27, 8),
27458 => conv_std_logic_vector(27, 8),
27459 => conv_std_logic_vector(28, 8),
27460 => conv_std_logic_vector(28, 8),
27461 => conv_std_logic_vector(28, 8),
27462 => conv_std_logic_vector(29, 8),
27463 => conv_std_logic_vector(29, 8),
27464 => conv_std_logic_vector(30, 8),
27465 => conv_std_logic_vector(30, 8),
27466 => conv_std_logic_vector(30, 8),
27467 => conv_std_logic_vector(31, 8),
27468 => conv_std_logic_vector(31, 8),
27469 => conv_std_logic_vector(32, 8),
27470 => conv_std_logic_vector(32, 8),
27471 => conv_std_logic_vector(33, 8),
27472 => conv_std_logic_vector(33, 8),
27473 => conv_std_logic_vector(33, 8),
27474 => conv_std_logic_vector(34, 8),
27475 => conv_std_logic_vector(34, 8),
27476 => conv_std_logic_vector(35, 8),
27477 => conv_std_logic_vector(35, 8),
27478 => conv_std_logic_vector(35, 8),
27479 => conv_std_logic_vector(36, 8),
27480 => conv_std_logic_vector(36, 8),
27481 => conv_std_logic_vector(37, 8),
27482 => conv_std_logic_vector(37, 8),
27483 => conv_std_logic_vector(38, 8),
27484 => conv_std_logic_vector(38, 8),
27485 => conv_std_logic_vector(38, 8),
27486 => conv_std_logic_vector(39, 8),
27487 => conv_std_logic_vector(39, 8),
27488 => conv_std_logic_vector(40, 8),
27489 => conv_std_logic_vector(40, 8),
27490 => conv_std_logic_vector(40, 8),
27491 => conv_std_logic_vector(41, 8),
27492 => conv_std_logic_vector(41, 8),
27493 => conv_std_logic_vector(42, 8),
27494 => conv_std_logic_vector(42, 8),
27495 => conv_std_logic_vector(43, 8),
27496 => conv_std_logic_vector(43, 8),
27497 => conv_std_logic_vector(43, 8),
27498 => conv_std_logic_vector(44, 8),
27499 => conv_std_logic_vector(44, 8),
27500 => conv_std_logic_vector(45, 8),
27501 => conv_std_logic_vector(45, 8),
27502 => conv_std_logic_vector(45, 8),
27503 => conv_std_logic_vector(46, 8),
27504 => conv_std_logic_vector(46, 8),
27505 => conv_std_logic_vector(47, 8),
27506 => conv_std_logic_vector(47, 8),
27507 => conv_std_logic_vector(48, 8),
27508 => conv_std_logic_vector(48, 8),
27509 => conv_std_logic_vector(48, 8),
27510 => conv_std_logic_vector(49, 8),
27511 => conv_std_logic_vector(49, 8),
27512 => conv_std_logic_vector(50, 8),
27513 => conv_std_logic_vector(50, 8),
27514 => conv_std_logic_vector(50, 8),
27515 => conv_std_logic_vector(51, 8),
27516 => conv_std_logic_vector(51, 8),
27517 => conv_std_logic_vector(52, 8),
27518 => conv_std_logic_vector(52, 8),
27519 => conv_std_logic_vector(53, 8),
27520 => conv_std_logic_vector(53, 8),
27521 => conv_std_logic_vector(53, 8),
27522 => conv_std_logic_vector(54, 8),
27523 => conv_std_logic_vector(54, 8),
27524 => conv_std_logic_vector(55, 8),
27525 => conv_std_logic_vector(55, 8),
27526 => conv_std_logic_vector(56, 8),
27527 => conv_std_logic_vector(56, 8),
27528 => conv_std_logic_vector(56, 8),
27529 => conv_std_logic_vector(57, 8),
27530 => conv_std_logic_vector(57, 8),
27531 => conv_std_logic_vector(58, 8),
27532 => conv_std_logic_vector(58, 8),
27533 => conv_std_logic_vector(58, 8),
27534 => conv_std_logic_vector(59, 8),
27535 => conv_std_logic_vector(59, 8),
27536 => conv_std_logic_vector(60, 8),
27537 => conv_std_logic_vector(60, 8),
27538 => conv_std_logic_vector(61, 8),
27539 => conv_std_logic_vector(61, 8),
27540 => conv_std_logic_vector(61, 8),
27541 => conv_std_logic_vector(62, 8),
27542 => conv_std_logic_vector(62, 8),
27543 => conv_std_logic_vector(63, 8),
27544 => conv_std_logic_vector(63, 8),
27545 => conv_std_logic_vector(63, 8),
27546 => conv_std_logic_vector(64, 8),
27547 => conv_std_logic_vector(64, 8),
27548 => conv_std_logic_vector(65, 8),
27549 => conv_std_logic_vector(65, 8),
27550 => conv_std_logic_vector(66, 8),
27551 => conv_std_logic_vector(66, 8),
27552 => conv_std_logic_vector(66, 8),
27553 => conv_std_logic_vector(67, 8),
27554 => conv_std_logic_vector(67, 8),
27555 => conv_std_logic_vector(68, 8),
27556 => conv_std_logic_vector(68, 8),
27557 => conv_std_logic_vector(68, 8),
27558 => conv_std_logic_vector(69, 8),
27559 => conv_std_logic_vector(69, 8),
27560 => conv_std_logic_vector(70, 8),
27561 => conv_std_logic_vector(70, 8),
27562 => conv_std_logic_vector(71, 8),
27563 => conv_std_logic_vector(71, 8),
27564 => conv_std_logic_vector(71, 8),
27565 => conv_std_logic_vector(72, 8),
27566 => conv_std_logic_vector(72, 8),
27567 => conv_std_logic_vector(73, 8),
27568 => conv_std_logic_vector(73, 8),
27569 => conv_std_logic_vector(73, 8),
27570 => conv_std_logic_vector(74, 8),
27571 => conv_std_logic_vector(74, 8),
27572 => conv_std_logic_vector(75, 8),
27573 => conv_std_logic_vector(75, 8),
27574 => conv_std_logic_vector(76, 8),
27575 => conv_std_logic_vector(76, 8),
27576 => conv_std_logic_vector(76, 8),
27577 => conv_std_logic_vector(77, 8),
27578 => conv_std_logic_vector(77, 8),
27579 => conv_std_logic_vector(78, 8),
27580 => conv_std_logic_vector(78, 8),
27581 => conv_std_logic_vector(78, 8),
27582 => conv_std_logic_vector(79, 8),
27583 => conv_std_logic_vector(79, 8),
27584 => conv_std_logic_vector(80, 8),
27585 => conv_std_logic_vector(80, 8),
27586 => conv_std_logic_vector(81, 8),
27587 => conv_std_logic_vector(81, 8),
27588 => conv_std_logic_vector(81, 8),
27589 => conv_std_logic_vector(82, 8),
27590 => conv_std_logic_vector(82, 8),
27591 => conv_std_logic_vector(83, 8),
27592 => conv_std_logic_vector(83, 8),
27593 => conv_std_logic_vector(84, 8),
27594 => conv_std_logic_vector(84, 8),
27595 => conv_std_logic_vector(84, 8),
27596 => conv_std_logic_vector(85, 8),
27597 => conv_std_logic_vector(85, 8),
27598 => conv_std_logic_vector(86, 8),
27599 => conv_std_logic_vector(86, 8),
27600 => conv_std_logic_vector(86, 8),
27601 => conv_std_logic_vector(87, 8),
27602 => conv_std_logic_vector(87, 8),
27603 => conv_std_logic_vector(88, 8),
27604 => conv_std_logic_vector(88, 8),
27605 => conv_std_logic_vector(89, 8),
27606 => conv_std_logic_vector(89, 8),
27607 => conv_std_logic_vector(89, 8),
27608 => conv_std_logic_vector(90, 8),
27609 => conv_std_logic_vector(90, 8),
27610 => conv_std_logic_vector(91, 8),
27611 => conv_std_logic_vector(91, 8),
27612 => conv_std_logic_vector(91, 8),
27613 => conv_std_logic_vector(92, 8),
27614 => conv_std_logic_vector(92, 8),
27615 => conv_std_logic_vector(93, 8),
27616 => conv_std_logic_vector(93, 8),
27617 => conv_std_logic_vector(94, 8),
27618 => conv_std_logic_vector(94, 8),
27619 => conv_std_logic_vector(94, 8),
27620 => conv_std_logic_vector(95, 8),
27621 => conv_std_logic_vector(95, 8),
27622 => conv_std_logic_vector(96, 8),
27623 => conv_std_logic_vector(96, 8),
27624 => conv_std_logic_vector(96, 8),
27625 => conv_std_logic_vector(97, 8),
27626 => conv_std_logic_vector(97, 8),
27627 => conv_std_logic_vector(98, 8),
27628 => conv_std_logic_vector(98, 8),
27629 => conv_std_logic_vector(99, 8),
27630 => conv_std_logic_vector(99, 8),
27631 => conv_std_logic_vector(99, 8),
27632 => conv_std_logic_vector(100, 8),
27633 => conv_std_logic_vector(100, 8),
27634 => conv_std_logic_vector(101, 8),
27635 => conv_std_logic_vector(101, 8),
27636 => conv_std_logic_vector(101, 8),
27637 => conv_std_logic_vector(102, 8),
27638 => conv_std_logic_vector(102, 8),
27639 => conv_std_logic_vector(103, 8),
27640 => conv_std_logic_vector(103, 8),
27641 => conv_std_logic_vector(104, 8),
27642 => conv_std_logic_vector(104, 8),
27643 => conv_std_logic_vector(104, 8),
27644 => conv_std_logic_vector(105, 8),
27645 => conv_std_logic_vector(105, 8),
27646 => conv_std_logic_vector(106, 8),
27647 => conv_std_logic_vector(106, 8),
27648 => conv_std_logic_vector(0, 8),
27649 => conv_std_logic_vector(0, 8),
27650 => conv_std_logic_vector(0, 8),
27651 => conv_std_logic_vector(1, 8),
27652 => conv_std_logic_vector(1, 8),
27653 => conv_std_logic_vector(2, 8),
27654 => conv_std_logic_vector(2, 8),
27655 => conv_std_logic_vector(2, 8),
27656 => conv_std_logic_vector(3, 8),
27657 => conv_std_logic_vector(3, 8),
27658 => conv_std_logic_vector(4, 8),
27659 => conv_std_logic_vector(4, 8),
27660 => conv_std_logic_vector(5, 8),
27661 => conv_std_logic_vector(5, 8),
27662 => conv_std_logic_vector(5, 8),
27663 => conv_std_logic_vector(6, 8),
27664 => conv_std_logic_vector(6, 8),
27665 => conv_std_logic_vector(7, 8),
27666 => conv_std_logic_vector(7, 8),
27667 => conv_std_logic_vector(8, 8),
27668 => conv_std_logic_vector(8, 8),
27669 => conv_std_logic_vector(8, 8),
27670 => conv_std_logic_vector(9, 8),
27671 => conv_std_logic_vector(9, 8),
27672 => conv_std_logic_vector(10, 8),
27673 => conv_std_logic_vector(10, 8),
27674 => conv_std_logic_vector(10, 8),
27675 => conv_std_logic_vector(11, 8),
27676 => conv_std_logic_vector(11, 8),
27677 => conv_std_logic_vector(12, 8),
27678 => conv_std_logic_vector(12, 8),
27679 => conv_std_logic_vector(13, 8),
27680 => conv_std_logic_vector(13, 8),
27681 => conv_std_logic_vector(13, 8),
27682 => conv_std_logic_vector(14, 8),
27683 => conv_std_logic_vector(14, 8),
27684 => conv_std_logic_vector(15, 8),
27685 => conv_std_logic_vector(15, 8),
27686 => conv_std_logic_vector(16, 8),
27687 => conv_std_logic_vector(16, 8),
27688 => conv_std_logic_vector(16, 8),
27689 => conv_std_logic_vector(17, 8),
27690 => conv_std_logic_vector(17, 8),
27691 => conv_std_logic_vector(18, 8),
27692 => conv_std_logic_vector(18, 8),
27693 => conv_std_logic_vector(18, 8),
27694 => conv_std_logic_vector(19, 8),
27695 => conv_std_logic_vector(19, 8),
27696 => conv_std_logic_vector(20, 8),
27697 => conv_std_logic_vector(20, 8),
27698 => conv_std_logic_vector(21, 8),
27699 => conv_std_logic_vector(21, 8),
27700 => conv_std_logic_vector(21, 8),
27701 => conv_std_logic_vector(22, 8),
27702 => conv_std_logic_vector(22, 8),
27703 => conv_std_logic_vector(23, 8),
27704 => conv_std_logic_vector(23, 8),
27705 => conv_std_logic_vector(24, 8),
27706 => conv_std_logic_vector(24, 8),
27707 => conv_std_logic_vector(24, 8),
27708 => conv_std_logic_vector(25, 8),
27709 => conv_std_logic_vector(25, 8),
27710 => conv_std_logic_vector(26, 8),
27711 => conv_std_logic_vector(26, 8),
27712 => conv_std_logic_vector(27, 8),
27713 => conv_std_logic_vector(27, 8),
27714 => conv_std_logic_vector(27, 8),
27715 => conv_std_logic_vector(28, 8),
27716 => conv_std_logic_vector(28, 8),
27717 => conv_std_logic_vector(29, 8),
27718 => conv_std_logic_vector(29, 8),
27719 => conv_std_logic_vector(29, 8),
27720 => conv_std_logic_vector(30, 8),
27721 => conv_std_logic_vector(30, 8),
27722 => conv_std_logic_vector(31, 8),
27723 => conv_std_logic_vector(31, 8),
27724 => conv_std_logic_vector(32, 8),
27725 => conv_std_logic_vector(32, 8),
27726 => conv_std_logic_vector(32, 8),
27727 => conv_std_logic_vector(33, 8),
27728 => conv_std_logic_vector(33, 8),
27729 => conv_std_logic_vector(34, 8),
27730 => conv_std_logic_vector(34, 8),
27731 => conv_std_logic_vector(35, 8),
27732 => conv_std_logic_vector(35, 8),
27733 => conv_std_logic_vector(35, 8),
27734 => conv_std_logic_vector(36, 8),
27735 => conv_std_logic_vector(36, 8),
27736 => conv_std_logic_vector(37, 8),
27737 => conv_std_logic_vector(37, 8),
27738 => conv_std_logic_vector(37, 8),
27739 => conv_std_logic_vector(38, 8),
27740 => conv_std_logic_vector(38, 8),
27741 => conv_std_logic_vector(39, 8),
27742 => conv_std_logic_vector(39, 8),
27743 => conv_std_logic_vector(40, 8),
27744 => conv_std_logic_vector(40, 8),
27745 => conv_std_logic_vector(40, 8),
27746 => conv_std_logic_vector(41, 8),
27747 => conv_std_logic_vector(41, 8),
27748 => conv_std_logic_vector(42, 8),
27749 => conv_std_logic_vector(42, 8),
27750 => conv_std_logic_vector(43, 8),
27751 => conv_std_logic_vector(43, 8),
27752 => conv_std_logic_vector(43, 8),
27753 => conv_std_logic_vector(44, 8),
27754 => conv_std_logic_vector(44, 8),
27755 => conv_std_logic_vector(45, 8),
27756 => conv_std_logic_vector(45, 8),
27757 => conv_std_logic_vector(45, 8),
27758 => conv_std_logic_vector(46, 8),
27759 => conv_std_logic_vector(46, 8),
27760 => conv_std_logic_vector(47, 8),
27761 => conv_std_logic_vector(47, 8),
27762 => conv_std_logic_vector(48, 8),
27763 => conv_std_logic_vector(48, 8),
27764 => conv_std_logic_vector(48, 8),
27765 => conv_std_logic_vector(49, 8),
27766 => conv_std_logic_vector(49, 8),
27767 => conv_std_logic_vector(50, 8),
27768 => conv_std_logic_vector(50, 8),
27769 => conv_std_logic_vector(51, 8),
27770 => conv_std_logic_vector(51, 8),
27771 => conv_std_logic_vector(51, 8),
27772 => conv_std_logic_vector(52, 8),
27773 => conv_std_logic_vector(52, 8),
27774 => conv_std_logic_vector(53, 8),
27775 => conv_std_logic_vector(53, 8),
27776 => conv_std_logic_vector(54, 8),
27777 => conv_std_logic_vector(54, 8),
27778 => conv_std_logic_vector(54, 8),
27779 => conv_std_logic_vector(55, 8),
27780 => conv_std_logic_vector(55, 8),
27781 => conv_std_logic_vector(56, 8),
27782 => conv_std_logic_vector(56, 8),
27783 => conv_std_logic_vector(56, 8),
27784 => conv_std_logic_vector(57, 8),
27785 => conv_std_logic_vector(57, 8),
27786 => conv_std_logic_vector(58, 8),
27787 => conv_std_logic_vector(58, 8),
27788 => conv_std_logic_vector(59, 8),
27789 => conv_std_logic_vector(59, 8),
27790 => conv_std_logic_vector(59, 8),
27791 => conv_std_logic_vector(60, 8),
27792 => conv_std_logic_vector(60, 8),
27793 => conv_std_logic_vector(61, 8),
27794 => conv_std_logic_vector(61, 8),
27795 => conv_std_logic_vector(62, 8),
27796 => conv_std_logic_vector(62, 8),
27797 => conv_std_logic_vector(62, 8),
27798 => conv_std_logic_vector(63, 8),
27799 => conv_std_logic_vector(63, 8),
27800 => conv_std_logic_vector(64, 8),
27801 => conv_std_logic_vector(64, 8),
27802 => conv_std_logic_vector(64, 8),
27803 => conv_std_logic_vector(65, 8),
27804 => conv_std_logic_vector(65, 8),
27805 => conv_std_logic_vector(66, 8),
27806 => conv_std_logic_vector(66, 8),
27807 => conv_std_logic_vector(67, 8),
27808 => conv_std_logic_vector(67, 8),
27809 => conv_std_logic_vector(67, 8),
27810 => conv_std_logic_vector(68, 8),
27811 => conv_std_logic_vector(68, 8),
27812 => conv_std_logic_vector(69, 8),
27813 => conv_std_logic_vector(69, 8),
27814 => conv_std_logic_vector(70, 8),
27815 => conv_std_logic_vector(70, 8),
27816 => conv_std_logic_vector(70, 8),
27817 => conv_std_logic_vector(71, 8),
27818 => conv_std_logic_vector(71, 8),
27819 => conv_std_logic_vector(72, 8),
27820 => conv_std_logic_vector(72, 8),
27821 => conv_std_logic_vector(72, 8),
27822 => conv_std_logic_vector(73, 8),
27823 => conv_std_logic_vector(73, 8),
27824 => conv_std_logic_vector(74, 8),
27825 => conv_std_logic_vector(74, 8),
27826 => conv_std_logic_vector(75, 8),
27827 => conv_std_logic_vector(75, 8),
27828 => conv_std_logic_vector(75, 8),
27829 => conv_std_logic_vector(76, 8),
27830 => conv_std_logic_vector(76, 8),
27831 => conv_std_logic_vector(77, 8),
27832 => conv_std_logic_vector(77, 8),
27833 => conv_std_logic_vector(78, 8),
27834 => conv_std_logic_vector(78, 8),
27835 => conv_std_logic_vector(78, 8),
27836 => conv_std_logic_vector(79, 8),
27837 => conv_std_logic_vector(79, 8),
27838 => conv_std_logic_vector(80, 8),
27839 => conv_std_logic_vector(80, 8),
27840 => conv_std_logic_vector(81, 8),
27841 => conv_std_logic_vector(81, 8),
27842 => conv_std_logic_vector(81, 8),
27843 => conv_std_logic_vector(82, 8),
27844 => conv_std_logic_vector(82, 8),
27845 => conv_std_logic_vector(83, 8),
27846 => conv_std_logic_vector(83, 8),
27847 => conv_std_logic_vector(83, 8),
27848 => conv_std_logic_vector(84, 8),
27849 => conv_std_logic_vector(84, 8),
27850 => conv_std_logic_vector(85, 8),
27851 => conv_std_logic_vector(85, 8),
27852 => conv_std_logic_vector(86, 8),
27853 => conv_std_logic_vector(86, 8),
27854 => conv_std_logic_vector(86, 8),
27855 => conv_std_logic_vector(87, 8),
27856 => conv_std_logic_vector(87, 8),
27857 => conv_std_logic_vector(88, 8),
27858 => conv_std_logic_vector(88, 8),
27859 => conv_std_logic_vector(89, 8),
27860 => conv_std_logic_vector(89, 8),
27861 => conv_std_logic_vector(89, 8),
27862 => conv_std_logic_vector(90, 8),
27863 => conv_std_logic_vector(90, 8),
27864 => conv_std_logic_vector(91, 8),
27865 => conv_std_logic_vector(91, 8),
27866 => conv_std_logic_vector(91, 8),
27867 => conv_std_logic_vector(92, 8),
27868 => conv_std_logic_vector(92, 8),
27869 => conv_std_logic_vector(93, 8),
27870 => conv_std_logic_vector(93, 8),
27871 => conv_std_logic_vector(94, 8),
27872 => conv_std_logic_vector(94, 8),
27873 => conv_std_logic_vector(94, 8),
27874 => conv_std_logic_vector(95, 8),
27875 => conv_std_logic_vector(95, 8),
27876 => conv_std_logic_vector(96, 8),
27877 => conv_std_logic_vector(96, 8),
27878 => conv_std_logic_vector(97, 8),
27879 => conv_std_logic_vector(97, 8),
27880 => conv_std_logic_vector(97, 8),
27881 => conv_std_logic_vector(98, 8),
27882 => conv_std_logic_vector(98, 8),
27883 => conv_std_logic_vector(99, 8),
27884 => conv_std_logic_vector(99, 8),
27885 => conv_std_logic_vector(99, 8),
27886 => conv_std_logic_vector(100, 8),
27887 => conv_std_logic_vector(100, 8),
27888 => conv_std_logic_vector(101, 8),
27889 => conv_std_logic_vector(101, 8),
27890 => conv_std_logic_vector(102, 8),
27891 => conv_std_logic_vector(102, 8),
27892 => conv_std_logic_vector(102, 8),
27893 => conv_std_logic_vector(103, 8),
27894 => conv_std_logic_vector(103, 8),
27895 => conv_std_logic_vector(104, 8),
27896 => conv_std_logic_vector(104, 8),
27897 => conv_std_logic_vector(105, 8),
27898 => conv_std_logic_vector(105, 8),
27899 => conv_std_logic_vector(105, 8),
27900 => conv_std_logic_vector(106, 8),
27901 => conv_std_logic_vector(106, 8),
27902 => conv_std_logic_vector(107, 8),
27903 => conv_std_logic_vector(107, 8),
27904 => conv_std_logic_vector(0, 8),
27905 => conv_std_logic_vector(0, 8),
27906 => conv_std_logic_vector(0, 8),
27907 => conv_std_logic_vector(1, 8),
27908 => conv_std_logic_vector(1, 8),
27909 => conv_std_logic_vector(2, 8),
27910 => conv_std_logic_vector(2, 8),
27911 => conv_std_logic_vector(2, 8),
27912 => conv_std_logic_vector(3, 8),
27913 => conv_std_logic_vector(3, 8),
27914 => conv_std_logic_vector(4, 8),
27915 => conv_std_logic_vector(4, 8),
27916 => conv_std_logic_vector(5, 8),
27917 => conv_std_logic_vector(5, 8),
27918 => conv_std_logic_vector(5, 8),
27919 => conv_std_logic_vector(6, 8),
27920 => conv_std_logic_vector(6, 8),
27921 => conv_std_logic_vector(7, 8),
27922 => conv_std_logic_vector(7, 8),
27923 => conv_std_logic_vector(8, 8),
27924 => conv_std_logic_vector(8, 8),
27925 => conv_std_logic_vector(8, 8),
27926 => conv_std_logic_vector(9, 8),
27927 => conv_std_logic_vector(9, 8),
27928 => conv_std_logic_vector(10, 8),
27929 => conv_std_logic_vector(10, 8),
27930 => conv_std_logic_vector(11, 8),
27931 => conv_std_logic_vector(11, 8),
27932 => conv_std_logic_vector(11, 8),
27933 => conv_std_logic_vector(12, 8),
27934 => conv_std_logic_vector(12, 8),
27935 => conv_std_logic_vector(13, 8),
27936 => conv_std_logic_vector(13, 8),
27937 => conv_std_logic_vector(14, 8),
27938 => conv_std_logic_vector(14, 8),
27939 => conv_std_logic_vector(14, 8),
27940 => conv_std_logic_vector(15, 8),
27941 => conv_std_logic_vector(15, 8),
27942 => conv_std_logic_vector(16, 8),
27943 => conv_std_logic_vector(16, 8),
27944 => conv_std_logic_vector(17, 8),
27945 => conv_std_logic_vector(17, 8),
27946 => conv_std_logic_vector(17, 8),
27947 => conv_std_logic_vector(18, 8),
27948 => conv_std_logic_vector(18, 8),
27949 => conv_std_logic_vector(19, 8),
27950 => conv_std_logic_vector(19, 8),
27951 => conv_std_logic_vector(20, 8),
27952 => conv_std_logic_vector(20, 8),
27953 => conv_std_logic_vector(20, 8),
27954 => conv_std_logic_vector(21, 8),
27955 => conv_std_logic_vector(21, 8),
27956 => conv_std_logic_vector(22, 8),
27957 => conv_std_logic_vector(22, 8),
27958 => conv_std_logic_vector(22, 8),
27959 => conv_std_logic_vector(23, 8),
27960 => conv_std_logic_vector(23, 8),
27961 => conv_std_logic_vector(24, 8),
27962 => conv_std_logic_vector(24, 8),
27963 => conv_std_logic_vector(25, 8),
27964 => conv_std_logic_vector(25, 8),
27965 => conv_std_logic_vector(25, 8),
27966 => conv_std_logic_vector(26, 8),
27967 => conv_std_logic_vector(26, 8),
27968 => conv_std_logic_vector(27, 8),
27969 => conv_std_logic_vector(27, 8),
27970 => conv_std_logic_vector(28, 8),
27971 => conv_std_logic_vector(28, 8),
27972 => conv_std_logic_vector(28, 8),
27973 => conv_std_logic_vector(29, 8),
27974 => conv_std_logic_vector(29, 8),
27975 => conv_std_logic_vector(30, 8),
27976 => conv_std_logic_vector(30, 8),
27977 => conv_std_logic_vector(31, 8),
27978 => conv_std_logic_vector(31, 8),
27979 => conv_std_logic_vector(31, 8),
27980 => conv_std_logic_vector(32, 8),
27981 => conv_std_logic_vector(32, 8),
27982 => conv_std_logic_vector(33, 8),
27983 => conv_std_logic_vector(33, 8),
27984 => conv_std_logic_vector(34, 8),
27985 => conv_std_logic_vector(34, 8),
27986 => conv_std_logic_vector(34, 8),
27987 => conv_std_logic_vector(35, 8),
27988 => conv_std_logic_vector(35, 8),
27989 => conv_std_logic_vector(36, 8),
27990 => conv_std_logic_vector(36, 8),
27991 => conv_std_logic_vector(37, 8),
27992 => conv_std_logic_vector(37, 8),
27993 => conv_std_logic_vector(37, 8),
27994 => conv_std_logic_vector(38, 8),
27995 => conv_std_logic_vector(38, 8),
27996 => conv_std_logic_vector(39, 8),
27997 => conv_std_logic_vector(39, 8),
27998 => conv_std_logic_vector(40, 8),
27999 => conv_std_logic_vector(40, 8),
28000 => conv_std_logic_vector(40, 8),
28001 => conv_std_logic_vector(41, 8),
28002 => conv_std_logic_vector(41, 8),
28003 => conv_std_logic_vector(42, 8),
28004 => conv_std_logic_vector(42, 8),
28005 => conv_std_logic_vector(43, 8),
28006 => conv_std_logic_vector(43, 8),
28007 => conv_std_logic_vector(43, 8),
28008 => conv_std_logic_vector(44, 8),
28009 => conv_std_logic_vector(44, 8),
28010 => conv_std_logic_vector(45, 8),
28011 => conv_std_logic_vector(45, 8),
28012 => conv_std_logic_vector(45, 8),
28013 => conv_std_logic_vector(46, 8),
28014 => conv_std_logic_vector(46, 8),
28015 => conv_std_logic_vector(47, 8),
28016 => conv_std_logic_vector(47, 8),
28017 => conv_std_logic_vector(48, 8),
28018 => conv_std_logic_vector(48, 8),
28019 => conv_std_logic_vector(48, 8),
28020 => conv_std_logic_vector(49, 8),
28021 => conv_std_logic_vector(49, 8),
28022 => conv_std_logic_vector(50, 8),
28023 => conv_std_logic_vector(50, 8),
28024 => conv_std_logic_vector(51, 8),
28025 => conv_std_logic_vector(51, 8),
28026 => conv_std_logic_vector(51, 8),
28027 => conv_std_logic_vector(52, 8),
28028 => conv_std_logic_vector(52, 8),
28029 => conv_std_logic_vector(53, 8),
28030 => conv_std_logic_vector(53, 8),
28031 => conv_std_logic_vector(54, 8),
28032 => conv_std_logic_vector(54, 8),
28033 => conv_std_logic_vector(54, 8),
28034 => conv_std_logic_vector(55, 8),
28035 => conv_std_logic_vector(55, 8),
28036 => conv_std_logic_vector(56, 8),
28037 => conv_std_logic_vector(56, 8),
28038 => conv_std_logic_vector(57, 8),
28039 => conv_std_logic_vector(57, 8),
28040 => conv_std_logic_vector(57, 8),
28041 => conv_std_logic_vector(58, 8),
28042 => conv_std_logic_vector(58, 8),
28043 => conv_std_logic_vector(59, 8),
28044 => conv_std_logic_vector(59, 8),
28045 => conv_std_logic_vector(60, 8),
28046 => conv_std_logic_vector(60, 8),
28047 => conv_std_logic_vector(60, 8),
28048 => conv_std_logic_vector(61, 8),
28049 => conv_std_logic_vector(61, 8),
28050 => conv_std_logic_vector(62, 8),
28051 => conv_std_logic_vector(62, 8),
28052 => conv_std_logic_vector(63, 8),
28053 => conv_std_logic_vector(63, 8),
28054 => conv_std_logic_vector(63, 8),
28055 => conv_std_logic_vector(64, 8),
28056 => conv_std_logic_vector(64, 8),
28057 => conv_std_logic_vector(65, 8),
28058 => conv_std_logic_vector(65, 8),
28059 => conv_std_logic_vector(65, 8),
28060 => conv_std_logic_vector(66, 8),
28061 => conv_std_logic_vector(66, 8),
28062 => conv_std_logic_vector(67, 8),
28063 => conv_std_logic_vector(67, 8),
28064 => conv_std_logic_vector(68, 8),
28065 => conv_std_logic_vector(68, 8),
28066 => conv_std_logic_vector(68, 8),
28067 => conv_std_logic_vector(69, 8),
28068 => conv_std_logic_vector(69, 8),
28069 => conv_std_logic_vector(70, 8),
28070 => conv_std_logic_vector(70, 8),
28071 => conv_std_logic_vector(71, 8),
28072 => conv_std_logic_vector(71, 8),
28073 => conv_std_logic_vector(71, 8),
28074 => conv_std_logic_vector(72, 8),
28075 => conv_std_logic_vector(72, 8),
28076 => conv_std_logic_vector(73, 8),
28077 => conv_std_logic_vector(73, 8),
28078 => conv_std_logic_vector(74, 8),
28079 => conv_std_logic_vector(74, 8),
28080 => conv_std_logic_vector(74, 8),
28081 => conv_std_logic_vector(75, 8),
28082 => conv_std_logic_vector(75, 8),
28083 => conv_std_logic_vector(76, 8),
28084 => conv_std_logic_vector(76, 8),
28085 => conv_std_logic_vector(77, 8),
28086 => conv_std_logic_vector(77, 8),
28087 => conv_std_logic_vector(77, 8),
28088 => conv_std_logic_vector(78, 8),
28089 => conv_std_logic_vector(78, 8),
28090 => conv_std_logic_vector(79, 8),
28091 => conv_std_logic_vector(79, 8),
28092 => conv_std_logic_vector(80, 8),
28093 => conv_std_logic_vector(80, 8),
28094 => conv_std_logic_vector(80, 8),
28095 => conv_std_logic_vector(81, 8),
28096 => conv_std_logic_vector(81, 8),
28097 => conv_std_logic_vector(82, 8),
28098 => conv_std_logic_vector(82, 8),
28099 => conv_std_logic_vector(83, 8),
28100 => conv_std_logic_vector(83, 8),
28101 => conv_std_logic_vector(83, 8),
28102 => conv_std_logic_vector(84, 8),
28103 => conv_std_logic_vector(84, 8),
28104 => conv_std_logic_vector(85, 8),
28105 => conv_std_logic_vector(85, 8),
28106 => conv_std_logic_vector(86, 8),
28107 => conv_std_logic_vector(86, 8),
28108 => conv_std_logic_vector(86, 8),
28109 => conv_std_logic_vector(87, 8),
28110 => conv_std_logic_vector(87, 8),
28111 => conv_std_logic_vector(88, 8),
28112 => conv_std_logic_vector(88, 8),
28113 => conv_std_logic_vector(88, 8),
28114 => conv_std_logic_vector(89, 8),
28115 => conv_std_logic_vector(89, 8),
28116 => conv_std_logic_vector(90, 8),
28117 => conv_std_logic_vector(90, 8),
28118 => conv_std_logic_vector(91, 8),
28119 => conv_std_logic_vector(91, 8),
28120 => conv_std_logic_vector(91, 8),
28121 => conv_std_logic_vector(92, 8),
28122 => conv_std_logic_vector(92, 8),
28123 => conv_std_logic_vector(93, 8),
28124 => conv_std_logic_vector(93, 8),
28125 => conv_std_logic_vector(94, 8),
28126 => conv_std_logic_vector(94, 8),
28127 => conv_std_logic_vector(94, 8),
28128 => conv_std_logic_vector(95, 8),
28129 => conv_std_logic_vector(95, 8),
28130 => conv_std_logic_vector(96, 8),
28131 => conv_std_logic_vector(96, 8),
28132 => conv_std_logic_vector(97, 8),
28133 => conv_std_logic_vector(97, 8),
28134 => conv_std_logic_vector(97, 8),
28135 => conv_std_logic_vector(98, 8),
28136 => conv_std_logic_vector(98, 8),
28137 => conv_std_logic_vector(99, 8),
28138 => conv_std_logic_vector(99, 8),
28139 => conv_std_logic_vector(100, 8),
28140 => conv_std_logic_vector(100, 8),
28141 => conv_std_logic_vector(100, 8),
28142 => conv_std_logic_vector(101, 8),
28143 => conv_std_logic_vector(101, 8),
28144 => conv_std_logic_vector(102, 8),
28145 => conv_std_logic_vector(102, 8),
28146 => conv_std_logic_vector(103, 8),
28147 => conv_std_logic_vector(103, 8),
28148 => conv_std_logic_vector(103, 8),
28149 => conv_std_logic_vector(104, 8),
28150 => conv_std_logic_vector(104, 8),
28151 => conv_std_logic_vector(105, 8),
28152 => conv_std_logic_vector(105, 8),
28153 => conv_std_logic_vector(106, 8),
28154 => conv_std_logic_vector(106, 8),
28155 => conv_std_logic_vector(106, 8),
28156 => conv_std_logic_vector(107, 8),
28157 => conv_std_logic_vector(107, 8),
28158 => conv_std_logic_vector(108, 8),
28159 => conv_std_logic_vector(108, 8),
28160 => conv_std_logic_vector(0, 8),
28161 => conv_std_logic_vector(0, 8),
28162 => conv_std_logic_vector(0, 8),
28163 => conv_std_logic_vector(1, 8),
28164 => conv_std_logic_vector(1, 8),
28165 => conv_std_logic_vector(2, 8),
28166 => conv_std_logic_vector(2, 8),
28167 => conv_std_logic_vector(3, 8),
28168 => conv_std_logic_vector(3, 8),
28169 => conv_std_logic_vector(3, 8),
28170 => conv_std_logic_vector(4, 8),
28171 => conv_std_logic_vector(4, 8),
28172 => conv_std_logic_vector(5, 8),
28173 => conv_std_logic_vector(5, 8),
28174 => conv_std_logic_vector(6, 8),
28175 => conv_std_logic_vector(6, 8),
28176 => conv_std_logic_vector(6, 8),
28177 => conv_std_logic_vector(7, 8),
28178 => conv_std_logic_vector(7, 8),
28179 => conv_std_logic_vector(8, 8),
28180 => conv_std_logic_vector(8, 8),
28181 => conv_std_logic_vector(9, 8),
28182 => conv_std_logic_vector(9, 8),
28183 => conv_std_logic_vector(9, 8),
28184 => conv_std_logic_vector(10, 8),
28185 => conv_std_logic_vector(10, 8),
28186 => conv_std_logic_vector(11, 8),
28187 => conv_std_logic_vector(11, 8),
28188 => conv_std_logic_vector(12, 8),
28189 => conv_std_logic_vector(12, 8),
28190 => conv_std_logic_vector(12, 8),
28191 => conv_std_logic_vector(13, 8),
28192 => conv_std_logic_vector(13, 8),
28193 => conv_std_logic_vector(14, 8),
28194 => conv_std_logic_vector(14, 8),
28195 => conv_std_logic_vector(15, 8),
28196 => conv_std_logic_vector(15, 8),
28197 => conv_std_logic_vector(15, 8),
28198 => conv_std_logic_vector(16, 8),
28199 => conv_std_logic_vector(16, 8),
28200 => conv_std_logic_vector(17, 8),
28201 => conv_std_logic_vector(17, 8),
28202 => conv_std_logic_vector(18, 8),
28203 => conv_std_logic_vector(18, 8),
28204 => conv_std_logic_vector(18, 8),
28205 => conv_std_logic_vector(19, 8),
28206 => conv_std_logic_vector(19, 8),
28207 => conv_std_logic_vector(20, 8),
28208 => conv_std_logic_vector(20, 8),
28209 => conv_std_logic_vector(21, 8),
28210 => conv_std_logic_vector(21, 8),
28211 => conv_std_logic_vector(21, 8),
28212 => conv_std_logic_vector(22, 8),
28213 => conv_std_logic_vector(22, 8),
28214 => conv_std_logic_vector(23, 8),
28215 => conv_std_logic_vector(23, 8),
28216 => conv_std_logic_vector(24, 8),
28217 => conv_std_logic_vector(24, 8),
28218 => conv_std_logic_vector(24, 8),
28219 => conv_std_logic_vector(25, 8),
28220 => conv_std_logic_vector(25, 8),
28221 => conv_std_logic_vector(26, 8),
28222 => conv_std_logic_vector(26, 8),
28223 => conv_std_logic_vector(27, 8),
28224 => conv_std_logic_vector(27, 8),
28225 => conv_std_logic_vector(27, 8),
28226 => conv_std_logic_vector(28, 8),
28227 => conv_std_logic_vector(28, 8),
28228 => conv_std_logic_vector(29, 8),
28229 => conv_std_logic_vector(29, 8),
28230 => conv_std_logic_vector(30, 8),
28231 => conv_std_logic_vector(30, 8),
28232 => conv_std_logic_vector(30, 8),
28233 => conv_std_logic_vector(31, 8),
28234 => conv_std_logic_vector(31, 8),
28235 => conv_std_logic_vector(32, 8),
28236 => conv_std_logic_vector(32, 8),
28237 => conv_std_logic_vector(33, 8),
28238 => conv_std_logic_vector(33, 8),
28239 => conv_std_logic_vector(33, 8),
28240 => conv_std_logic_vector(34, 8),
28241 => conv_std_logic_vector(34, 8),
28242 => conv_std_logic_vector(35, 8),
28243 => conv_std_logic_vector(35, 8),
28244 => conv_std_logic_vector(36, 8),
28245 => conv_std_logic_vector(36, 8),
28246 => conv_std_logic_vector(36, 8),
28247 => conv_std_logic_vector(37, 8),
28248 => conv_std_logic_vector(37, 8),
28249 => conv_std_logic_vector(38, 8),
28250 => conv_std_logic_vector(38, 8),
28251 => conv_std_logic_vector(39, 8),
28252 => conv_std_logic_vector(39, 8),
28253 => conv_std_logic_vector(39, 8),
28254 => conv_std_logic_vector(40, 8),
28255 => conv_std_logic_vector(40, 8),
28256 => conv_std_logic_vector(41, 8),
28257 => conv_std_logic_vector(41, 8),
28258 => conv_std_logic_vector(42, 8),
28259 => conv_std_logic_vector(42, 8),
28260 => conv_std_logic_vector(42, 8),
28261 => conv_std_logic_vector(43, 8),
28262 => conv_std_logic_vector(43, 8),
28263 => conv_std_logic_vector(44, 8),
28264 => conv_std_logic_vector(44, 8),
28265 => conv_std_logic_vector(45, 8),
28266 => conv_std_logic_vector(45, 8),
28267 => conv_std_logic_vector(45, 8),
28268 => conv_std_logic_vector(46, 8),
28269 => conv_std_logic_vector(46, 8),
28270 => conv_std_logic_vector(47, 8),
28271 => conv_std_logic_vector(47, 8),
28272 => conv_std_logic_vector(48, 8),
28273 => conv_std_logic_vector(48, 8),
28274 => conv_std_logic_vector(48, 8),
28275 => conv_std_logic_vector(49, 8),
28276 => conv_std_logic_vector(49, 8),
28277 => conv_std_logic_vector(50, 8),
28278 => conv_std_logic_vector(50, 8),
28279 => conv_std_logic_vector(51, 8),
28280 => conv_std_logic_vector(51, 8),
28281 => conv_std_logic_vector(51, 8),
28282 => conv_std_logic_vector(52, 8),
28283 => conv_std_logic_vector(52, 8),
28284 => conv_std_logic_vector(53, 8),
28285 => conv_std_logic_vector(53, 8),
28286 => conv_std_logic_vector(54, 8),
28287 => conv_std_logic_vector(54, 8),
28288 => conv_std_logic_vector(55, 8),
28289 => conv_std_logic_vector(55, 8),
28290 => conv_std_logic_vector(55, 8),
28291 => conv_std_logic_vector(56, 8),
28292 => conv_std_logic_vector(56, 8),
28293 => conv_std_logic_vector(57, 8),
28294 => conv_std_logic_vector(57, 8),
28295 => conv_std_logic_vector(58, 8),
28296 => conv_std_logic_vector(58, 8),
28297 => conv_std_logic_vector(58, 8),
28298 => conv_std_logic_vector(59, 8),
28299 => conv_std_logic_vector(59, 8),
28300 => conv_std_logic_vector(60, 8),
28301 => conv_std_logic_vector(60, 8),
28302 => conv_std_logic_vector(61, 8),
28303 => conv_std_logic_vector(61, 8),
28304 => conv_std_logic_vector(61, 8),
28305 => conv_std_logic_vector(62, 8),
28306 => conv_std_logic_vector(62, 8),
28307 => conv_std_logic_vector(63, 8),
28308 => conv_std_logic_vector(63, 8),
28309 => conv_std_logic_vector(64, 8),
28310 => conv_std_logic_vector(64, 8),
28311 => conv_std_logic_vector(64, 8),
28312 => conv_std_logic_vector(65, 8),
28313 => conv_std_logic_vector(65, 8),
28314 => conv_std_logic_vector(66, 8),
28315 => conv_std_logic_vector(66, 8),
28316 => conv_std_logic_vector(67, 8),
28317 => conv_std_logic_vector(67, 8),
28318 => conv_std_logic_vector(67, 8),
28319 => conv_std_logic_vector(68, 8),
28320 => conv_std_logic_vector(68, 8),
28321 => conv_std_logic_vector(69, 8),
28322 => conv_std_logic_vector(69, 8),
28323 => conv_std_logic_vector(70, 8),
28324 => conv_std_logic_vector(70, 8),
28325 => conv_std_logic_vector(70, 8),
28326 => conv_std_logic_vector(71, 8),
28327 => conv_std_logic_vector(71, 8),
28328 => conv_std_logic_vector(72, 8),
28329 => conv_std_logic_vector(72, 8),
28330 => conv_std_logic_vector(73, 8),
28331 => conv_std_logic_vector(73, 8),
28332 => conv_std_logic_vector(73, 8),
28333 => conv_std_logic_vector(74, 8),
28334 => conv_std_logic_vector(74, 8),
28335 => conv_std_logic_vector(75, 8),
28336 => conv_std_logic_vector(75, 8),
28337 => conv_std_logic_vector(76, 8),
28338 => conv_std_logic_vector(76, 8),
28339 => conv_std_logic_vector(76, 8),
28340 => conv_std_logic_vector(77, 8),
28341 => conv_std_logic_vector(77, 8),
28342 => conv_std_logic_vector(78, 8),
28343 => conv_std_logic_vector(78, 8),
28344 => conv_std_logic_vector(79, 8),
28345 => conv_std_logic_vector(79, 8),
28346 => conv_std_logic_vector(79, 8),
28347 => conv_std_logic_vector(80, 8),
28348 => conv_std_logic_vector(80, 8),
28349 => conv_std_logic_vector(81, 8),
28350 => conv_std_logic_vector(81, 8),
28351 => conv_std_logic_vector(82, 8),
28352 => conv_std_logic_vector(82, 8),
28353 => conv_std_logic_vector(82, 8),
28354 => conv_std_logic_vector(83, 8),
28355 => conv_std_logic_vector(83, 8),
28356 => conv_std_logic_vector(84, 8),
28357 => conv_std_logic_vector(84, 8),
28358 => conv_std_logic_vector(85, 8),
28359 => conv_std_logic_vector(85, 8),
28360 => conv_std_logic_vector(85, 8),
28361 => conv_std_logic_vector(86, 8),
28362 => conv_std_logic_vector(86, 8),
28363 => conv_std_logic_vector(87, 8),
28364 => conv_std_logic_vector(87, 8),
28365 => conv_std_logic_vector(88, 8),
28366 => conv_std_logic_vector(88, 8),
28367 => conv_std_logic_vector(88, 8),
28368 => conv_std_logic_vector(89, 8),
28369 => conv_std_logic_vector(89, 8),
28370 => conv_std_logic_vector(90, 8),
28371 => conv_std_logic_vector(90, 8),
28372 => conv_std_logic_vector(91, 8),
28373 => conv_std_logic_vector(91, 8),
28374 => conv_std_logic_vector(91, 8),
28375 => conv_std_logic_vector(92, 8),
28376 => conv_std_logic_vector(92, 8),
28377 => conv_std_logic_vector(93, 8),
28378 => conv_std_logic_vector(93, 8),
28379 => conv_std_logic_vector(94, 8),
28380 => conv_std_logic_vector(94, 8),
28381 => conv_std_logic_vector(94, 8),
28382 => conv_std_logic_vector(95, 8),
28383 => conv_std_logic_vector(95, 8),
28384 => conv_std_logic_vector(96, 8),
28385 => conv_std_logic_vector(96, 8),
28386 => conv_std_logic_vector(97, 8),
28387 => conv_std_logic_vector(97, 8),
28388 => conv_std_logic_vector(97, 8),
28389 => conv_std_logic_vector(98, 8),
28390 => conv_std_logic_vector(98, 8),
28391 => conv_std_logic_vector(99, 8),
28392 => conv_std_logic_vector(99, 8),
28393 => conv_std_logic_vector(100, 8),
28394 => conv_std_logic_vector(100, 8),
28395 => conv_std_logic_vector(100, 8),
28396 => conv_std_logic_vector(101, 8),
28397 => conv_std_logic_vector(101, 8),
28398 => conv_std_logic_vector(102, 8),
28399 => conv_std_logic_vector(102, 8),
28400 => conv_std_logic_vector(103, 8),
28401 => conv_std_logic_vector(103, 8),
28402 => conv_std_logic_vector(103, 8),
28403 => conv_std_logic_vector(104, 8),
28404 => conv_std_logic_vector(104, 8),
28405 => conv_std_logic_vector(105, 8),
28406 => conv_std_logic_vector(105, 8),
28407 => conv_std_logic_vector(106, 8),
28408 => conv_std_logic_vector(106, 8),
28409 => conv_std_logic_vector(106, 8),
28410 => conv_std_logic_vector(107, 8),
28411 => conv_std_logic_vector(107, 8),
28412 => conv_std_logic_vector(108, 8),
28413 => conv_std_logic_vector(108, 8),
28414 => conv_std_logic_vector(109, 8),
28415 => conv_std_logic_vector(109, 8),
28416 => conv_std_logic_vector(0, 8),
28417 => conv_std_logic_vector(0, 8),
28418 => conv_std_logic_vector(0, 8),
28419 => conv_std_logic_vector(1, 8),
28420 => conv_std_logic_vector(1, 8),
28421 => conv_std_logic_vector(2, 8),
28422 => conv_std_logic_vector(2, 8),
28423 => conv_std_logic_vector(3, 8),
28424 => conv_std_logic_vector(3, 8),
28425 => conv_std_logic_vector(3, 8),
28426 => conv_std_logic_vector(4, 8),
28427 => conv_std_logic_vector(4, 8),
28428 => conv_std_logic_vector(5, 8),
28429 => conv_std_logic_vector(5, 8),
28430 => conv_std_logic_vector(6, 8),
28431 => conv_std_logic_vector(6, 8),
28432 => conv_std_logic_vector(6, 8),
28433 => conv_std_logic_vector(7, 8),
28434 => conv_std_logic_vector(7, 8),
28435 => conv_std_logic_vector(8, 8),
28436 => conv_std_logic_vector(8, 8),
28437 => conv_std_logic_vector(9, 8),
28438 => conv_std_logic_vector(9, 8),
28439 => conv_std_logic_vector(9, 8),
28440 => conv_std_logic_vector(10, 8),
28441 => conv_std_logic_vector(10, 8),
28442 => conv_std_logic_vector(11, 8),
28443 => conv_std_logic_vector(11, 8),
28444 => conv_std_logic_vector(12, 8),
28445 => conv_std_logic_vector(12, 8),
28446 => conv_std_logic_vector(13, 8),
28447 => conv_std_logic_vector(13, 8),
28448 => conv_std_logic_vector(13, 8),
28449 => conv_std_logic_vector(14, 8),
28450 => conv_std_logic_vector(14, 8),
28451 => conv_std_logic_vector(15, 8),
28452 => conv_std_logic_vector(15, 8),
28453 => conv_std_logic_vector(16, 8),
28454 => conv_std_logic_vector(16, 8),
28455 => conv_std_logic_vector(16, 8),
28456 => conv_std_logic_vector(17, 8),
28457 => conv_std_logic_vector(17, 8),
28458 => conv_std_logic_vector(18, 8),
28459 => conv_std_logic_vector(18, 8),
28460 => conv_std_logic_vector(19, 8),
28461 => conv_std_logic_vector(19, 8),
28462 => conv_std_logic_vector(19, 8),
28463 => conv_std_logic_vector(20, 8),
28464 => conv_std_logic_vector(20, 8),
28465 => conv_std_logic_vector(21, 8),
28466 => conv_std_logic_vector(21, 8),
28467 => conv_std_logic_vector(22, 8),
28468 => conv_std_logic_vector(22, 8),
28469 => conv_std_logic_vector(22, 8),
28470 => conv_std_logic_vector(23, 8),
28471 => conv_std_logic_vector(23, 8),
28472 => conv_std_logic_vector(24, 8),
28473 => conv_std_logic_vector(24, 8),
28474 => conv_std_logic_vector(25, 8),
28475 => conv_std_logic_vector(25, 8),
28476 => conv_std_logic_vector(26, 8),
28477 => conv_std_logic_vector(26, 8),
28478 => conv_std_logic_vector(26, 8),
28479 => conv_std_logic_vector(27, 8),
28480 => conv_std_logic_vector(27, 8),
28481 => conv_std_logic_vector(28, 8),
28482 => conv_std_logic_vector(28, 8),
28483 => conv_std_logic_vector(29, 8),
28484 => conv_std_logic_vector(29, 8),
28485 => conv_std_logic_vector(29, 8),
28486 => conv_std_logic_vector(30, 8),
28487 => conv_std_logic_vector(30, 8),
28488 => conv_std_logic_vector(31, 8),
28489 => conv_std_logic_vector(31, 8),
28490 => conv_std_logic_vector(32, 8),
28491 => conv_std_logic_vector(32, 8),
28492 => conv_std_logic_vector(32, 8),
28493 => conv_std_logic_vector(33, 8),
28494 => conv_std_logic_vector(33, 8),
28495 => conv_std_logic_vector(34, 8),
28496 => conv_std_logic_vector(34, 8),
28497 => conv_std_logic_vector(35, 8),
28498 => conv_std_logic_vector(35, 8),
28499 => conv_std_logic_vector(35, 8),
28500 => conv_std_logic_vector(36, 8),
28501 => conv_std_logic_vector(36, 8),
28502 => conv_std_logic_vector(37, 8),
28503 => conv_std_logic_vector(37, 8),
28504 => conv_std_logic_vector(38, 8),
28505 => conv_std_logic_vector(38, 8),
28506 => conv_std_logic_vector(39, 8),
28507 => conv_std_logic_vector(39, 8),
28508 => conv_std_logic_vector(39, 8),
28509 => conv_std_logic_vector(40, 8),
28510 => conv_std_logic_vector(40, 8),
28511 => conv_std_logic_vector(41, 8),
28512 => conv_std_logic_vector(41, 8),
28513 => conv_std_logic_vector(42, 8),
28514 => conv_std_logic_vector(42, 8),
28515 => conv_std_logic_vector(42, 8),
28516 => conv_std_logic_vector(43, 8),
28517 => conv_std_logic_vector(43, 8),
28518 => conv_std_logic_vector(44, 8),
28519 => conv_std_logic_vector(44, 8),
28520 => conv_std_logic_vector(45, 8),
28521 => conv_std_logic_vector(45, 8),
28522 => conv_std_logic_vector(45, 8),
28523 => conv_std_logic_vector(46, 8),
28524 => conv_std_logic_vector(46, 8),
28525 => conv_std_logic_vector(47, 8),
28526 => conv_std_logic_vector(47, 8),
28527 => conv_std_logic_vector(48, 8),
28528 => conv_std_logic_vector(48, 8),
28529 => conv_std_logic_vector(48, 8),
28530 => conv_std_logic_vector(49, 8),
28531 => conv_std_logic_vector(49, 8),
28532 => conv_std_logic_vector(50, 8),
28533 => conv_std_logic_vector(50, 8),
28534 => conv_std_logic_vector(51, 8),
28535 => conv_std_logic_vector(51, 8),
28536 => conv_std_logic_vector(52, 8),
28537 => conv_std_logic_vector(52, 8),
28538 => conv_std_logic_vector(52, 8),
28539 => conv_std_logic_vector(53, 8),
28540 => conv_std_logic_vector(53, 8),
28541 => conv_std_logic_vector(54, 8),
28542 => conv_std_logic_vector(54, 8),
28543 => conv_std_logic_vector(55, 8),
28544 => conv_std_logic_vector(55, 8),
28545 => conv_std_logic_vector(55, 8),
28546 => conv_std_logic_vector(56, 8),
28547 => conv_std_logic_vector(56, 8),
28548 => conv_std_logic_vector(57, 8),
28549 => conv_std_logic_vector(57, 8),
28550 => conv_std_logic_vector(58, 8),
28551 => conv_std_logic_vector(58, 8),
28552 => conv_std_logic_vector(58, 8),
28553 => conv_std_logic_vector(59, 8),
28554 => conv_std_logic_vector(59, 8),
28555 => conv_std_logic_vector(60, 8),
28556 => conv_std_logic_vector(60, 8),
28557 => conv_std_logic_vector(61, 8),
28558 => conv_std_logic_vector(61, 8),
28559 => conv_std_logic_vector(62, 8),
28560 => conv_std_logic_vector(62, 8),
28561 => conv_std_logic_vector(62, 8),
28562 => conv_std_logic_vector(63, 8),
28563 => conv_std_logic_vector(63, 8),
28564 => conv_std_logic_vector(64, 8),
28565 => conv_std_logic_vector(64, 8),
28566 => conv_std_logic_vector(65, 8),
28567 => conv_std_logic_vector(65, 8),
28568 => conv_std_logic_vector(65, 8),
28569 => conv_std_logic_vector(66, 8),
28570 => conv_std_logic_vector(66, 8),
28571 => conv_std_logic_vector(67, 8),
28572 => conv_std_logic_vector(67, 8),
28573 => conv_std_logic_vector(68, 8),
28574 => conv_std_logic_vector(68, 8),
28575 => conv_std_logic_vector(68, 8),
28576 => conv_std_logic_vector(69, 8),
28577 => conv_std_logic_vector(69, 8),
28578 => conv_std_logic_vector(70, 8),
28579 => conv_std_logic_vector(70, 8),
28580 => conv_std_logic_vector(71, 8),
28581 => conv_std_logic_vector(71, 8),
28582 => conv_std_logic_vector(71, 8),
28583 => conv_std_logic_vector(72, 8),
28584 => conv_std_logic_vector(72, 8),
28585 => conv_std_logic_vector(73, 8),
28586 => conv_std_logic_vector(73, 8),
28587 => conv_std_logic_vector(74, 8),
28588 => conv_std_logic_vector(74, 8),
28589 => conv_std_logic_vector(75, 8),
28590 => conv_std_logic_vector(75, 8),
28591 => conv_std_logic_vector(75, 8),
28592 => conv_std_logic_vector(76, 8),
28593 => conv_std_logic_vector(76, 8),
28594 => conv_std_logic_vector(77, 8),
28595 => conv_std_logic_vector(77, 8),
28596 => conv_std_logic_vector(78, 8),
28597 => conv_std_logic_vector(78, 8),
28598 => conv_std_logic_vector(78, 8),
28599 => conv_std_logic_vector(79, 8),
28600 => conv_std_logic_vector(79, 8),
28601 => conv_std_logic_vector(80, 8),
28602 => conv_std_logic_vector(80, 8),
28603 => conv_std_logic_vector(81, 8),
28604 => conv_std_logic_vector(81, 8),
28605 => conv_std_logic_vector(81, 8),
28606 => conv_std_logic_vector(82, 8),
28607 => conv_std_logic_vector(82, 8),
28608 => conv_std_logic_vector(83, 8),
28609 => conv_std_logic_vector(83, 8),
28610 => conv_std_logic_vector(84, 8),
28611 => conv_std_logic_vector(84, 8),
28612 => conv_std_logic_vector(84, 8),
28613 => conv_std_logic_vector(85, 8),
28614 => conv_std_logic_vector(85, 8),
28615 => conv_std_logic_vector(86, 8),
28616 => conv_std_logic_vector(86, 8),
28617 => conv_std_logic_vector(87, 8),
28618 => conv_std_logic_vector(87, 8),
28619 => conv_std_logic_vector(88, 8),
28620 => conv_std_logic_vector(88, 8),
28621 => conv_std_logic_vector(88, 8),
28622 => conv_std_logic_vector(89, 8),
28623 => conv_std_logic_vector(89, 8),
28624 => conv_std_logic_vector(90, 8),
28625 => conv_std_logic_vector(90, 8),
28626 => conv_std_logic_vector(91, 8),
28627 => conv_std_logic_vector(91, 8),
28628 => conv_std_logic_vector(91, 8),
28629 => conv_std_logic_vector(92, 8),
28630 => conv_std_logic_vector(92, 8),
28631 => conv_std_logic_vector(93, 8),
28632 => conv_std_logic_vector(93, 8),
28633 => conv_std_logic_vector(94, 8),
28634 => conv_std_logic_vector(94, 8),
28635 => conv_std_logic_vector(94, 8),
28636 => conv_std_logic_vector(95, 8),
28637 => conv_std_logic_vector(95, 8),
28638 => conv_std_logic_vector(96, 8),
28639 => conv_std_logic_vector(96, 8),
28640 => conv_std_logic_vector(97, 8),
28641 => conv_std_logic_vector(97, 8),
28642 => conv_std_logic_vector(97, 8),
28643 => conv_std_logic_vector(98, 8),
28644 => conv_std_logic_vector(98, 8),
28645 => conv_std_logic_vector(99, 8),
28646 => conv_std_logic_vector(99, 8),
28647 => conv_std_logic_vector(100, 8),
28648 => conv_std_logic_vector(100, 8),
28649 => conv_std_logic_vector(101, 8),
28650 => conv_std_logic_vector(101, 8),
28651 => conv_std_logic_vector(101, 8),
28652 => conv_std_logic_vector(102, 8),
28653 => conv_std_logic_vector(102, 8),
28654 => conv_std_logic_vector(103, 8),
28655 => conv_std_logic_vector(103, 8),
28656 => conv_std_logic_vector(104, 8),
28657 => conv_std_logic_vector(104, 8),
28658 => conv_std_logic_vector(104, 8),
28659 => conv_std_logic_vector(105, 8),
28660 => conv_std_logic_vector(105, 8),
28661 => conv_std_logic_vector(106, 8),
28662 => conv_std_logic_vector(106, 8),
28663 => conv_std_logic_vector(107, 8),
28664 => conv_std_logic_vector(107, 8),
28665 => conv_std_logic_vector(107, 8),
28666 => conv_std_logic_vector(108, 8),
28667 => conv_std_logic_vector(108, 8),
28668 => conv_std_logic_vector(109, 8),
28669 => conv_std_logic_vector(109, 8),
28670 => conv_std_logic_vector(110, 8),
28671 => conv_std_logic_vector(110, 8),
28672 => conv_std_logic_vector(0, 8),
28673 => conv_std_logic_vector(0, 8),
28674 => conv_std_logic_vector(0, 8),
28675 => conv_std_logic_vector(1, 8),
28676 => conv_std_logic_vector(1, 8),
28677 => conv_std_logic_vector(2, 8),
28678 => conv_std_logic_vector(2, 8),
28679 => conv_std_logic_vector(3, 8),
28680 => conv_std_logic_vector(3, 8),
28681 => conv_std_logic_vector(3, 8),
28682 => conv_std_logic_vector(4, 8),
28683 => conv_std_logic_vector(4, 8),
28684 => conv_std_logic_vector(5, 8),
28685 => conv_std_logic_vector(5, 8),
28686 => conv_std_logic_vector(6, 8),
28687 => conv_std_logic_vector(6, 8),
28688 => conv_std_logic_vector(7, 8),
28689 => conv_std_logic_vector(7, 8),
28690 => conv_std_logic_vector(7, 8),
28691 => conv_std_logic_vector(8, 8),
28692 => conv_std_logic_vector(8, 8),
28693 => conv_std_logic_vector(9, 8),
28694 => conv_std_logic_vector(9, 8),
28695 => conv_std_logic_vector(10, 8),
28696 => conv_std_logic_vector(10, 8),
28697 => conv_std_logic_vector(10, 8),
28698 => conv_std_logic_vector(11, 8),
28699 => conv_std_logic_vector(11, 8),
28700 => conv_std_logic_vector(12, 8),
28701 => conv_std_logic_vector(12, 8),
28702 => conv_std_logic_vector(13, 8),
28703 => conv_std_logic_vector(13, 8),
28704 => conv_std_logic_vector(14, 8),
28705 => conv_std_logic_vector(14, 8),
28706 => conv_std_logic_vector(14, 8),
28707 => conv_std_logic_vector(15, 8),
28708 => conv_std_logic_vector(15, 8),
28709 => conv_std_logic_vector(16, 8),
28710 => conv_std_logic_vector(16, 8),
28711 => conv_std_logic_vector(17, 8),
28712 => conv_std_logic_vector(17, 8),
28713 => conv_std_logic_vector(17, 8),
28714 => conv_std_logic_vector(18, 8),
28715 => conv_std_logic_vector(18, 8),
28716 => conv_std_logic_vector(19, 8),
28717 => conv_std_logic_vector(19, 8),
28718 => conv_std_logic_vector(20, 8),
28719 => conv_std_logic_vector(20, 8),
28720 => conv_std_logic_vector(21, 8),
28721 => conv_std_logic_vector(21, 8),
28722 => conv_std_logic_vector(21, 8),
28723 => conv_std_logic_vector(22, 8),
28724 => conv_std_logic_vector(22, 8),
28725 => conv_std_logic_vector(23, 8),
28726 => conv_std_logic_vector(23, 8),
28727 => conv_std_logic_vector(24, 8),
28728 => conv_std_logic_vector(24, 8),
28729 => conv_std_logic_vector(24, 8),
28730 => conv_std_logic_vector(25, 8),
28731 => conv_std_logic_vector(25, 8),
28732 => conv_std_logic_vector(26, 8),
28733 => conv_std_logic_vector(26, 8),
28734 => conv_std_logic_vector(27, 8),
28735 => conv_std_logic_vector(27, 8),
28736 => conv_std_logic_vector(28, 8),
28737 => conv_std_logic_vector(28, 8),
28738 => conv_std_logic_vector(28, 8),
28739 => conv_std_logic_vector(29, 8),
28740 => conv_std_logic_vector(29, 8),
28741 => conv_std_logic_vector(30, 8),
28742 => conv_std_logic_vector(30, 8),
28743 => conv_std_logic_vector(31, 8),
28744 => conv_std_logic_vector(31, 8),
28745 => conv_std_logic_vector(31, 8),
28746 => conv_std_logic_vector(32, 8),
28747 => conv_std_logic_vector(32, 8),
28748 => conv_std_logic_vector(33, 8),
28749 => conv_std_logic_vector(33, 8),
28750 => conv_std_logic_vector(34, 8),
28751 => conv_std_logic_vector(34, 8),
28752 => conv_std_logic_vector(35, 8),
28753 => conv_std_logic_vector(35, 8),
28754 => conv_std_logic_vector(35, 8),
28755 => conv_std_logic_vector(36, 8),
28756 => conv_std_logic_vector(36, 8),
28757 => conv_std_logic_vector(37, 8),
28758 => conv_std_logic_vector(37, 8),
28759 => conv_std_logic_vector(38, 8),
28760 => conv_std_logic_vector(38, 8),
28761 => conv_std_logic_vector(38, 8),
28762 => conv_std_logic_vector(39, 8),
28763 => conv_std_logic_vector(39, 8),
28764 => conv_std_logic_vector(40, 8),
28765 => conv_std_logic_vector(40, 8),
28766 => conv_std_logic_vector(41, 8),
28767 => conv_std_logic_vector(41, 8),
28768 => conv_std_logic_vector(42, 8),
28769 => conv_std_logic_vector(42, 8),
28770 => conv_std_logic_vector(42, 8),
28771 => conv_std_logic_vector(43, 8),
28772 => conv_std_logic_vector(43, 8),
28773 => conv_std_logic_vector(44, 8),
28774 => conv_std_logic_vector(44, 8),
28775 => conv_std_logic_vector(45, 8),
28776 => conv_std_logic_vector(45, 8),
28777 => conv_std_logic_vector(45, 8),
28778 => conv_std_logic_vector(46, 8),
28779 => conv_std_logic_vector(46, 8),
28780 => conv_std_logic_vector(47, 8),
28781 => conv_std_logic_vector(47, 8),
28782 => conv_std_logic_vector(48, 8),
28783 => conv_std_logic_vector(48, 8),
28784 => conv_std_logic_vector(49, 8),
28785 => conv_std_logic_vector(49, 8),
28786 => conv_std_logic_vector(49, 8),
28787 => conv_std_logic_vector(50, 8),
28788 => conv_std_logic_vector(50, 8),
28789 => conv_std_logic_vector(51, 8),
28790 => conv_std_logic_vector(51, 8),
28791 => conv_std_logic_vector(52, 8),
28792 => conv_std_logic_vector(52, 8),
28793 => conv_std_logic_vector(52, 8),
28794 => conv_std_logic_vector(53, 8),
28795 => conv_std_logic_vector(53, 8),
28796 => conv_std_logic_vector(54, 8),
28797 => conv_std_logic_vector(54, 8),
28798 => conv_std_logic_vector(55, 8),
28799 => conv_std_logic_vector(55, 8),
28800 => conv_std_logic_vector(56, 8),
28801 => conv_std_logic_vector(56, 8),
28802 => conv_std_logic_vector(56, 8),
28803 => conv_std_logic_vector(57, 8),
28804 => conv_std_logic_vector(57, 8),
28805 => conv_std_logic_vector(58, 8),
28806 => conv_std_logic_vector(58, 8),
28807 => conv_std_logic_vector(59, 8),
28808 => conv_std_logic_vector(59, 8),
28809 => conv_std_logic_vector(59, 8),
28810 => conv_std_logic_vector(60, 8),
28811 => conv_std_logic_vector(60, 8),
28812 => conv_std_logic_vector(61, 8),
28813 => conv_std_logic_vector(61, 8),
28814 => conv_std_logic_vector(62, 8),
28815 => conv_std_logic_vector(62, 8),
28816 => conv_std_logic_vector(63, 8),
28817 => conv_std_logic_vector(63, 8),
28818 => conv_std_logic_vector(63, 8),
28819 => conv_std_logic_vector(64, 8),
28820 => conv_std_logic_vector(64, 8),
28821 => conv_std_logic_vector(65, 8),
28822 => conv_std_logic_vector(65, 8),
28823 => conv_std_logic_vector(66, 8),
28824 => conv_std_logic_vector(66, 8),
28825 => conv_std_logic_vector(66, 8),
28826 => conv_std_logic_vector(67, 8),
28827 => conv_std_logic_vector(67, 8),
28828 => conv_std_logic_vector(68, 8),
28829 => conv_std_logic_vector(68, 8),
28830 => conv_std_logic_vector(69, 8),
28831 => conv_std_logic_vector(69, 8),
28832 => conv_std_logic_vector(70, 8),
28833 => conv_std_logic_vector(70, 8),
28834 => conv_std_logic_vector(70, 8),
28835 => conv_std_logic_vector(71, 8),
28836 => conv_std_logic_vector(71, 8),
28837 => conv_std_logic_vector(72, 8),
28838 => conv_std_logic_vector(72, 8),
28839 => conv_std_logic_vector(73, 8),
28840 => conv_std_logic_vector(73, 8),
28841 => conv_std_logic_vector(73, 8),
28842 => conv_std_logic_vector(74, 8),
28843 => conv_std_logic_vector(74, 8),
28844 => conv_std_logic_vector(75, 8),
28845 => conv_std_logic_vector(75, 8),
28846 => conv_std_logic_vector(76, 8),
28847 => conv_std_logic_vector(76, 8),
28848 => conv_std_logic_vector(77, 8),
28849 => conv_std_logic_vector(77, 8),
28850 => conv_std_logic_vector(77, 8),
28851 => conv_std_logic_vector(78, 8),
28852 => conv_std_logic_vector(78, 8),
28853 => conv_std_logic_vector(79, 8),
28854 => conv_std_logic_vector(79, 8),
28855 => conv_std_logic_vector(80, 8),
28856 => conv_std_logic_vector(80, 8),
28857 => conv_std_logic_vector(80, 8),
28858 => conv_std_logic_vector(81, 8),
28859 => conv_std_logic_vector(81, 8),
28860 => conv_std_logic_vector(82, 8),
28861 => conv_std_logic_vector(82, 8),
28862 => conv_std_logic_vector(83, 8),
28863 => conv_std_logic_vector(83, 8),
28864 => conv_std_logic_vector(84, 8),
28865 => conv_std_logic_vector(84, 8),
28866 => conv_std_logic_vector(84, 8),
28867 => conv_std_logic_vector(85, 8),
28868 => conv_std_logic_vector(85, 8),
28869 => conv_std_logic_vector(86, 8),
28870 => conv_std_logic_vector(86, 8),
28871 => conv_std_logic_vector(87, 8),
28872 => conv_std_logic_vector(87, 8),
28873 => conv_std_logic_vector(87, 8),
28874 => conv_std_logic_vector(88, 8),
28875 => conv_std_logic_vector(88, 8),
28876 => conv_std_logic_vector(89, 8),
28877 => conv_std_logic_vector(89, 8),
28878 => conv_std_logic_vector(90, 8),
28879 => conv_std_logic_vector(90, 8),
28880 => conv_std_logic_vector(91, 8),
28881 => conv_std_logic_vector(91, 8),
28882 => conv_std_logic_vector(91, 8),
28883 => conv_std_logic_vector(92, 8),
28884 => conv_std_logic_vector(92, 8),
28885 => conv_std_logic_vector(93, 8),
28886 => conv_std_logic_vector(93, 8),
28887 => conv_std_logic_vector(94, 8),
28888 => conv_std_logic_vector(94, 8),
28889 => conv_std_logic_vector(94, 8),
28890 => conv_std_logic_vector(95, 8),
28891 => conv_std_logic_vector(95, 8),
28892 => conv_std_logic_vector(96, 8),
28893 => conv_std_logic_vector(96, 8),
28894 => conv_std_logic_vector(97, 8),
28895 => conv_std_logic_vector(97, 8),
28896 => conv_std_logic_vector(98, 8),
28897 => conv_std_logic_vector(98, 8),
28898 => conv_std_logic_vector(98, 8),
28899 => conv_std_logic_vector(99, 8),
28900 => conv_std_logic_vector(99, 8),
28901 => conv_std_logic_vector(100, 8),
28902 => conv_std_logic_vector(100, 8),
28903 => conv_std_logic_vector(101, 8),
28904 => conv_std_logic_vector(101, 8),
28905 => conv_std_logic_vector(101, 8),
28906 => conv_std_logic_vector(102, 8),
28907 => conv_std_logic_vector(102, 8),
28908 => conv_std_logic_vector(103, 8),
28909 => conv_std_logic_vector(103, 8),
28910 => conv_std_logic_vector(104, 8),
28911 => conv_std_logic_vector(104, 8),
28912 => conv_std_logic_vector(105, 8),
28913 => conv_std_logic_vector(105, 8),
28914 => conv_std_logic_vector(105, 8),
28915 => conv_std_logic_vector(106, 8),
28916 => conv_std_logic_vector(106, 8),
28917 => conv_std_logic_vector(107, 8),
28918 => conv_std_logic_vector(107, 8),
28919 => conv_std_logic_vector(108, 8),
28920 => conv_std_logic_vector(108, 8),
28921 => conv_std_logic_vector(108, 8),
28922 => conv_std_logic_vector(109, 8),
28923 => conv_std_logic_vector(109, 8),
28924 => conv_std_logic_vector(110, 8),
28925 => conv_std_logic_vector(110, 8),
28926 => conv_std_logic_vector(111, 8),
28927 => conv_std_logic_vector(111, 8),
28928 => conv_std_logic_vector(0, 8),
28929 => conv_std_logic_vector(0, 8),
28930 => conv_std_logic_vector(0, 8),
28931 => conv_std_logic_vector(1, 8),
28932 => conv_std_logic_vector(1, 8),
28933 => conv_std_logic_vector(2, 8),
28934 => conv_std_logic_vector(2, 8),
28935 => conv_std_logic_vector(3, 8),
28936 => conv_std_logic_vector(3, 8),
28937 => conv_std_logic_vector(3, 8),
28938 => conv_std_logic_vector(4, 8),
28939 => conv_std_logic_vector(4, 8),
28940 => conv_std_logic_vector(5, 8),
28941 => conv_std_logic_vector(5, 8),
28942 => conv_std_logic_vector(6, 8),
28943 => conv_std_logic_vector(6, 8),
28944 => conv_std_logic_vector(7, 8),
28945 => conv_std_logic_vector(7, 8),
28946 => conv_std_logic_vector(7, 8),
28947 => conv_std_logic_vector(8, 8),
28948 => conv_std_logic_vector(8, 8),
28949 => conv_std_logic_vector(9, 8),
28950 => conv_std_logic_vector(9, 8),
28951 => conv_std_logic_vector(10, 8),
28952 => conv_std_logic_vector(10, 8),
28953 => conv_std_logic_vector(11, 8),
28954 => conv_std_logic_vector(11, 8),
28955 => conv_std_logic_vector(11, 8),
28956 => conv_std_logic_vector(12, 8),
28957 => conv_std_logic_vector(12, 8),
28958 => conv_std_logic_vector(13, 8),
28959 => conv_std_logic_vector(13, 8),
28960 => conv_std_logic_vector(14, 8),
28961 => conv_std_logic_vector(14, 8),
28962 => conv_std_logic_vector(15, 8),
28963 => conv_std_logic_vector(15, 8),
28964 => conv_std_logic_vector(15, 8),
28965 => conv_std_logic_vector(16, 8),
28966 => conv_std_logic_vector(16, 8),
28967 => conv_std_logic_vector(17, 8),
28968 => conv_std_logic_vector(17, 8),
28969 => conv_std_logic_vector(18, 8),
28970 => conv_std_logic_vector(18, 8),
28971 => conv_std_logic_vector(18, 8),
28972 => conv_std_logic_vector(19, 8),
28973 => conv_std_logic_vector(19, 8),
28974 => conv_std_logic_vector(20, 8),
28975 => conv_std_logic_vector(20, 8),
28976 => conv_std_logic_vector(21, 8),
28977 => conv_std_logic_vector(21, 8),
28978 => conv_std_logic_vector(22, 8),
28979 => conv_std_logic_vector(22, 8),
28980 => conv_std_logic_vector(22, 8),
28981 => conv_std_logic_vector(23, 8),
28982 => conv_std_logic_vector(23, 8),
28983 => conv_std_logic_vector(24, 8),
28984 => conv_std_logic_vector(24, 8),
28985 => conv_std_logic_vector(25, 8),
28986 => conv_std_logic_vector(25, 8),
28987 => conv_std_logic_vector(26, 8),
28988 => conv_std_logic_vector(26, 8),
28989 => conv_std_logic_vector(26, 8),
28990 => conv_std_logic_vector(27, 8),
28991 => conv_std_logic_vector(27, 8),
28992 => conv_std_logic_vector(28, 8),
28993 => conv_std_logic_vector(28, 8),
28994 => conv_std_logic_vector(29, 8),
28995 => conv_std_logic_vector(29, 8),
28996 => conv_std_logic_vector(30, 8),
28997 => conv_std_logic_vector(30, 8),
28998 => conv_std_logic_vector(30, 8),
28999 => conv_std_logic_vector(31, 8),
29000 => conv_std_logic_vector(31, 8),
29001 => conv_std_logic_vector(32, 8),
29002 => conv_std_logic_vector(32, 8),
29003 => conv_std_logic_vector(33, 8),
29004 => conv_std_logic_vector(33, 8),
29005 => conv_std_logic_vector(33, 8),
29006 => conv_std_logic_vector(34, 8),
29007 => conv_std_logic_vector(34, 8),
29008 => conv_std_logic_vector(35, 8),
29009 => conv_std_logic_vector(35, 8),
29010 => conv_std_logic_vector(36, 8),
29011 => conv_std_logic_vector(36, 8),
29012 => conv_std_logic_vector(37, 8),
29013 => conv_std_logic_vector(37, 8),
29014 => conv_std_logic_vector(37, 8),
29015 => conv_std_logic_vector(38, 8),
29016 => conv_std_logic_vector(38, 8),
29017 => conv_std_logic_vector(39, 8),
29018 => conv_std_logic_vector(39, 8),
29019 => conv_std_logic_vector(40, 8),
29020 => conv_std_logic_vector(40, 8),
29021 => conv_std_logic_vector(41, 8),
29022 => conv_std_logic_vector(41, 8),
29023 => conv_std_logic_vector(41, 8),
29024 => conv_std_logic_vector(42, 8),
29025 => conv_std_logic_vector(42, 8),
29026 => conv_std_logic_vector(43, 8),
29027 => conv_std_logic_vector(43, 8),
29028 => conv_std_logic_vector(44, 8),
29029 => conv_std_logic_vector(44, 8),
29030 => conv_std_logic_vector(45, 8),
29031 => conv_std_logic_vector(45, 8),
29032 => conv_std_logic_vector(45, 8),
29033 => conv_std_logic_vector(46, 8),
29034 => conv_std_logic_vector(46, 8),
29035 => conv_std_logic_vector(47, 8),
29036 => conv_std_logic_vector(47, 8),
29037 => conv_std_logic_vector(48, 8),
29038 => conv_std_logic_vector(48, 8),
29039 => conv_std_logic_vector(48, 8),
29040 => conv_std_logic_vector(49, 8),
29041 => conv_std_logic_vector(49, 8),
29042 => conv_std_logic_vector(50, 8),
29043 => conv_std_logic_vector(50, 8),
29044 => conv_std_logic_vector(51, 8),
29045 => conv_std_logic_vector(51, 8),
29046 => conv_std_logic_vector(52, 8),
29047 => conv_std_logic_vector(52, 8),
29048 => conv_std_logic_vector(52, 8),
29049 => conv_std_logic_vector(53, 8),
29050 => conv_std_logic_vector(53, 8),
29051 => conv_std_logic_vector(54, 8),
29052 => conv_std_logic_vector(54, 8),
29053 => conv_std_logic_vector(55, 8),
29054 => conv_std_logic_vector(55, 8),
29055 => conv_std_logic_vector(56, 8),
29056 => conv_std_logic_vector(56, 8),
29057 => conv_std_logic_vector(56, 8),
29058 => conv_std_logic_vector(57, 8),
29059 => conv_std_logic_vector(57, 8),
29060 => conv_std_logic_vector(58, 8),
29061 => conv_std_logic_vector(58, 8),
29062 => conv_std_logic_vector(59, 8),
29063 => conv_std_logic_vector(59, 8),
29064 => conv_std_logic_vector(60, 8),
29065 => conv_std_logic_vector(60, 8),
29066 => conv_std_logic_vector(60, 8),
29067 => conv_std_logic_vector(61, 8),
29068 => conv_std_logic_vector(61, 8),
29069 => conv_std_logic_vector(62, 8),
29070 => conv_std_logic_vector(62, 8),
29071 => conv_std_logic_vector(63, 8),
29072 => conv_std_logic_vector(63, 8),
29073 => conv_std_logic_vector(64, 8),
29074 => conv_std_logic_vector(64, 8),
29075 => conv_std_logic_vector(64, 8),
29076 => conv_std_logic_vector(65, 8),
29077 => conv_std_logic_vector(65, 8),
29078 => conv_std_logic_vector(66, 8),
29079 => conv_std_logic_vector(66, 8),
29080 => conv_std_logic_vector(67, 8),
29081 => conv_std_logic_vector(67, 8),
29082 => conv_std_logic_vector(67, 8),
29083 => conv_std_logic_vector(68, 8),
29084 => conv_std_logic_vector(68, 8),
29085 => conv_std_logic_vector(69, 8),
29086 => conv_std_logic_vector(69, 8),
29087 => conv_std_logic_vector(70, 8),
29088 => conv_std_logic_vector(70, 8),
29089 => conv_std_logic_vector(71, 8),
29090 => conv_std_logic_vector(71, 8),
29091 => conv_std_logic_vector(71, 8),
29092 => conv_std_logic_vector(72, 8),
29093 => conv_std_logic_vector(72, 8),
29094 => conv_std_logic_vector(73, 8),
29095 => conv_std_logic_vector(73, 8),
29096 => conv_std_logic_vector(74, 8),
29097 => conv_std_logic_vector(74, 8),
29098 => conv_std_logic_vector(75, 8),
29099 => conv_std_logic_vector(75, 8),
29100 => conv_std_logic_vector(75, 8),
29101 => conv_std_logic_vector(76, 8),
29102 => conv_std_logic_vector(76, 8),
29103 => conv_std_logic_vector(77, 8),
29104 => conv_std_logic_vector(77, 8),
29105 => conv_std_logic_vector(78, 8),
29106 => conv_std_logic_vector(78, 8),
29107 => conv_std_logic_vector(79, 8),
29108 => conv_std_logic_vector(79, 8),
29109 => conv_std_logic_vector(79, 8),
29110 => conv_std_logic_vector(80, 8),
29111 => conv_std_logic_vector(80, 8),
29112 => conv_std_logic_vector(81, 8),
29113 => conv_std_logic_vector(81, 8),
29114 => conv_std_logic_vector(82, 8),
29115 => conv_std_logic_vector(82, 8),
29116 => conv_std_logic_vector(82, 8),
29117 => conv_std_logic_vector(83, 8),
29118 => conv_std_logic_vector(83, 8),
29119 => conv_std_logic_vector(84, 8),
29120 => conv_std_logic_vector(84, 8),
29121 => conv_std_logic_vector(85, 8),
29122 => conv_std_logic_vector(85, 8),
29123 => conv_std_logic_vector(86, 8),
29124 => conv_std_logic_vector(86, 8),
29125 => conv_std_logic_vector(86, 8),
29126 => conv_std_logic_vector(87, 8),
29127 => conv_std_logic_vector(87, 8),
29128 => conv_std_logic_vector(88, 8),
29129 => conv_std_logic_vector(88, 8),
29130 => conv_std_logic_vector(89, 8),
29131 => conv_std_logic_vector(89, 8),
29132 => conv_std_logic_vector(90, 8),
29133 => conv_std_logic_vector(90, 8),
29134 => conv_std_logic_vector(90, 8),
29135 => conv_std_logic_vector(91, 8),
29136 => conv_std_logic_vector(91, 8),
29137 => conv_std_logic_vector(92, 8),
29138 => conv_std_logic_vector(92, 8),
29139 => conv_std_logic_vector(93, 8),
29140 => conv_std_logic_vector(93, 8),
29141 => conv_std_logic_vector(94, 8),
29142 => conv_std_logic_vector(94, 8),
29143 => conv_std_logic_vector(94, 8),
29144 => conv_std_logic_vector(95, 8),
29145 => conv_std_logic_vector(95, 8),
29146 => conv_std_logic_vector(96, 8),
29147 => conv_std_logic_vector(96, 8),
29148 => conv_std_logic_vector(97, 8),
29149 => conv_std_logic_vector(97, 8),
29150 => conv_std_logic_vector(97, 8),
29151 => conv_std_logic_vector(98, 8),
29152 => conv_std_logic_vector(98, 8),
29153 => conv_std_logic_vector(99, 8),
29154 => conv_std_logic_vector(99, 8),
29155 => conv_std_logic_vector(100, 8),
29156 => conv_std_logic_vector(100, 8),
29157 => conv_std_logic_vector(101, 8),
29158 => conv_std_logic_vector(101, 8),
29159 => conv_std_logic_vector(101, 8),
29160 => conv_std_logic_vector(102, 8),
29161 => conv_std_logic_vector(102, 8),
29162 => conv_std_logic_vector(103, 8),
29163 => conv_std_logic_vector(103, 8),
29164 => conv_std_logic_vector(104, 8),
29165 => conv_std_logic_vector(104, 8),
29166 => conv_std_logic_vector(105, 8),
29167 => conv_std_logic_vector(105, 8),
29168 => conv_std_logic_vector(105, 8),
29169 => conv_std_logic_vector(106, 8),
29170 => conv_std_logic_vector(106, 8),
29171 => conv_std_logic_vector(107, 8),
29172 => conv_std_logic_vector(107, 8),
29173 => conv_std_logic_vector(108, 8),
29174 => conv_std_logic_vector(108, 8),
29175 => conv_std_logic_vector(109, 8),
29176 => conv_std_logic_vector(109, 8),
29177 => conv_std_logic_vector(109, 8),
29178 => conv_std_logic_vector(110, 8),
29179 => conv_std_logic_vector(110, 8),
29180 => conv_std_logic_vector(111, 8),
29181 => conv_std_logic_vector(111, 8),
29182 => conv_std_logic_vector(112, 8),
29183 => conv_std_logic_vector(112, 8),
29184 => conv_std_logic_vector(0, 8),
29185 => conv_std_logic_vector(0, 8),
29186 => conv_std_logic_vector(0, 8),
29187 => conv_std_logic_vector(1, 8),
29188 => conv_std_logic_vector(1, 8),
29189 => conv_std_logic_vector(2, 8),
29190 => conv_std_logic_vector(2, 8),
29191 => conv_std_logic_vector(3, 8),
29192 => conv_std_logic_vector(3, 8),
29193 => conv_std_logic_vector(4, 8),
29194 => conv_std_logic_vector(4, 8),
29195 => conv_std_logic_vector(4, 8),
29196 => conv_std_logic_vector(5, 8),
29197 => conv_std_logic_vector(5, 8),
29198 => conv_std_logic_vector(6, 8),
29199 => conv_std_logic_vector(6, 8),
29200 => conv_std_logic_vector(7, 8),
29201 => conv_std_logic_vector(7, 8),
29202 => conv_std_logic_vector(8, 8),
29203 => conv_std_logic_vector(8, 8),
29204 => conv_std_logic_vector(8, 8),
29205 => conv_std_logic_vector(9, 8),
29206 => conv_std_logic_vector(9, 8),
29207 => conv_std_logic_vector(10, 8),
29208 => conv_std_logic_vector(10, 8),
29209 => conv_std_logic_vector(11, 8),
29210 => conv_std_logic_vector(11, 8),
29211 => conv_std_logic_vector(12, 8),
29212 => conv_std_logic_vector(12, 8),
29213 => conv_std_logic_vector(12, 8),
29214 => conv_std_logic_vector(13, 8),
29215 => conv_std_logic_vector(13, 8),
29216 => conv_std_logic_vector(14, 8),
29217 => conv_std_logic_vector(14, 8),
29218 => conv_std_logic_vector(15, 8),
29219 => conv_std_logic_vector(15, 8),
29220 => conv_std_logic_vector(16, 8),
29221 => conv_std_logic_vector(16, 8),
29222 => conv_std_logic_vector(16, 8),
29223 => conv_std_logic_vector(17, 8),
29224 => conv_std_logic_vector(17, 8),
29225 => conv_std_logic_vector(18, 8),
29226 => conv_std_logic_vector(18, 8),
29227 => conv_std_logic_vector(19, 8),
29228 => conv_std_logic_vector(19, 8),
29229 => conv_std_logic_vector(20, 8),
29230 => conv_std_logic_vector(20, 8),
29231 => conv_std_logic_vector(20, 8),
29232 => conv_std_logic_vector(21, 8),
29233 => conv_std_logic_vector(21, 8),
29234 => conv_std_logic_vector(22, 8),
29235 => conv_std_logic_vector(22, 8),
29236 => conv_std_logic_vector(23, 8),
29237 => conv_std_logic_vector(23, 8),
29238 => conv_std_logic_vector(24, 8),
29239 => conv_std_logic_vector(24, 8),
29240 => conv_std_logic_vector(24, 8),
29241 => conv_std_logic_vector(25, 8),
29242 => conv_std_logic_vector(25, 8),
29243 => conv_std_logic_vector(26, 8),
29244 => conv_std_logic_vector(26, 8),
29245 => conv_std_logic_vector(27, 8),
29246 => conv_std_logic_vector(27, 8),
29247 => conv_std_logic_vector(28, 8),
29248 => conv_std_logic_vector(28, 8),
29249 => conv_std_logic_vector(28, 8),
29250 => conv_std_logic_vector(29, 8),
29251 => conv_std_logic_vector(29, 8),
29252 => conv_std_logic_vector(30, 8),
29253 => conv_std_logic_vector(30, 8),
29254 => conv_std_logic_vector(31, 8),
29255 => conv_std_logic_vector(31, 8),
29256 => conv_std_logic_vector(32, 8),
29257 => conv_std_logic_vector(32, 8),
29258 => conv_std_logic_vector(32, 8),
29259 => conv_std_logic_vector(33, 8),
29260 => conv_std_logic_vector(33, 8),
29261 => conv_std_logic_vector(34, 8),
29262 => conv_std_logic_vector(34, 8),
29263 => conv_std_logic_vector(35, 8),
29264 => conv_std_logic_vector(35, 8),
29265 => conv_std_logic_vector(36, 8),
29266 => conv_std_logic_vector(36, 8),
29267 => conv_std_logic_vector(36, 8),
29268 => conv_std_logic_vector(37, 8),
29269 => conv_std_logic_vector(37, 8),
29270 => conv_std_logic_vector(38, 8),
29271 => conv_std_logic_vector(38, 8),
29272 => conv_std_logic_vector(39, 8),
29273 => conv_std_logic_vector(39, 8),
29274 => conv_std_logic_vector(40, 8),
29275 => conv_std_logic_vector(40, 8),
29276 => conv_std_logic_vector(40, 8),
29277 => conv_std_logic_vector(41, 8),
29278 => conv_std_logic_vector(41, 8),
29279 => conv_std_logic_vector(42, 8),
29280 => conv_std_logic_vector(42, 8),
29281 => conv_std_logic_vector(43, 8),
29282 => conv_std_logic_vector(43, 8),
29283 => conv_std_logic_vector(44, 8),
29284 => conv_std_logic_vector(44, 8),
29285 => conv_std_logic_vector(44, 8),
29286 => conv_std_logic_vector(45, 8),
29287 => conv_std_logic_vector(45, 8),
29288 => conv_std_logic_vector(46, 8),
29289 => conv_std_logic_vector(46, 8),
29290 => conv_std_logic_vector(47, 8),
29291 => conv_std_logic_vector(47, 8),
29292 => conv_std_logic_vector(48, 8),
29293 => conv_std_logic_vector(48, 8),
29294 => conv_std_logic_vector(48, 8),
29295 => conv_std_logic_vector(49, 8),
29296 => conv_std_logic_vector(49, 8),
29297 => conv_std_logic_vector(50, 8),
29298 => conv_std_logic_vector(50, 8),
29299 => conv_std_logic_vector(51, 8),
29300 => conv_std_logic_vector(51, 8),
29301 => conv_std_logic_vector(52, 8),
29302 => conv_std_logic_vector(52, 8),
29303 => conv_std_logic_vector(52, 8),
29304 => conv_std_logic_vector(53, 8),
29305 => conv_std_logic_vector(53, 8),
29306 => conv_std_logic_vector(54, 8),
29307 => conv_std_logic_vector(54, 8),
29308 => conv_std_logic_vector(55, 8),
29309 => conv_std_logic_vector(55, 8),
29310 => conv_std_logic_vector(56, 8),
29311 => conv_std_logic_vector(56, 8),
29312 => conv_std_logic_vector(57, 8),
29313 => conv_std_logic_vector(57, 8),
29314 => conv_std_logic_vector(57, 8),
29315 => conv_std_logic_vector(58, 8),
29316 => conv_std_logic_vector(58, 8),
29317 => conv_std_logic_vector(59, 8),
29318 => conv_std_logic_vector(59, 8),
29319 => conv_std_logic_vector(60, 8),
29320 => conv_std_logic_vector(60, 8),
29321 => conv_std_logic_vector(61, 8),
29322 => conv_std_logic_vector(61, 8),
29323 => conv_std_logic_vector(61, 8),
29324 => conv_std_logic_vector(62, 8),
29325 => conv_std_logic_vector(62, 8),
29326 => conv_std_logic_vector(63, 8),
29327 => conv_std_logic_vector(63, 8),
29328 => conv_std_logic_vector(64, 8),
29329 => conv_std_logic_vector(64, 8),
29330 => conv_std_logic_vector(65, 8),
29331 => conv_std_logic_vector(65, 8),
29332 => conv_std_logic_vector(65, 8),
29333 => conv_std_logic_vector(66, 8),
29334 => conv_std_logic_vector(66, 8),
29335 => conv_std_logic_vector(67, 8),
29336 => conv_std_logic_vector(67, 8),
29337 => conv_std_logic_vector(68, 8),
29338 => conv_std_logic_vector(68, 8),
29339 => conv_std_logic_vector(69, 8),
29340 => conv_std_logic_vector(69, 8),
29341 => conv_std_logic_vector(69, 8),
29342 => conv_std_logic_vector(70, 8),
29343 => conv_std_logic_vector(70, 8),
29344 => conv_std_logic_vector(71, 8),
29345 => conv_std_logic_vector(71, 8),
29346 => conv_std_logic_vector(72, 8),
29347 => conv_std_logic_vector(72, 8),
29348 => conv_std_logic_vector(73, 8),
29349 => conv_std_logic_vector(73, 8),
29350 => conv_std_logic_vector(73, 8),
29351 => conv_std_logic_vector(74, 8),
29352 => conv_std_logic_vector(74, 8),
29353 => conv_std_logic_vector(75, 8),
29354 => conv_std_logic_vector(75, 8),
29355 => conv_std_logic_vector(76, 8),
29356 => conv_std_logic_vector(76, 8),
29357 => conv_std_logic_vector(77, 8),
29358 => conv_std_logic_vector(77, 8),
29359 => conv_std_logic_vector(77, 8),
29360 => conv_std_logic_vector(78, 8),
29361 => conv_std_logic_vector(78, 8),
29362 => conv_std_logic_vector(79, 8),
29363 => conv_std_logic_vector(79, 8),
29364 => conv_std_logic_vector(80, 8),
29365 => conv_std_logic_vector(80, 8),
29366 => conv_std_logic_vector(81, 8),
29367 => conv_std_logic_vector(81, 8),
29368 => conv_std_logic_vector(81, 8),
29369 => conv_std_logic_vector(82, 8),
29370 => conv_std_logic_vector(82, 8),
29371 => conv_std_logic_vector(83, 8),
29372 => conv_std_logic_vector(83, 8),
29373 => conv_std_logic_vector(84, 8),
29374 => conv_std_logic_vector(84, 8),
29375 => conv_std_logic_vector(85, 8),
29376 => conv_std_logic_vector(85, 8),
29377 => conv_std_logic_vector(85, 8),
29378 => conv_std_logic_vector(86, 8),
29379 => conv_std_logic_vector(86, 8),
29380 => conv_std_logic_vector(87, 8),
29381 => conv_std_logic_vector(87, 8),
29382 => conv_std_logic_vector(88, 8),
29383 => conv_std_logic_vector(88, 8),
29384 => conv_std_logic_vector(89, 8),
29385 => conv_std_logic_vector(89, 8),
29386 => conv_std_logic_vector(89, 8),
29387 => conv_std_logic_vector(90, 8),
29388 => conv_std_logic_vector(90, 8),
29389 => conv_std_logic_vector(91, 8),
29390 => conv_std_logic_vector(91, 8),
29391 => conv_std_logic_vector(92, 8),
29392 => conv_std_logic_vector(92, 8),
29393 => conv_std_logic_vector(93, 8),
29394 => conv_std_logic_vector(93, 8),
29395 => conv_std_logic_vector(93, 8),
29396 => conv_std_logic_vector(94, 8),
29397 => conv_std_logic_vector(94, 8),
29398 => conv_std_logic_vector(95, 8),
29399 => conv_std_logic_vector(95, 8),
29400 => conv_std_logic_vector(96, 8),
29401 => conv_std_logic_vector(96, 8),
29402 => conv_std_logic_vector(97, 8),
29403 => conv_std_logic_vector(97, 8),
29404 => conv_std_logic_vector(97, 8),
29405 => conv_std_logic_vector(98, 8),
29406 => conv_std_logic_vector(98, 8),
29407 => conv_std_logic_vector(99, 8),
29408 => conv_std_logic_vector(99, 8),
29409 => conv_std_logic_vector(100, 8),
29410 => conv_std_logic_vector(100, 8),
29411 => conv_std_logic_vector(101, 8),
29412 => conv_std_logic_vector(101, 8),
29413 => conv_std_logic_vector(101, 8),
29414 => conv_std_logic_vector(102, 8),
29415 => conv_std_logic_vector(102, 8),
29416 => conv_std_logic_vector(103, 8),
29417 => conv_std_logic_vector(103, 8),
29418 => conv_std_logic_vector(104, 8),
29419 => conv_std_logic_vector(104, 8),
29420 => conv_std_logic_vector(105, 8),
29421 => conv_std_logic_vector(105, 8),
29422 => conv_std_logic_vector(105, 8),
29423 => conv_std_logic_vector(106, 8),
29424 => conv_std_logic_vector(106, 8),
29425 => conv_std_logic_vector(107, 8),
29426 => conv_std_logic_vector(107, 8),
29427 => conv_std_logic_vector(108, 8),
29428 => conv_std_logic_vector(108, 8),
29429 => conv_std_logic_vector(109, 8),
29430 => conv_std_logic_vector(109, 8),
29431 => conv_std_logic_vector(109, 8),
29432 => conv_std_logic_vector(110, 8),
29433 => conv_std_logic_vector(110, 8),
29434 => conv_std_logic_vector(111, 8),
29435 => conv_std_logic_vector(111, 8),
29436 => conv_std_logic_vector(112, 8),
29437 => conv_std_logic_vector(112, 8),
29438 => conv_std_logic_vector(113, 8),
29439 => conv_std_logic_vector(113, 8),
29440 => conv_std_logic_vector(0, 8),
29441 => conv_std_logic_vector(0, 8),
29442 => conv_std_logic_vector(0, 8),
29443 => conv_std_logic_vector(1, 8),
29444 => conv_std_logic_vector(1, 8),
29445 => conv_std_logic_vector(2, 8),
29446 => conv_std_logic_vector(2, 8),
29447 => conv_std_logic_vector(3, 8),
29448 => conv_std_logic_vector(3, 8),
29449 => conv_std_logic_vector(4, 8),
29450 => conv_std_logic_vector(4, 8),
29451 => conv_std_logic_vector(4, 8),
29452 => conv_std_logic_vector(5, 8),
29453 => conv_std_logic_vector(5, 8),
29454 => conv_std_logic_vector(6, 8),
29455 => conv_std_logic_vector(6, 8),
29456 => conv_std_logic_vector(7, 8),
29457 => conv_std_logic_vector(7, 8),
29458 => conv_std_logic_vector(8, 8),
29459 => conv_std_logic_vector(8, 8),
29460 => conv_std_logic_vector(8, 8),
29461 => conv_std_logic_vector(9, 8),
29462 => conv_std_logic_vector(9, 8),
29463 => conv_std_logic_vector(10, 8),
29464 => conv_std_logic_vector(10, 8),
29465 => conv_std_logic_vector(11, 8),
29466 => conv_std_logic_vector(11, 8),
29467 => conv_std_logic_vector(12, 8),
29468 => conv_std_logic_vector(12, 8),
29469 => conv_std_logic_vector(13, 8),
29470 => conv_std_logic_vector(13, 8),
29471 => conv_std_logic_vector(13, 8),
29472 => conv_std_logic_vector(14, 8),
29473 => conv_std_logic_vector(14, 8),
29474 => conv_std_logic_vector(15, 8),
29475 => conv_std_logic_vector(15, 8),
29476 => conv_std_logic_vector(16, 8),
29477 => conv_std_logic_vector(16, 8),
29478 => conv_std_logic_vector(17, 8),
29479 => conv_std_logic_vector(17, 8),
29480 => conv_std_logic_vector(17, 8),
29481 => conv_std_logic_vector(18, 8),
29482 => conv_std_logic_vector(18, 8),
29483 => conv_std_logic_vector(19, 8),
29484 => conv_std_logic_vector(19, 8),
29485 => conv_std_logic_vector(20, 8),
29486 => conv_std_logic_vector(20, 8),
29487 => conv_std_logic_vector(21, 8),
29488 => conv_std_logic_vector(21, 8),
29489 => conv_std_logic_vector(22, 8),
29490 => conv_std_logic_vector(22, 8),
29491 => conv_std_logic_vector(22, 8),
29492 => conv_std_logic_vector(23, 8),
29493 => conv_std_logic_vector(23, 8),
29494 => conv_std_logic_vector(24, 8),
29495 => conv_std_logic_vector(24, 8),
29496 => conv_std_logic_vector(25, 8),
29497 => conv_std_logic_vector(25, 8),
29498 => conv_std_logic_vector(26, 8),
29499 => conv_std_logic_vector(26, 8),
29500 => conv_std_logic_vector(26, 8),
29501 => conv_std_logic_vector(27, 8),
29502 => conv_std_logic_vector(27, 8),
29503 => conv_std_logic_vector(28, 8),
29504 => conv_std_logic_vector(28, 8),
29505 => conv_std_logic_vector(29, 8),
29506 => conv_std_logic_vector(29, 8),
29507 => conv_std_logic_vector(30, 8),
29508 => conv_std_logic_vector(30, 8),
29509 => conv_std_logic_vector(30, 8),
29510 => conv_std_logic_vector(31, 8),
29511 => conv_std_logic_vector(31, 8),
29512 => conv_std_logic_vector(32, 8),
29513 => conv_std_logic_vector(32, 8),
29514 => conv_std_logic_vector(33, 8),
29515 => conv_std_logic_vector(33, 8),
29516 => conv_std_logic_vector(34, 8),
29517 => conv_std_logic_vector(34, 8),
29518 => conv_std_logic_vector(35, 8),
29519 => conv_std_logic_vector(35, 8),
29520 => conv_std_logic_vector(35, 8),
29521 => conv_std_logic_vector(36, 8),
29522 => conv_std_logic_vector(36, 8),
29523 => conv_std_logic_vector(37, 8),
29524 => conv_std_logic_vector(37, 8),
29525 => conv_std_logic_vector(38, 8),
29526 => conv_std_logic_vector(38, 8),
29527 => conv_std_logic_vector(39, 8),
29528 => conv_std_logic_vector(39, 8),
29529 => conv_std_logic_vector(39, 8),
29530 => conv_std_logic_vector(40, 8),
29531 => conv_std_logic_vector(40, 8),
29532 => conv_std_logic_vector(41, 8),
29533 => conv_std_logic_vector(41, 8),
29534 => conv_std_logic_vector(42, 8),
29535 => conv_std_logic_vector(42, 8),
29536 => conv_std_logic_vector(43, 8),
29537 => conv_std_logic_vector(43, 8),
29538 => conv_std_logic_vector(44, 8),
29539 => conv_std_logic_vector(44, 8),
29540 => conv_std_logic_vector(44, 8),
29541 => conv_std_logic_vector(45, 8),
29542 => conv_std_logic_vector(45, 8),
29543 => conv_std_logic_vector(46, 8),
29544 => conv_std_logic_vector(46, 8),
29545 => conv_std_logic_vector(47, 8),
29546 => conv_std_logic_vector(47, 8),
29547 => conv_std_logic_vector(48, 8),
29548 => conv_std_logic_vector(48, 8),
29549 => conv_std_logic_vector(48, 8),
29550 => conv_std_logic_vector(49, 8),
29551 => conv_std_logic_vector(49, 8),
29552 => conv_std_logic_vector(50, 8),
29553 => conv_std_logic_vector(50, 8),
29554 => conv_std_logic_vector(51, 8),
29555 => conv_std_logic_vector(51, 8),
29556 => conv_std_logic_vector(52, 8),
29557 => conv_std_logic_vector(52, 8),
29558 => conv_std_logic_vector(53, 8),
29559 => conv_std_logic_vector(53, 8),
29560 => conv_std_logic_vector(53, 8),
29561 => conv_std_logic_vector(54, 8),
29562 => conv_std_logic_vector(54, 8),
29563 => conv_std_logic_vector(55, 8),
29564 => conv_std_logic_vector(55, 8),
29565 => conv_std_logic_vector(56, 8),
29566 => conv_std_logic_vector(56, 8),
29567 => conv_std_logic_vector(57, 8),
29568 => conv_std_logic_vector(57, 8),
29569 => conv_std_logic_vector(57, 8),
29570 => conv_std_logic_vector(58, 8),
29571 => conv_std_logic_vector(58, 8),
29572 => conv_std_logic_vector(59, 8),
29573 => conv_std_logic_vector(59, 8),
29574 => conv_std_logic_vector(60, 8),
29575 => conv_std_logic_vector(60, 8),
29576 => conv_std_logic_vector(61, 8),
29577 => conv_std_logic_vector(61, 8),
29578 => conv_std_logic_vector(61, 8),
29579 => conv_std_logic_vector(62, 8),
29580 => conv_std_logic_vector(62, 8),
29581 => conv_std_logic_vector(63, 8),
29582 => conv_std_logic_vector(63, 8),
29583 => conv_std_logic_vector(64, 8),
29584 => conv_std_logic_vector(64, 8),
29585 => conv_std_logic_vector(65, 8),
29586 => conv_std_logic_vector(65, 8),
29587 => conv_std_logic_vector(66, 8),
29588 => conv_std_logic_vector(66, 8),
29589 => conv_std_logic_vector(66, 8),
29590 => conv_std_logic_vector(67, 8),
29591 => conv_std_logic_vector(67, 8),
29592 => conv_std_logic_vector(68, 8),
29593 => conv_std_logic_vector(68, 8),
29594 => conv_std_logic_vector(69, 8),
29595 => conv_std_logic_vector(69, 8),
29596 => conv_std_logic_vector(70, 8),
29597 => conv_std_logic_vector(70, 8),
29598 => conv_std_logic_vector(70, 8),
29599 => conv_std_logic_vector(71, 8),
29600 => conv_std_logic_vector(71, 8),
29601 => conv_std_logic_vector(72, 8),
29602 => conv_std_logic_vector(72, 8),
29603 => conv_std_logic_vector(73, 8),
29604 => conv_std_logic_vector(73, 8),
29605 => conv_std_logic_vector(74, 8),
29606 => conv_std_logic_vector(74, 8),
29607 => conv_std_logic_vector(75, 8),
29608 => conv_std_logic_vector(75, 8),
29609 => conv_std_logic_vector(75, 8),
29610 => conv_std_logic_vector(76, 8),
29611 => conv_std_logic_vector(76, 8),
29612 => conv_std_logic_vector(77, 8),
29613 => conv_std_logic_vector(77, 8),
29614 => conv_std_logic_vector(78, 8),
29615 => conv_std_logic_vector(78, 8),
29616 => conv_std_logic_vector(79, 8),
29617 => conv_std_logic_vector(79, 8),
29618 => conv_std_logic_vector(79, 8),
29619 => conv_std_logic_vector(80, 8),
29620 => conv_std_logic_vector(80, 8),
29621 => conv_std_logic_vector(81, 8),
29622 => conv_std_logic_vector(81, 8),
29623 => conv_std_logic_vector(82, 8),
29624 => conv_std_logic_vector(82, 8),
29625 => conv_std_logic_vector(83, 8),
29626 => conv_std_logic_vector(83, 8),
29627 => conv_std_logic_vector(84, 8),
29628 => conv_std_logic_vector(84, 8),
29629 => conv_std_logic_vector(84, 8),
29630 => conv_std_logic_vector(85, 8),
29631 => conv_std_logic_vector(85, 8),
29632 => conv_std_logic_vector(86, 8),
29633 => conv_std_logic_vector(86, 8),
29634 => conv_std_logic_vector(87, 8),
29635 => conv_std_logic_vector(87, 8),
29636 => conv_std_logic_vector(88, 8),
29637 => conv_std_logic_vector(88, 8),
29638 => conv_std_logic_vector(88, 8),
29639 => conv_std_logic_vector(89, 8),
29640 => conv_std_logic_vector(89, 8),
29641 => conv_std_logic_vector(90, 8),
29642 => conv_std_logic_vector(90, 8),
29643 => conv_std_logic_vector(91, 8),
29644 => conv_std_logic_vector(91, 8),
29645 => conv_std_logic_vector(92, 8),
29646 => conv_std_logic_vector(92, 8),
29647 => conv_std_logic_vector(92, 8),
29648 => conv_std_logic_vector(93, 8),
29649 => conv_std_logic_vector(93, 8),
29650 => conv_std_logic_vector(94, 8),
29651 => conv_std_logic_vector(94, 8),
29652 => conv_std_logic_vector(95, 8),
29653 => conv_std_logic_vector(95, 8),
29654 => conv_std_logic_vector(96, 8),
29655 => conv_std_logic_vector(96, 8),
29656 => conv_std_logic_vector(97, 8),
29657 => conv_std_logic_vector(97, 8),
29658 => conv_std_logic_vector(97, 8),
29659 => conv_std_logic_vector(98, 8),
29660 => conv_std_logic_vector(98, 8),
29661 => conv_std_logic_vector(99, 8),
29662 => conv_std_logic_vector(99, 8),
29663 => conv_std_logic_vector(100, 8),
29664 => conv_std_logic_vector(100, 8),
29665 => conv_std_logic_vector(101, 8),
29666 => conv_std_logic_vector(101, 8),
29667 => conv_std_logic_vector(101, 8),
29668 => conv_std_logic_vector(102, 8),
29669 => conv_std_logic_vector(102, 8),
29670 => conv_std_logic_vector(103, 8),
29671 => conv_std_logic_vector(103, 8),
29672 => conv_std_logic_vector(104, 8),
29673 => conv_std_logic_vector(104, 8),
29674 => conv_std_logic_vector(105, 8),
29675 => conv_std_logic_vector(105, 8),
29676 => conv_std_logic_vector(106, 8),
29677 => conv_std_logic_vector(106, 8),
29678 => conv_std_logic_vector(106, 8),
29679 => conv_std_logic_vector(107, 8),
29680 => conv_std_logic_vector(107, 8),
29681 => conv_std_logic_vector(108, 8),
29682 => conv_std_logic_vector(108, 8),
29683 => conv_std_logic_vector(109, 8),
29684 => conv_std_logic_vector(109, 8),
29685 => conv_std_logic_vector(110, 8),
29686 => conv_std_logic_vector(110, 8),
29687 => conv_std_logic_vector(110, 8),
29688 => conv_std_logic_vector(111, 8),
29689 => conv_std_logic_vector(111, 8),
29690 => conv_std_logic_vector(112, 8),
29691 => conv_std_logic_vector(112, 8),
29692 => conv_std_logic_vector(113, 8),
29693 => conv_std_logic_vector(113, 8),
29694 => conv_std_logic_vector(114, 8),
29695 => conv_std_logic_vector(114, 8),
29696 => conv_std_logic_vector(0, 8),
29697 => conv_std_logic_vector(0, 8),
29698 => conv_std_logic_vector(0, 8),
29699 => conv_std_logic_vector(1, 8),
29700 => conv_std_logic_vector(1, 8),
29701 => conv_std_logic_vector(2, 8),
29702 => conv_std_logic_vector(2, 8),
29703 => conv_std_logic_vector(3, 8),
29704 => conv_std_logic_vector(3, 8),
29705 => conv_std_logic_vector(4, 8),
29706 => conv_std_logic_vector(4, 8),
29707 => conv_std_logic_vector(4, 8),
29708 => conv_std_logic_vector(5, 8),
29709 => conv_std_logic_vector(5, 8),
29710 => conv_std_logic_vector(6, 8),
29711 => conv_std_logic_vector(6, 8),
29712 => conv_std_logic_vector(7, 8),
29713 => conv_std_logic_vector(7, 8),
29714 => conv_std_logic_vector(8, 8),
29715 => conv_std_logic_vector(8, 8),
29716 => conv_std_logic_vector(9, 8),
29717 => conv_std_logic_vector(9, 8),
29718 => conv_std_logic_vector(9, 8),
29719 => conv_std_logic_vector(10, 8),
29720 => conv_std_logic_vector(10, 8),
29721 => conv_std_logic_vector(11, 8),
29722 => conv_std_logic_vector(11, 8),
29723 => conv_std_logic_vector(12, 8),
29724 => conv_std_logic_vector(12, 8),
29725 => conv_std_logic_vector(13, 8),
29726 => conv_std_logic_vector(13, 8),
29727 => conv_std_logic_vector(14, 8),
29728 => conv_std_logic_vector(14, 8),
29729 => conv_std_logic_vector(14, 8),
29730 => conv_std_logic_vector(15, 8),
29731 => conv_std_logic_vector(15, 8),
29732 => conv_std_logic_vector(16, 8),
29733 => conv_std_logic_vector(16, 8),
29734 => conv_std_logic_vector(17, 8),
29735 => conv_std_logic_vector(17, 8),
29736 => conv_std_logic_vector(18, 8),
29737 => conv_std_logic_vector(18, 8),
29738 => conv_std_logic_vector(19, 8),
29739 => conv_std_logic_vector(19, 8),
29740 => conv_std_logic_vector(19, 8),
29741 => conv_std_logic_vector(20, 8),
29742 => conv_std_logic_vector(20, 8),
29743 => conv_std_logic_vector(21, 8),
29744 => conv_std_logic_vector(21, 8),
29745 => conv_std_logic_vector(22, 8),
29746 => conv_std_logic_vector(22, 8),
29747 => conv_std_logic_vector(23, 8),
29748 => conv_std_logic_vector(23, 8),
29749 => conv_std_logic_vector(24, 8),
29750 => conv_std_logic_vector(24, 8),
29751 => conv_std_logic_vector(24, 8),
29752 => conv_std_logic_vector(25, 8),
29753 => conv_std_logic_vector(25, 8),
29754 => conv_std_logic_vector(26, 8),
29755 => conv_std_logic_vector(26, 8),
29756 => conv_std_logic_vector(27, 8),
29757 => conv_std_logic_vector(27, 8),
29758 => conv_std_logic_vector(28, 8),
29759 => conv_std_logic_vector(28, 8),
29760 => conv_std_logic_vector(29, 8),
29761 => conv_std_logic_vector(29, 8),
29762 => conv_std_logic_vector(29, 8),
29763 => conv_std_logic_vector(30, 8),
29764 => conv_std_logic_vector(30, 8),
29765 => conv_std_logic_vector(31, 8),
29766 => conv_std_logic_vector(31, 8),
29767 => conv_std_logic_vector(32, 8),
29768 => conv_std_logic_vector(32, 8),
29769 => conv_std_logic_vector(33, 8),
29770 => conv_std_logic_vector(33, 8),
29771 => conv_std_logic_vector(33, 8),
29772 => conv_std_logic_vector(34, 8),
29773 => conv_std_logic_vector(34, 8),
29774 => conv_std_logic_vector(35, 8),
29775 => conv_std_logic_vector(35, 8),
29776 => conv_std_logic_vector(36, 8),
29777 => conv_std_logic_vector(36, 8),
29778 => conv_std_logic_vector(37, 8),
29779 => conv_std_logic_vector(37, 8),
29780 => conv_std_logic_vector(38, 8),
29781 => conv_std_logic_vector(38, 8),
29782 => conv_std_logic_vector(38, 8),
29783 => conv_std_logic_vector(39, 8),
29784 => conv_std_logic_vector(39, 8),
29785 => conv_std_logic_vector(40, 8),
29786 => conv_std_logic_vector(40, 8),
29787 => conv_std_logic_vector(41, 8),
29788 => conv_std_logic_vector(41, 8),
29789 => conv_std_logic_vector(42, 8),
29790 => conv_std_logic_vector(42, 8),
29791 => conv_std_logic_vector(43, 8),
29792 => conv_std_logic_vector(43, 8),
29793 => conv_std_logic_vector(43, 8),
29794 => conv_std_logic_vector(44, 8),
29795 => conv_std_logic_vector(44, 8),
29796 => conv_std_logic_vector(45, 8),
29797 => conv_std_logic_vector(45, 8),
29798 => conv_std_logic_vector(46, 8),
29799 => conv_std_logic_vector(46, 8),
29800 => conv_std_logic_vector(47, 8),
29801 => conv_std_logic_vector(47, 8),
29802 => conv_std_logic_vector(48, 8),
29803 => conv_std_logic_vector(48, 8),
29804 => conv_std_logic_vector(48, 8),
29805 => conv_std_logic_vector(49, 8),
29806 => conv_std_logic_vector(49, 8),
29807 => conv_std_logic_vector(50, 8),
29808 => conv_std_logic_vector(50, 8),
29809 => conv_std_logic_vector(51, 8),
29810 => conv_std_logic_vector(51, 8),
29811 => conv_std_logic_vector(52, 8),
29812 => conv_std_logic_vector(52, 8),
29813 => conv_std_logic_vector(53, 8),
29814 => conv_std_logic_vector(53, 8),
29815 => conv_std_logic_vector(53, 8),
29816 => conv_std_logic_vector(54, 8),
29817 => conv_std_logic_vector(54, 8),
29818 => conv_std_logic_vector(55, 8),
29819 => conv_std_logic_vector(55, 8),
29820 => conv_std_logic_vector(56, 8),
29821 => conv_std_logic_vector(56, 8),
29822 => conv_std_logic_vector(57, 8),
29823 => conv_std_logic_vector(57, 8),
29824 => conv_std_logic_vector(58, 8),
29825 => conv_std_logic_vector(58, 8),
29826 => conv_std_logic_vector(58, 8),
29827 => conv_std_logic_vector(59, 8),
29828 => conv_std_logic_vector(59, 8),
29829 => conv_std_logic_vector(60, 8),
29830 => conv_std_logic_vector(60, 8),
29831 => conv_std_logic_vector(61, 8),
29832 => conv_std_logic_vector(61, 8),
29833 => conv_std_logic_vector(62, 8),
29834 => conv_std_logic_vector(62, 8),
29835 => conv_std_logic_vector(62, 8),
29836 => conv_std_logic_vector(63, 8),
29837 => conv_std_logic_vector(63, 8),
29838 => conv_std_logic_vector(64, 8),
29839 => conv_std_logic_vector(64, 8),
29840 => conv_std_logic_vector(65, 8),
29841 => conv_std_logic_vector(65, 8),
29842 => conv_std_logic_vector(66, 8),
29843 => conv_std_logic_vector(66, 8),
29844 => conv_std_logic_vector(67, 8),
29845 => conv_std_logic_vector(67, 8),
29846 => conv_std_logic_vector(67, 8),
29847 => conv_std_logic_vector(68, 8),
29848 => conv_std_logic_vector(68, 8),
29849 => conv_std_logic_vector(69, 8),
29850 => conv_std_logic_vector(69, 8),
29851 => conv_std_logic_vector(70, 8),
29852 => conv_std_logic_vector(70, 8),
29853 => conv_std_logic_vector(71, 8),
29854 => conv_std_logic_vector(71, 8),
29855 => conv_std_logic_vector(72, 8),
29856 => conv_std_logic_vector(72, 8),
29857 => conv_std_logic_vector(72, 8),
29858 => conv_std_logic_vector(73, 8),
29859 => conv_std_logic_vector(73, 8),
29860 => conv_std_logic_vector(74, 8),
29861 => conv_std_logic_vector(74, 8),
29862 => conv_std_logic_vector(75, 8),
29863 => conv_std_logic_vector(75, 8),
29864 => conv_std_logic_vector(76, 8),
29865 => conv_std_logic_vector(76, 8),
29866 => conv_std_logic_vector(77, 8),
29867 => conv_std_logic_vector(77, 8),
29868 => conv_std_logic_vector(77, 8),
29869 => conv_std_logic_vector(78, 8),
29870 => conv_std_logic_vector(78, 8),
29871 => conv_std_logic_vector(79, 8),
29872 => conv_std_logic_vector(79, 8),
29873 => conv_std_logic_vector(80, 8),
29874 => conv_std_logic_vector(80, 8),
29875 => conv_std_logic_vector(81, 8),
29876 => conv_std_logic_vector(81, 8),
29877 => conv_std_logic_vector(82, 8),
29878 => conv_std_logic_vector(82, 8),
29879 => conv_std_logic_vector(82, 8),
29880 => conv_std_logic_vector(83, 8),
29881 => conv_std_logic_vector(83, 8),
29882 => conv_std_logic_vector(84, 8),
29883 => conv_std_logic_vector(84, 8),
29884 => conv_std_logic_vector(85, 8),
29885 => conv_std_logic_vector(85, 8),
29886 => conv_std_logic_vector(86, 8),
29887 => conv_std_logic_vector(86, 8),
29888 => conv_std_logic_vector(87, 8),
29889 => conv_std_logic_vector(87, 8),
29890 => conv_std_logic_vector(87, 8),
29891 => conv_std_logic_vector(88, 8),
29892 => conv_std_logic_vector(88, 8),
29893 => conv_std_logic_vector(89, 8),
29894 => conv_std_logic_vector(89, 8),
29895 => conv_std_logic_vector(90, 8),
29896 => conv_std_logic_vector(90, 8),
29897 => conv_std_logic_vector(91, 8),
29898 => conv_std_logic_vector(91, 8),
29899 => conv_std_logic_vector(91, 8),
29900 => conv_std_logic_vector(92, 8),
29901 => conv_std_logic_vector(92, 8),
29902 => conv_std_logic_vector(93, 8),
29903 => conv_std_logic_vector(93, 8),
29904 => conv_std_logic_vector(94, 8),
29905 => conv_std_logic_vector(94, 8),
29906 => conv_std_logic_vector(95, 8),
29907 => conv_std_logic_vector(95, 8),
29908 => conv_std_logic_vector(96, 8),
29909 => conv_std_logic_vector(96, 8),
29910 => conv_std_logic_vector(96, 8),
29911 => conv_std_logic_vector(97, 8),
29912 => conv_std_logic_vector(97, 8),
29913 => conv_std_logic_vector(98, 8),
29914 => conv_std_logic_vector(98, 8),
29915 => conv_std_logic_vector(99, 8),
29916 => conv_std_logic_vector(99, 8),
29917 => conv_std_logic_vector(100, 8),
29918 => conv_std_logic_vector(100, 8),
29919 => conv_std_logic_vector(101, 8),
29920 => conv_std_logic_vector(101, 8),
29921 => conv_std_logic_vector(101, 8),
29922 => conv_std_logic_vector(102, 8),
29923 => conv_std_logic_vector(102, 8),
29924 => conv_std_logic_vector(103, 8),
29925 => conv_std_logic_vector(103, 8),
29926 => conv_std_logic_vector(104, 8),
29927 => conv_std_logic_vector(104, 8),
29928 => conv_std_logic_vector(105, 8),
29929 => conv_std_logic_vector(105, 8),
29930 => conv_std_logic_vector(106, 8),
29931 => conv_std_logic_vector(106, 8),
29932 => conv_std_logic_vector(106, 8),
29933 => conv_std_logic_vector(107, 8),
29934 => conv_std_logic_vector(107, 8),
29935 => conv_std_logic_vector(108, 8),
29936 => conv_std_logic_vector(108, 8),
29937 => conv_std_logic_vector(109, 8),
29938 => conv_std_logic_vector(109, 8),
29939 => conv_std_logic_vector(110, 8),
29940 => conv_std_logic_vector(110, 8),
29941 => conv_std_logic_vector(111, 8),
29942 => conv_std_logic_vector(111, 8),
29943 => conv_std_logic_vector(111, 8),
29944 => conv_std_logic_vector(112, 8),
29945 => conv_std_logic_vector(112, 8),
29946 => conv_std_logic_vector(113, 8),
29947 => conv_std_logic_vector(113, 8),
29948 => conv_std_logic_vector(114, 8),
29949 => conv_std_logic_vector(114, 8),
29950 => conv_std_logic_vector(115, 8),
29951 => conv_std_logic_vector(115, 8),
29952 => conv_std_logic_vector(0, 8),
29953 => conv_std_logic_vector(0, 8),
29954 => conv_std_logic_vector(0, 8),
29955 => conv_std_logic_vector(1, 8),
29956 => conv_std_logic_vector(1, 8),
29957 => conv_std_logic_vector(2, 8),
29958 => conv_std_logic_vector(2, 8),
29959 => conv_std_logic_vector(3, 8),
29960 => conv_std_logic_vector(3, 8),
29961 => conv_std_logic_vector(4, 8),
29962 => conv_std_logic_vector(4, 8),
29963 => conv_std_logic_vector(5, 8),
29964 => conv_std_logic_vector(5, 8),
29965 => conv_std_logic_vector(5, 8),
29966 => conv_std_logic_vector(6, 8),
29967 => conv_std_logic_vector(6, 8),
29968 => conv_std_logic_vector(7, 8),
29969 => conv_std_logic_vector(7, 8),
29970 => conv_std_logic_vector(8, 8),
29971 => conv_std_logic_vector(8, 8),
29972 => conv_std_logic_vector(9, 8),
29973 => conv_std_logic_vector(9, 8),
29974 => conv_std_logic_vector(10, 8),
29975 => conv_std_logic_vector(10, 8),
29976 => conv_std_logic_vector(10, 8),
29977 => conv_std_logic_vector(11, 8),
29978 => conv_std_logic_vector(11, 8),
29979 => conv_std_logic_vector(12, 8),
29980 => conv_std_logic_vector(12, 8),
29981 => conv_std_logic_vector(13, 8),
29982 => conv_std_logic_vector(13, 8),
29983 => conv_std_logic_vector(14, 8),
29984 => conv_std_logic_vector(14, 8),
29985 => conv_std_logic_vector(15, 8),
29986 => conv_std_logic_vector(15, 8),
29987 => conv_std_logic_vector(15, 8),
29988 => conv_std_logic_vector(16, 8),
29989 => conv_std_logic_vector(16, 8),
29990 => conv_std_logic_vector(17, 8),
29991 => conv_std_logic_vector(17, 8),
29992 => conv_std_logic_vector(18, 8),
29993 => conv_std_logic_vector(18, 8),
29994 => conv_std_logic_vector(19, 8),
29995 => conv_std_logic_vector(19, 8),
29996 => conv_std_logic_vector(20, 8),
29997 => conv_std_logic_vector(20, 8),
29998 => conv_std_logic_vector(21, 8),
29999 => conv_std_logic_vector(21, 8),
30000 => conv_std_logic_vector(21, 8),
30001 => conv_std_logic_vector(22, 8),
30002 => conv_std_logic_vector(22, 8),
30003 => conv_std_logic_vector(23, 8),
30004 => conv_std_logic_vector(23, 8),
30005 => conv_std_logic_vector(24, 8),
30006 => conv_std_logic_vector(24, 8),
30007 => conv_std_logic_vector(25, 8),
30008 => conv_std_logic_vector(25, 8),
30009 => conv_std_logic_vector(26, 8),
30010 => conv_std_logic_vector(26, 8),
30011 => conv_std_logic_vector(26, 8),
30012 => conv_std_logic_vector(27, 8),
30013 => conv_std_logic_vector(27, 8),
30014 => conv_std_logic_vector(28, 8),
30015 => conv_std_logic_vector(28, 8),
30016 => conv_std_logic_vector(29, 8),
30017 => conv_std_logic_vector(29, 8),
30018 => conv_std_logic_vector(30, 8),
30019 => conv_std_logic_vector(30, 8),
30020 => conv_std_logic_vector(31, 8),
30021 => conv_std_logic_vector(31, 8),
30022 => conv_std_logic_vector(31, 8),
30023 => conv_std_logic_vector(32, 8),
30024 => conv_std_logic_vector(32, 8),
30025 => conv_std_logic_vector(33, 8),
30026 => conv_std_logic_vector(33, 8),
30027 => conv_std_logic_vector(34, 8),
30028 => conv_std_logic_vector(34, 8),
30029 => conv_std_logic_vector(35, 8),
30030 => conv_std_logic_vector(35, 8),
30031 => conv_std_logic_vector(36, 8),
30032 => conv_std_logic_vector(36, 8),
30033 => conv_std_logic_vector(37, 8),
30034 => conv_std_logic_vector(37, 8),
30035 => conv_std_logic_vector(37, 8),
30036 => conv_std_logic_vector(38, 8),
30037 => conv_std_logic_vector(38, 8),
30038 => conv_std_logic_vector(39, 8),
30039 => conv_std_logic_vector(39, 8),
30040 => conv_std_logic_vector(40, 8),
30041 => conv_std_logic_vector(40, 8),
30042 => conv_std_logic_vector(41, 8),
30043 => conv_std_logic_vector(41, 8),
30044 => conv_std_logic_vector(42, 8),
30045 => conv_std_logic_vector(42, 8),
30046 => conv_std_logic_vector(42, 8),
30047 => conv_std_logic_vector(43, 8),
30048 => conv_std_logic_vector(43, 8),
30049 => conv_std_logic_vector(44, 8),
30050 => conv_std_logic_vector(44, 8),
30051 => conv_std_logic_vector(45, 8),
30052 => conv_std_logic_vector(45, 8),
30053 => conv_std_logic_vector(46, 8),
30054 => conv_std_logic_vector(46, 8),
30055 => conv_std_logic_vector(47, 8),
30056 => conv_std_logic_vector(47, 8),
30057 => conv_std_logic_vector(47, 8),
30058 => conv_std_logic_vector(48, 8),
30059 => conv_std_logic_vector(48, 8),
30060 => conv_std_logic_vector(49, 8),
30061 => conv_std_logic_vector(49, 8),
30062 => conv_std_logic_vector(50, 8),
30063 => conv_std_logic_vector(50, 8),
30064 => conv_std_logic_vector(51, 8),
30065 => conv_std_logic_vector(51, 8),
30066 => conv_std_logic_vector(52, 8),
30067 => conv_std_logic_vector(52, 8),
30068 => conv_std_logic_vector(53, 8),
30069 => conv_std_logic_vector(53, 8),
30070 => conv_std_logic_vector(53, 8),
30071 => conv_std_logic_vector(54, 8),
30072 => conv_std_logic_vector(54, 8),
30073 => conv_std_logic_vector(55, 8),
30074 => conv_std_logic_vector(55, 8),
30075 => conv_std_logic_vector(56, 8),
30076 => conv_std_logic_vector(56, 8),
30077 => conv_std_logic_vector(57, 8),
30078 => conv_std_logic_vector(57, 8),
30079 => conv_std_logic_vector(58, 8),
30080 => conv_std_logic_vector(58, 8),
30081 => conv_std_logic_vector(58, 8),
30082 => conv_std_logic_vector(59, 8),
30083 => conv_std_logic_vector(59, 8),
30084 => conv_std_logic_vector(60, 8),
30085 => conv_std_logic_vector(60, 8),
30086 => conv_std_logic_vector(61, 8),
30087 => conv_std_logic_vector(61, 8),
30088 => conv_std_logic_vector(62, 8),
30089 => conv_std_logic_vector(62, 8),
30090 => conv_std_logic_vector(63, 8),
30091 => conv_std_logic_vector(63, 8),
30092 => conv_std_logic_vector(63, 8),
30093 => conv_std_logic_vector(64, 8),
30094 => conv_std_logic_vector(64, 8),
30095 => conv_std_logic_vector(65, 8),
30096 => conv_std_logic_vector(65, 8),
30097 => conv_std_logic_vector(66, 8),
30098 => conv_std_logic_vector(66, 8),
30099 => conv_std_logic_vector(67, 8),
30100 => conv_std_logic_vector(67, 8),
30101 => conv_std_logic_vector(68, 8),
30102 => conv_std_logic_vector(68, 8),
30103 => conv_std_logic_vector(69, 8),
30104 => conv_std_logic_vector(69, 8),
30105 => conv_std_logic_vector(69, 8),
30106 => conv_std_logic_vector(70, 8),
30107 => conv_std_logic_vector(70, 8),
30108 => conv_std_logic_vector(71, 8),
30109 => conv_std_logic_vector(71, 8),
30110 => conv_std_logic_vector(72, 8),
30111 => conv_std_logic_vector(72, 8),
30112 => conv_std_logic_vector(73, 8),
30113 => conv_std_logic_vector(73, 8),
30114 => conv_std_logic_vector(74, 8),
30115 => conv_std_logic_vector(74, 8),
30116 => conv_std_logic_vector(74, 8),
30117 => conv_std_logic_vector(75, 8),
30118 => conv_std_logic_vector(75, 8),
30119 => conv_std_logic_vector(76, 8),
30120 => conv_std_logic_vector(76, 8),
30121 => conv_std_logic_vector(77, 8),
30122 => conv_std_logic_vector(77, 8),
30123 => conv_std_logic_vector(78, 8),
30124 => conv_std_logic_vector(78, 8),
30125 => conv_std_logic_vector(79, 8),
30126 => conv_std_logic_vector(79, 8),
30127 => conv_std_logic_vector(79, 8),
30128 => conv_std_logic_vector(80, 8),
30129 => conv_std_logic_vector(80, 8),
30130 => conv_std_logic_vector(81, 8),
30131 => conv_std_logic_vector(81, 8),
30132 => conv_std_logic_vector(82, 8),
30133 => conv_std_logic_vector(82, 8),
30134 => conv_std_logic_vector(83, 8),
30135 => conv_std_logic_vector(83, 8),
30136 => conv_std_logic_vector(84, 8),
30137 => conv_std_logic_vector(84, 8),
30138 => conv_std_logic_vector(85, 8),
30139 => conv_std_logic_vector(85, 8),
30140 => conv_std_logic_vector(85, 8),
30141 => conv_std_logic_vector(86, 8),
30142 => conv_std_logic_vector(86, 8),
30143 => conv_std_logic_vector(87, 8),
30144 => conv_std_logic_vector(87, 8),
30145 => conv_std_logic_vector(88, 8),
30146 => conv_std_logic_vector(88, 8),
30147 => conv_std_logic_vector(89, 8),
30148 => conv_std_logic_vector(89, 8),
30149 => conv_std_logic_vector(90, 8),
30150 => conv_std_logic_vector(90, 8),
30151 => conv_std_logic_vector(90, 8),
30152 => conv_std_logic_vector(91, 8),
30153 => conv_std_logic_vector(91, 8),
30154 => conv_std_logic_vector(92, 8),
30155 => conv_std_logic_vector(92, 8),
30156 => conv_std_logic_vector(93, 8),
30157 => conv_std_logic_vector(93, 8),
30158 => conv_std_logic_vector(94, 8),
30159 => conv_std_logic_vector(94, 8),
30160 => conv_std_logic_vector(95, 8),
30161 => conv_std_logic_vector(95, 8),
30162 => conv_std_logic_vector(95, 8),
30163 => conv_std_logic_vector(96, 8),
30164 => conv_std_logic_vector(96, 8),
30165 => conv_std_logic_vector(97, 8),
30166 => conv_std_logic_vector(97, 8),
30167 => conv_std_logic_vector(98, 8),
30168 => conv_std_logic_vector(98, 8),
30169 => conv_std_logic_vector(99, 8),
30170 => conv_std_logic_vector(99, 8),
30171 => conv_std_logic_vector(100, 8),
30172 => conv_std_logic_vector(100, 8),
30173 => conv_std_logic_vector(101, 8),
30174 => conv_std_logic_vector(101, 8),
30175 => conv_std_logic_vector(101, 8),
30176 => conv_std_logic_vector(102, 8),
30177 => conv_std_logic_vector(102, 8),
30178 => conv_std_logic_vector(103, 8),
30179 => conv_std_logic_vector(103, 8),
30180 => conv_std_logic_vector(104, 8),
30181 => conv_std_logic_vector(104, 8),
30182 => conv_std_logic_vector(105, 8),
30183 => conv_std_logic_vector(105, 8),
30184 => conv_std_logic_vector(106, 8),
30185 => conv_std_logic_vector(106, 8),
30186 => conv_std_logic_vector(106, 8),
30187 => conv_std_logic_vector(107, 8),
30188 => conv_std_logic_vector(107, 8),
30189 => conv_std_logic_vector(108, 8),
30190 => conv_std_logic_vector(108, 8),
30191 => conv_std_logic_vector(109, 8),
30192 => conv_std_logic_vector(109, 8),
30193 => conv_std_logic_vector(110, 8),
30194 => conv_std_logic_vector(110, 8),
30195 => conv_std_logic_vector(111, 8),
30196 => conv_std_logic_vector(111, 8),
30197 => conv_std_logic_vector(111, 8),
30198 => conv_std_logic_vector(112, 8),
30199 => conv_std_logic_vector(112, 8),
30200 => conv_std_logic_vector(113, 8),
30201 => conv_std_logic_vector(113, 8),
30202 => conv_std_logic_vector(114, 8),
30203 => conv_std_logic_vector(114, 8),
30204 => conv_std_logic_vector(115, 8),
30205 => conv_std_logic_vector(115, 8),
30206 => conv_std_logic_vector(116, 8),
30207 => conv_std_logic_vector(116, 8),
30208 => conv_std_logic_vector(0, 8),
30209 => conv_std_logic_vector(0, 8),
30210 => conv_std_logic_vector(0, 8),
30211 => conv_std_logic_vector(1, 8),
30212 => conv_std_logic_vector(1, 8),
30213 => conv_std_logic_vector(2, 8),
30214 => conv_std_logic_vector(2, 8),
30215 => conv_std_logic_vector(3, 8),
30216 => conv_std_logic_vector(3, 8),
30217 => conv_std_logic_vector(4, 8),
30218 => conv_std_logic_vector(4, 8),
30219 => conv_std_logic_vector(5, 8),
30220 => conv_std_logic_vector(5, 8),
30221 => conv_std_logic_vector(5, 8),
30222 => conv_std_logic_vector(6, 8),
30223 => conv_std_logic_vector(6, 8),
30224 => conv_std_logic_vector(7, 8),
30225 => conv_std_logic_vector(7, 8),
30226 => conv_std_logic_vector(8, 8),
30227 => conv_std_logic_vector(8, 8),
30228 => conv_std_logic_vector(9, 8),
30229 => conv_std_logic_vector(9, 8),
30230 => conv_std_logic_vector(10, 8),
30231 => conv_std_logic_vector(10, 8),
30232 => conv_std_logic_vector(11, 8),
30233 => conv_std_logic_vector(11, 8),
30234 => conv_std_logic_vector(11, 8),
30235 => conv_std_logic_vector(12, 8),
30236 => conv_std_logic_vector(12, 8),
30237 => conv_std_logic_vector(13, 8),
30238 => conv_std_logic_vector(13, 8),
30239 => conv_std_logic_vector(14, 8),
30240 => conv_std_logic_vector(14, 8),
30241 => conv_std_logic_vector(15, 8),
30242 => conv_std_logic_vector(15, 8),
30243 => conv_std_logic_vector(16, 8),
30244 => conv_std_logic_vector(16, 8),
30245 => conv_std_logic_vector(17, 8),
30246 => conv_std_logic_vector(17, 8),
30247 => conv_std_logic_vector(17, 8),
30248 => conv_std_logic_vector(18, 8),
30249 => conv_std_logic_vector(18, 8),
30250 => conv_std_logic_vector(19, 8),
30251 => conv_std_logic_vector(19, 8),
30252 => conv_std_logic_vector(20, 8),
30253 => conv_std_logic_vector(20, 8),
30254 => conv_std_logic_vector(21, 8),
30255 => conv_std_logic_vector(21, 8),
30256 => conv_std_logic_vector(22, 8),
30257 => conv_std_logic_vector(22, 8),
30258 => conv_std_logic_vector(23, 8),
30259 => conv_std_logic_vector(23, 8),
30260 => conv_std_logic_vector(23, 8),
30261 => conv_std_logic_vector(24, 8),
30262 => conv_std_logic_vector(24, 8),
30263 => conv_std_logic_vector(25, 8),
30264 => conv_std_logic_vector(25, 8),
30265 => conv_std_logic_vector(26, 8),
30266 => conv_std_logic_vector(26, 8),
30267 => conv_std_logic_vector(27, 8),
30268 => conv_std_logic_vector(27, 8),
30269 => conv_std_logic_vector(28, 8),
30270 => conv_std_logic_vector(28, 8),
30271 => conv_std_logic_vector(29, 8),
30272 => conv_std_logic_vector(29, 8),
30273 => conv_std_logic_vector(29, 8),
30274 => conv_std_logic_vector(30, 8),
30275 => conv_std_logic_vector(30, 8),
30276 => conv_std_logic_vector(31, 8),
30277 => conv_std_logic_vector(31, 8),
30278 => conv_std_logic_vector(32, 8),
30279 => conv_std_logic_vector(32, 8),
30280 => conv_std_logic_vector(33, 8),
30281 => conv_std_logic_vector(33, 8),
30282 => conv_std_logic_vector(34, 8),
30283 => conv_std_logic_vector(34, 8),
30284 => conv_std_logic_vector(35, 8),
30285 => conv_std_logic_vector(35, 8),
30286 => conv_std_logic_vector(35, 8),
30287 => conv_std_logic_vector(36, 8),
30288 => conv_std_logic_vector(36, 8),
30289 => conv_std_logic_vector(37, 8),
30290 => conv_std_logic_vector(37, 8),
30291 => conv_std_logic_vector(38, 8),
30292 => conv_std_logic_vector(38, 8),
30293 => conv_std_logic_vector(39, 8),
30294 => conv_std_logic_vector(39, 8),
30295 => conv_std_logic_vector(40, 8),
30296 => conv_std_logic_vector(40, 8),
30297 => conv_std_logic_vector(41, 8),
30298 => conv_std_logic_vector(41, 8),
30299 => conv_std_logic_vector(41, 8),
30300 => conv_std_logic_vector(42, 8),
30301 => conv_std_logic_vector(42, 8),
30302 => conv_std_logic_vector(43, 8),
30303 => conv_std_logic_vector(43, 8),
30304 => conv_std_logic_vector(44, 8),
30305 => conv_std_logic_vector(44, 8),
30306 => conv_std_logic_vector(45, 8),
30307 => conv_std_logic_vector(45, 8),
30308 => conv_std_logic_vector(46, 8),
30309 => conv_std_logic_vector(46, 8),
30310 => conv_std_logic_vector(47, 8),
30311 => conv_std_logic_vector(47, 8),
30312 => conv_std_logic_vector(47, 8),
30313 => conv_std_logic_vector(48, 8),
30314 => conv_std_logic_vector(48, 8),
30315 => conv_std_logic_vector(49, 8),
30316 => conv_std_logic_vector(49, 8),
30317 => conv_std_logic_vector(50, 8),
30318 => conv_std_logic_vector(50, 8),
30319 => conv_std_logic_vector(51, 8),
30320 => conv_std_logic_vector(51, 8),
30321 => conv_std_logic_vector(52, 8),
30322 => conv_std_logic_vector(52, 8),
30323 => conv_std_logic_vector(53, 8),
30324 => conv_std_logic_vector(53, 8),
30325 => conv_std_logic_vector(53, 8),
30326 => conv_std_logic_vector(54, 8),
30327 => conv_std_logic_vector(54, 8),
30328 => conv_std_logic_vector(55, 8),
30329 => conv_std_logic_vector(55, 8),
30330 => conv_std_logic_vector(56, 8),
30331 => conv_std_logic_vector(56, 8),
30332 => conv_std_logic_vector(57, 8),
30333 => conv_std_logic_vector(57, 8),
30334 => conv_std_logic_vector(58, 8),
30335 => conv_std_logic_vector(58, 8),
30336 => conv_std_logic_vector(59, 8),
30337 => conv_std_logic_vector(59, 8),
30338 => conv_std_logic_vector(59, 8),
30339 => conv_std_logic_vector(60, 8),
30340 => conv_std_logic_vector(60, 8),
30341 => conv_std_logic_vector(61, 8),
30342 => conv_std_logic_vector(61, 8),
30343 => conv_std_logic_vector(62, 8),
30344 => conv_std_logic_vector(62, 8),
30345 => conv_std_logic_vector(63, 8),
30346 => conv_std_logic_vector(63, 8),
30347 => conv_std_logic_vector(64, 8),
30348 => conv_std_logic_vector(64, 8),
30349 => conv_std_logic_vector(64, 8),
30350 => conv_std_logic_vector(65, 8),
30351 => conv_std_logic_vector(65, 8),
30352 => conv_std_logic_vector(66, 8),
30353 => conv_std_logic_vector(66, 8),
30354 => conv_std_logic_vector(67, 8),
30355 => conv_std_logic_vector(67, 8),
30356 => conv_std_logic_vector(68, 8),
30357 => conv_std_logic_vector(68, 8),
30358 => conv_std_logic_vector(69, 8),
30359 => conv_std_logic_vector(69, 8),
30360 => conv_std_logic_vector(70, 8),
30361 => conv_std_logic_vector(70, 8),
30362 => conv_std_logic_vector(70, 8),
30363 => conv_std_logic_vector(71, 8),
30364 => conv_std_logic_vector(71, 8),
30365 => conv_std_logic_vector(72, 8),
30366 => conv_std_logic_vector(72, 8),
30367 => conv_std_logic_vector(73, 8),
30368 => conv_std_logic_vector(73, 8),
30369 => conv_std_logic_vector(74, 8),
30370 => conv_std_logic_vector(74, 8),
30371 => conv_std_logic_vector(75, 8),
30372 => conv_std_logic_vector(75, 8),
30373 => conv_std_logic_vector(76, 8),
30374 => conv_std_logic_vector(76, 8),
30375 => conv_std_logic_vector(76, 8),
30376 => conv_std_logic_vector(77, 8),
30377 => conv_std_logic_vector(77, 8),
30378 => conv_std_logic_vector(78, 8),
30379 => conv_std_logic_vector(78, 8),
30380 => conv_std_logic_vector(79, 8),
30381 => conv_std_logic_vector(79, 8),
30382 => conv_std_logic_vector(80, 8),
30383 => conv_std_logic_vector(80, 8),
30384 => conv_std_logic_vector(81, 8),
30385 => conv_std_logic_vector(81, 8),
30386 => conv_std_logic_vector(82, 8),
30387 => conv_std_logic_vector(82, 8),
30388 => conv_std_logic_vector(82, 8),
30389 => conv_std_logic_vector(83, 8),
30390 => conv_std_logic_vector(83, 8),
30391 => conv_std_logic_vector(84, 8),
30392 => conv_std_logic_vector(84, 8),
30393 => conv_std_logic_vector(85, 8),
30394 => conv_std_logic_vector(85, 8),
30395 => conv_std_logic_vector(86, 8),
30396 => conv_std_logic_vector(86, 8),
30397 => conv_std_logic_vector(87, 8),
30398 => conv_std_logic_vector(87, 8),
30399 => conv_std_logic_vector(88, 8),
30400 => conv_std_logic_vector(88, 8),
30401 => conv_std_logic_vector(88, 8),
30402 => conv_std_logic_vector(89, 8),
30403 => conv_std_logic_vector(89, 8),
30404 => conv_std_logic_vector(90, 8),
30405 => conv_std_logic_vector(90, 8),
30406 => conv_std_logic_vector(91, 8),
30407 => conv_std_logic_vector(91, 8),
30408 => conv_std_logic_vector(92, 8),
30409 => conv_std_logic_vector(92, 8),
30410 => conv_std_logic_vector(93, 8),
30411 => conv_std_logic_vector(93, 8),
30412 => conv_std_logic_vector(94, 8),
30413 => conv_std_logic_vector(94, 8),
30414 => conv_std_logic_vector(94, 8),
30415 => conv_std_logic_vector(95, 8),
30416 => conv_std_logic_vector(95, 8),
30417 => conv_std_logic_vector(96, 8),
30418 => conv_std_logic_vector(96, 8),
30419 => conv_std_logic_vector(97, 8),
30420 => conv_std_logic_vector(97, 8),
30421 => conv_std_logic_vector(98, 8),
30422 => conv_std_logic_vector(98, 8),
30423 => conv_std_logic_vector(99, 8),
30424 => conv_std_logic_vector(99, 8),
30425 => conv_std_logic_vector(100, 8),
30426 => conv_std_logic_vector(100, 8),
30427 => conv_std_logic_vector(100, 8),
30428 => conv_std_logic_vector(101, 8),
30429 => conv_std_logic_vector(101, 8),
30430 => conv_std_logic_vector(102, 8),
30431 => conv_std_logic_vector(102, 8),
30432 => conv_std_logic_vector(103, 8),
30433 => conv_std_logic_vector(103, 8),
30434 => conv_std_logic_vector(104, 8),
30435 => conv_std_logic_vector(104, 8),
30436 => conv_std_logic_vector(105, 8),
30437 => conv_std_logic_vector(105, 8),
30438 => conv_std_logic_vector(106, 8),
30439 => conv_std_logic_vector(106, 8),
30440 => conv_std_logic_vector(106, 8),
30441 => conv_std_logic_vector(107, 8),
30442 => conv_std_logic_vector(107, 8),
30443 => conv_std_logic_vector(108, 8),
30444 => conv_std_logic_vector(108, 8),
30445 => conv_std_logic_vector(109, 8),
30446 => conv_std_logic_vector(109, 8),
30447 => conv_std_logic_vector(110, 8),
30448 => conv_std_logic_vector(110, 8),
30449 => conv_std_logic_vector(111, 8),
30450 => conv_std_logic_vector(111, 8),
30451 => conv_std_logic_vector(112, 8),
30452 => conv_std_logic_vector(112, 8),
30453 => conv_std_logic_vector(112, 8),
30454 => conv_std_logic_vector(113, 8),
30455 => conv_std_logic_vector(113, 8),
30456 => conv_std_logic_vector(114, 8),
30457 => conv_std_logic_vector(114, 8),
30458 => conv_std_logic_vector(115, 8),
30459 => conv_std_logic_vector(115, 8),
30460 => conv_std_logic_vector(116, 8),
30461 => conv_std_logic_vector(116, 8),
30462 => conv_std_logic_vector(117, 8),
30463 => conv_std_logic_vector(117, 8),
30464 => conv_std_logic_vector(0, 8),
30465 => conv_std_logic_vector(0, 8),
30466 => conv_std_logic_vector(0, 8),
30467 => conv_std_logic_vector(1, 8),
30468 => conv_std_logic_vector(1, 8),
30469 => conv_std_logic_vector(2, 8),
30470 => conv_std_logic_vector(2, 8),
30471 => conv_std_logic_vector(3, 8),
30472 => conv_std_logic_vector(3, 8),
30473 => conv_std_logic_vector(4, 8),
30474 => conv_std_logic_vector(4, 8),
30475 => conv_std_logic_vector(5, 8),
30476 => conv_std_logic_vector(5, 8),
30477 => conv_std_logic_vector(6, 8),
30478 => conv_std_logic_vector(6, 8),
30479 => conv_std_logic_vector(6, 8),
30480 => conv_std_logic_vector(7, 8),
30481 => conv_std_logic_vector(7, 8),
30482 => conv_std_logic_vector(8, 8),
30483 => conv_std_logic_vector(8, 8),
30484 => conv_std_logic_vector(9, 8),
30485 => conv_std_logic_vector(9, 8),
30486 => conv_std_logic_vector(10, 8),
30487 => conv_std_logic_vector(10, 8),
30488 => conv_std_logic_vector(11, 8),
30489 => conv_std_logic_vector(11, 8),
30490 => conv_std_logic_vector(12, 8),
30491 => conv_std_logic_vector(12, 8),
30492 => conv_std_logic_vector(13, 8),
30493 => conv_std_logic_vector(13, 8),
30494 => conv_std_logic_vector(13, 8),
30495 => conv_std_logic_vector(14, 8),
30496 => conv_std_logic_vector(14, 8),
30497 => conv_std_logic_vector(15, 8),
30498 => conv_std_logic_vector(15, 8),
30499 => conv_std_logic_vector(16, 8),
30500 => conv_std_logic_vector(16, 8),
30501 => conv_std_logic_vector(17, 8),
30502 => conv_std_logic_vector(17, 8),
30503 => conv_std_logic_vector(18, 8),
30504 => conv_std_logic_vector(18, 8),
30505 => conv_std_logic_vector(19, 8),
30506 => conv_std_logic_vector(19, 8),
30507 => conv_std_logic_vector(19, 8),
30508 => conv_std_logic_vector(20, 8),
30509 => conv_std_logic_vector(20, 8),
30510 => conv_std_logic_vector(21, 8),
30511 => conv_std_logic_vector(21, 8),
30512 => conv_std_logic_vector(22, 8),
30513 => conv_std_logic_vector(22, 8),
30514 => conv_std_logic_vector(23, 8),
30515 => conv_std_logic_vector(23, 8),
30516 => conv_std_logic_vector(24, 8),
30517 => conv_std_logic_vector(24, 8),
30518 => conv_std_logic_vector(25, 8),
30519 => conv_std_logic_vector(25, 8),
30520 => conv_std_logic_vector(26, 8),
30521 => conv_std_logic_vector(26, 8),
30522 => conv_std_logic_vector(26, 8),
30523 => conv_std_logic_vector(27, 8),
30524 => conv_std_logic_vector(27, 8),
30525 => conv_std_logic_vector(28, 8),
30526 => conv_std_logic_vector(28, 8),
30527 => conv_std_logic_vector(29, 8),
30528 => conv_std_logic_vector(29, 8),
30529 => conv_std_logic_vector(30, 8),
30530 => conv_std_logic_vector(30, 8),
30531 => conv_std_logic_vector(31, 8),
30532 => conv_std_logic_vector(31, 8),
30533 => conv_std_logic_vector(32, 8),
30534 => conv_std_logic_vector(32, 8),
30535 => conv_std_logic_vector(33, 8),
30536 => conv_std_logic_vector(33, 8),
30537 => conv_std_logic_vector(33, 8),
30538 => conv_std_logic_vector(34, 8),
30539 => conv_std_logic_vector(34, 8),
30540 => conv_std_logic_vector(35, 8),
30541 => conv_std_logic_vector(35, 8),
30542 => conv_std_logic_vector(36, 8),
30543 => conv_std_logic_vector(36, 8),
30544 => conv_std_logic_vector(37, 8),
30545 => conv_std_logic_vector(37, 8),
30546 => conv_std_logic_vector(38, 8),
30547 => conv_std_logic_vector(38, 8),
30548 => conv_std_logic_vector(39, 8),
30549 => conv_std_logic_vector(39, 8),
30550 => conv_std_logic_vector(39, 8),
30551 => conv_std_logic_vector(40, 8),
30552 => conv_std_logic_vector(40, 8),
30553 => conv_std_logic_vector(41, 8),
30554 => conv_std_logic_vector(41, 8),
30555 => conv_std_logic_vector(42, 8),
30556 => conv_std_logic_vector(42, 8),
30557 => conv_std_logic_vector(43, 8),
30558 => conv_std_logic_vector(43, 8),
30559 => conv_std_logic_vector(44, 8),
30560 => conv_std_logic_vector(44, 8),
30561 => conv_std_logic_vector(45, 8),
30562 => conv_std_logic_vector(45, 8),
30563 => conv_std_logic_vector(46, 8),
30564 => conv_std_logic_vector(46, 8),
30565 => conv_std_logic_vector(46, 8),
30566 => conv_std_logic_vector(47, 8),
30567 => conv_std_logic_vector(47, 8),
30568 => conv_std_logic_vector(48, 8),
30569 => conv_std_logic_vector(48, 8),
30570 => conv_std_logic_vector(49, 8),
30571 => conv_std_logic_vector(49, 8),
30572 => conv_std_logic_vector(50, 8),
30573 => conv_std_logic_vector(50, 8),
30574 => conv_std_logic_vector(51, 8),
30575 => conv_std_logic_vector(51, 8),
30576 => conv_std_logic_vector(52, 8),
30577 => conv_std_logic_vector(52, 8),
30578 => conv_std_logic_vector(52, 8),
30579 => conv_std_logic_vector(53, 8),
30580 => conv_std_logic_vector(53, 8),
30581 => conv_std_logic_vector(54, 8),
30582 => conv_std_logic_vector(54, 8),
30583 => conv_std_logic_vector(55, 8),
30584 => conv_std_logic_vector(55, 8),
30585 => conv_std_logic_vector(56, 8),
30586 => conv_std_logic_vector(56, 8),
30587 => conv_std_logic_vector(57, 8),
30588 => conv_std_logic_vector(57, 8),
30589 => conv_std_logic_vector(58, 8),
30590 => conv_std_logic_vector(58, 8),
30591 => conv_std_logic_vector(59, 8),
30592 => conv_std_logic_vector(59, 8),
30593 => conv_std_logic_vector(59, 8),
30594 => conv_std_logic_vector(60, 8),
30595 => conv_std_logic_vector(60, 8),
30596 => conv_std_logic_vector(61, 8),
30597 => conv_std_logic_vector(61, 8),
30598 => conv_std_logic_vector(62, 8),
30599 => conv_std_logic_vector(62, 8),
30600 => conv_std_logic_vector(63, 8),
30601 => conv_std_logic_vector(63, 8),
30602 => conv_std_logic_vector(64, 8),
30603 => conv_std_logic_vector(64, 8),
30604 => conv_std_logic_vector(65, 8),
30605 => conv_std_logic_vector(65, 8),
30606 => conv_std_logic_vector(66, 8),
30607 => conv_std_logic_vector(66, 8),
30608 => conv_std_logic_vector(66, 8),
30609 => conv_std_logic_vector(67, 8),
30610 => conv_std_logic_vector(67, 8),
30611 => conv_std_logic_vector(68, 8),
30612 => conv_std_logic_vector(68, 8),
30613 => conv_std_logic_vector(69, 8),
30614 => conv_std_logic_vector(69, 8),
30615 => conv_std_logic_vector(70, 8),
30616 => conv_std_logic_vector(70, 8),
30617 => conv_std_logic_vector(71, 8),
30618 => conv_std_logic_vector(71, 8),
30619 => conv_std_logic_vector(72, 8),
30620 => conv_std_logic_vector(72, 8),
30621 => conv_std_logic_vector(72, 8),
30622 => conv_std_logic_vector(73, 8),
30623 => conv_std_logic_vector(73, 8),
30624 => conv_std_logic_vector(74, 8),
30625 => conv_std_logic_vector(74, 8),
30626 => conv_std_logic_vector(75, 8),
30627 => conv_std_logic_vector(75, 8),
30628 => conv_std_logic_vector(76, 8),
30629 => conv_std_logic_vector(76, 8),
30630 => conv_std_logic_vector(77, 8),
30631 => conv_std_logic_vector(77, 8),
30632 => conv_std_logic_vector(78, 8),
30633 => conv_std_logic_vector(78, 8),
30634 => conv_std_logic_vector(79, 8),
30635 => conv_std_logic_vector(79, 8),
30636 => conv_std_logic_vector(79, 8),
30637 => conv_std_logic_vector(80, 8),
30638 => conv_std_logic_vector(80, 8),
30639 => conv_std_logic_vector(81, 8),
30640 => conv_std_logic_vector(81, 8),
30641 => conv_std_logic_vector(82, 8),
30642 => conv_std_logic_vector(82, 8),
30643 => conv_std_logic_vector(83, 8),
30644 => conv_std_logic_vector(83, 8),
30645 => conv_std_logic_vector(84, 8),
30646 => conv_std_logic_vector(84, 8),
30647 => conv_std_logic_vector(85, 8),
30648 => conv_std_logic_vector(85, 8),
30649 => conv_std_logic_vector(85, 8),
30650 => conv_std_logic_vector(86, 8),
30651 => conv_std_logic_vector(86, 8),
30652 => conv_std_logic_vector(87, 8),
30653 => conv_std_logic_vector(87, 8),
30654 => conv_std_logic_vector(88, 8),
30655 => conv_std_logic_vector(88, 8),
30656 => conv_std_logic_vector(89, 8),
30657 => conv_std_logic_vector(89, 8),
30658 => conv_std_logic_vector(90, 8),
30659 => conv_std_logic_vector(90, 8),
30660 => conv_std_logic_vector(91, 8),
30661 => conv_std_logic_vector(91, 8),
30662 => conv_std_logic_vector(92, 8),
30663 => conv_std_logic_vector(92, 8),
30664 => conv_std_logic_vector(92, 8),
30665 => conv_std_logic_vector(93, 8),
30666 => conv_std_logic_vector(93, 8),
30667 => conv_std_logic_vector(94, 8),
30668 => conv_std_logic_vector(94, 8),
30669 => conv_std_logic_vector(95, 8),
30670 => conv_std_logic_vector(95, 8),
30671 => conv_std_logic_vector(96, 8),
30672 => conv_std_logic_vector(96, 8),
30673 => conv_std_logic_vector(97, 8),
30674 => conv_std_logic_vector(97, 8),
30675 => conv_std_logic_vector(98, 8),
30676 => conv_std_logic_vector(98, 8),
30677 => conv_std_logic_vector(99, 8),
30678 => conv_std_logic_vector(99, 8),
30679 => conv_std_logic_vector(99, 8),
30680 => conv_std_logic_vector(100, 8),
30681 => conv_std_logic_vector(100, 8),
30682 => conv_std_logic_vector(101, 8),
30683 => conv_std_logic_vector(101, 8),
30684 => conv_std_logic_vector(102, 8),
30685 => conv_std_logic_vector(102, 8),
30686 => conv_std_logic_vector(103, 8),
30687 => conv_std_logic_vector(103, 8),
30688 => conv_std_logic_vector(104, 8),
30689 => conv_std_logic_vector(104, 8),
30690 => conv_std_logic_vector(105, 8),
30691 => conv_std_logic_vector(105, 8),
30692 => conv_std_logic_vector(105, 8),
30693 => conv_std_logic_vector(106, 8),
30694 => conv_std_logic_vector(106, 8),
30695 => conv_std_logic_vector(107, 8),
30696 => conv_std_logic_vector(107, 8),
30697 => conv_std_logic_vector(108, 8),
30698 => conv_std_logic_vector(108, 8),
30699 => conv_std_logic_vector(109, 8),
30700 => conv_std_logic_vector(109, 8),
30701 => conv_std_logic_vector(110, 8),
30702 => conv_std_logic_vector(110, 8),
30703 => conv_std_logic_vector(111, 8),
30704 => conv_std_logic_vector(111, 8),
30705 => conv_std_logic_vector(112, 8),
30706 => conv_std_logic_vector(112, 8),
30707 => conv_std_logic_vector(112, 8),
30708 => conv_std_logic_vector(113, 8),
30709 => conv_std_logic_vector(113, 8),
30710 => conv_std_logic_vector(114, 8),
30711 => conv_std_logic_vector(114, 8),
30712 => conv_std_logic_vector(115, 8),
30713 => conv_std_logic_vector(115, 8),
30714 => conv_std_logic_vector(116, 8),
30715 => conv_std_logic_vector(116, 8),
30716 => conv_std_logic_vector(117, 8),
30717 => conv_std_logic_vector(117, 8),
30718 => conv_std_logic_vector(118, 8),
30719 => conv_std_logic_vector(118, 8),
30720 => conv_std_logic_vector(0, 8),
30721 => conv_std_logic_vector(0, 8),
30722 => conv_std_logic_vector(0, 8),
30723 => conv_std_logic_vector(1, 8),
30724 => conv_std_logic_vector(1, 8),
30725 => conv_std_logic_vector(2, 8),
30726 => conv_std_logic_vector(2, 8),
30727 => conv_std_logic_vector(3, 8),
30728 => conv_std_logic_vector(3, 8),
30729 => conv_std_logic_vector(4, 8),
30730 => conv_std_logic_vector(4, 8),
30731 => conv_std_logic_vector(5, 8),
30732 => conv_std_logic_vector(5, 8),
30733 => conv_std_logic_vector(6, 8),
30734 => conv_std_logic_vector(6, 8),
30735 => conv_std_logic_vector(7, 8),
30736 => conv_std_logic_vector(7, 8),
30737 => conv_std_logic_vector(7, 8),
30738 => conv_std_logic_vector(8, 8),
30739 => conv_std_logic_vector(8, 8),
30740 => conv_std_logic_vector(9, 8),
30741 => conv_std_logic_vector(9, 8),
30742 => conv_std_logic_vector(10, 8),
30743 => conv_std_logic_vector(10, 8),
30744 => conv_std_logic_vector(11, 8),
30745 => conv_std_logic_vector(11, 8),
30746 => conv_std_logic_vector(12, 8),
30747 => conv_std_logic_vector(12, 8),
30748 => conv_std_logic_vector(13, 8),
30749 => conv_std_logic_vector(13, 8),
30750 => conv_std_logic_vector(14, 8),
30751 => conv_std_logic_vector(14, 8),
30752 => conv_std_logic_vector(15, 8),
30753 => conv_std_logic_vector(15, 8),
30754 => conv_std_logic_vector(15, 8),
30755 => conv_std_logic_vector(16, 8),
30756 => conv_std_logic_vector(16, 8),
30757 => conv_std_logic_vector(17, 8),
30758 => conv_std_logic_vector(17, 8),
30759 => conv_std_logic_vector(18, 8),
30760 => conv_std_logic_vector(18, 8),
30761 => conv_std_logic_vector(19, 8),
30762 => conv_std_logic_vector(19, 8),
30763 => conv_std_logic_vector(20, 8),
30764 => conv_std_logic_vector(20, 8),
30765 => conv_std_logic_vector(21, 8),
30766 => conv_std_logic_vector(21, 8),
30767 => conv_std_logic_vector(22, 8),
30768 => conv_std_logic_vector(22, 8),
30769 => conv_std_logic_vector(22, 8),
30770 => conv_std_logic_vector(23, 8),
30771 => conv_std_logic_vector(23, 8),
30772 => conv_std_logic_vector(24, 8),
30773 => conv_std_logic_vector(24, 8),
30774 => conv_std_logic_vector(25, 8),
30775 => conv_std_logic_vector(25, 8),
30776 => conv_std_logic_vector(26, 8),
30777 => conv_std_logic_vector(26, 8),
30778 => conv_std_logic_vector(27, 8),
30779 => conv_std_logic_vector(27, 8),
30780 => conv_std_logic_vector(28, 8),
30781 => conv_std_logic_vector(28, 8),
30782 => conv_std_logic_vector(29, 8),
30783 => conv_std_logic_vector(29, 8),
30784 => conv_std_logic_vector(30, 8),
30785 => conv_std_logic_vector(30, 8),
30786 => conv_std_logic_vector(30, 8),
30787 => conv_std_logic_vector(31, 8),
30788 => conv_std_logic_vector(31, 8),
30789 => conv_std_logic_vector(32, 8),
30790 => conv_std_logic_vector(32, 8),
30791 => conv_std_logic_vector(33, 8),
30792 => conv_std_logic_vector(33, 8),
30793 => conv_std_logic_vector(34, 8),
30794 => conv_std_logic_vector(34, 8),
30795 => conv_std_logic_vector(35, 8),
30796 => conv_std_logic_vector(35, 8),
30797 => conv_std_logic_vector(36, 8),
30798 => conv_std_logic_vector(36, 8),
30799 => conv_std_logic_vector(37, 8),
30800 => conv_std_logic_vector(37, 8),
30801 => conv_std_logic_vector(37, 8),
30802 => conv_std_logic_vector(38, 8),
30803 => conv_std_logic_vector(38, 8),
30804 => conv_std_logic_vector(39, 8),
30805 => conv_std_logic_vector(39, 8),
30806 => conv_std_logic_vector(40, 8),
30807 => conv_std_logic_vector(40, 8),
30808 => conv_std_logic_vector(41, 8),
30809 => conv_std_logic_vector(41, 8),
30810 => conv_std_logic_vector(42, 8),
30811 => conv_std_logic_vector(42, 8),
30812 => conv_std_logic_vector(43, 8),
30813 => conv_std_logic_vector(43, 8),
30814 => conv_std_logic_vector(44, 8),
30815 => conv_std_logic_vector(44, 8),
30816 => conv_std_logic_vector(45, 8),
30817 => conv_std_logic_vector(45, 8),
30818 => conv_std_logic_vector(45, 8),
30819 => conv_std_logic_vector(46, 8),
30820 => conv_std_logic_vector(46, 8),
30821 => conv_std_logic_vector(47, 8),
30822 => conv_std_logic_vector(47, 8),
30823 => conv_std_logic_vector(48, 8),
30824 => conv_std_logic_vector(48, 8),
30825 => conv_std_logic_vector(49, 8),
30826 => conv_std_logic_vector(49, 8),
30827 => conv_std_logic_vector(50, 8),
30828 => conv_std_logic_vector(50, 8),
30829 => conv_std_logic_vector(51, 8),
30830 => conv_std_logic_vector(51, 8),
30831 => conv_std_logic_vector(52, 8),
30832 => conv_std_logic_vector(52, 8),
30833 => conv_std_logic_vector(52, 8),
30834 => conv_std_logic_vector(53, 8),
30835 => conv_std_logic_vector(53, 8),
30836 => conv_std_logic_vector(54, 8),
30837 => conv_std_logic_vector(54, 8),
30838 => conv_std_logic_vector(55, 8),
30839 => conv_std_logic_vector(55, 8),
30840 => conv_std_logic_vector(56, 8),
30841 => conv_std_logic_vector(56, 8),
30842 => conv_std_logic_vector(57, 8),
30843 => conv_std_logic_vector(57, 8),
30844 => conv_std_logic_vector(58, 8),
30845 => conv_std_logic_vector(58, 8),
30846 => conv_std_logic_vector(59, 8),
30847 => conv_std_logic_vector(59, 8),
30848 => conv_std_logic_vector(60, 8),
30849 => conv_std_logic_vector(60, 8),
30850 => conv_std_logic_vector(60, 8),
30851 => conv_std_logic_vector(61, 8),
30852 => conv_std_logic_vector(61, 8),
30853 => conv_std_logic_vector(62, 8),
30854 => conv_std_logic_vector(62, 8),
30855 => conv_std_logic_vector(63, 8),
30856 => conv_std_logic_vector(63, 8),
30857 => conv_std_logic_vector(64, 8),
30858 => conv_std_logic_vector(64, 8),
30859 => conv_std_logic_vector(65, 8),
30860 => conv_std_logic_vector(65, 8),
30861 => conv_std_logic_vector(66, 8),
30862 => conv_std_logic_vector(66, 8),
30863 => conv_std_logic_vector(67, 8),
30864 => conv_std_logic_vector(67, 8),
30865 => conv_std_logic_vector(67, 8),
30866 => conv_std_logic_vector(68, 8),
30867 => conv_std_logic_vector(68, 8),
30868 => conv_std_logic_vector(69, 8),
30869 => conv_std_logic_vector(69, 8),
30870 => conv_std_logic_vector(70, 8),
30871 => conv_std_logic_vector(70, 8),
30872 => conv_std_logic_vector(71, 8),
30873 => conv_std_logic_vector(71, 8),
30874 => conv_std_logic_vector(72, 8),
30875 => conv_std_logic_vector(72, 8),
30876 => conv_std_logic_vector(73, 8),
30877 => conv_std_logic_vector(73, 8),
30878 => conv_std_logic_vector(74, 8),
30879 => conv_std_logic_vector(74, 8),
30880 => conv_std_logic_vector(75, 8),
30881 => conv_std_logic_vector(75, 8),
30882 => conv_std_logic_vector(75, 8),
30883 => conv_std_logic_vector(76, 8),
30884 => conv_std_logic_vector(76, 8),
30885 => conv_std_logic_vector(77, 8),
30886 => conv_std_logic_vector(77, 8),
30887 => conv_std_logic_vector(78, 8),
30888 => conv_std_logic_vector(78, 8),
30889 => conv_std_logic_vector(79, 8),
30890 => conv_std_logic_vector(79, 8),
30891 => conv_std_logic_vector(80, 8),
30892 => conv_std_logic_vector(80, 8),
30893 => conv_std_logic_vector(81, 8),
30894 => conv_std_logic_vector(81, 8),
30895 => conv_std_logic_vector(82, 8),
30896 => conv_std_logic_vector(82, 8),
30897 => conv_std_logic_vector(82, 8),
30898 => conv_std_logic_vector(83, 8),
30899 => conv_std_logic_vector(83, 8),
30900 => conv_std_logic_vector(84, 8),
30901 => conv_std_logic_vector(84, 8),
30902 => conv_std_logic_vector(85, 8),
30903 => conv_std_logic_vector(85, 8),
30904 => conv_std_logic_vector(86, 8),
30905 => conv_std_logic_vector(86, 8),
30906 => conv_std_logic_vector(87, 8),
30907 => conv_std_logic_vector(87, 8),
30908 => conv_std_logic_vector(88, 8),
30909 => conv_std_logic_vector(88, 8),
30910 => conv_std_logic_vector(89, 8),
30911 => conv_std_logic_vector(89, 8),
30912 => conv_std_logic_vector(90, 8),
30913 => conv_std_logic_vector(90, 8),
30914 => conv_std_logic_vector(90, 8),
30915 => conv_std_logic_vector(91, 8),
30916 => conv_std_logic_vector(91, 8),
30917 => conv_std_logic_vector(92, 8),
30918 => conv_std_logic_vector(92, 8),
30919 => conv_std_logic_vector(93, 8),
30920 => conv_std_logic_vector(93, 8),
30921 => conv_std_logic_vector(94, 8),
30922 => conv_std_logic_vector(94, 8),
30923 => conv_std_logic_vector(95, 8),
30924 => conv_std_logic_vector(95, 8),
30925 => conv_std_logic_vector(96, 8),
30926 => conv_std_logic_vector(96, 8),
30927 => conv_std_logic_vector(97, 8),
30928 => conv_std_logic_vector(97, 8),
30929 => conv_std_logic_vector(97, 8),
30930 => conv_std_logic_vector(98, 8),
30931 => conv_std_logic_vector(98, 8),
30932 => conv_std_logic_vector(99, 8),
30933 => conv_std_logic_vector(99, 8),
30934 => conv_std_logic_vector(100, 8),
30935 => conv_std_logic_vector(100, 8),
30936 => conv_std_logic_vector(101, 8),
30937 => conv_std_logic_vector(101, 8),
30938 => conv_std_logic_vector(102, 8),
30939 => conv_std_logic_vector(102, 8),
30940 => conv_std_logic_vector(103, 8),
30941 => conv_std_logic_vector(103, 8),
30942 => conv_std_logic_vector(104, 8),
30943 => conv_std_logic_vector(104, 8),
30944 => conv_std_logic_vector(105, 8),
30945 => conv_std_logic_vector(105, 8),
30946 => conv_std_logic_vector(105, 8),
30947 => conv_std_logic_vector(106, 8),
30948 => conv_std_logic_vector(106, 8),
30949 => conv_std_logic_vector(107, 8),
30950 => conv_std_logic_vector(107, 8),
30951 => conv_std_logic_vector(108, 8),
30952 => conv_std_logic_vector(108, 8),
30953 => conv_std_logic_vector(109, 8),
30954 => conv_std_logic_vector(109, 8),
30955 => conv_std_logic_vector(110, 8),
30956 => conv_std_logic_vector(110, 8),
30957 => conv_std_logic_vector(111, 8),
30958 => conv_std_logic_vector(111, 8),
30959 => conv_std_logic_vector(112, 8),
30960 => conv_std_logic_vector(112, 8),
30961 => conv_std_logic_vector(112, 8),
30962 => conv_std_logic_vector(113, 8),
30963 => conv_std_logic_vector(113, 8),
30964 => conv_std_logic_vector(114, 8),
30965 => conv_std_logic_vector(114, 8),
30966 => conv_std_logic_vector(115, 8),
30967 => conv_std_logic_vector(115, 8),
30968 => conv_std_logic_vector(116, 8),
30969 => conv_std_logic_vector(116, 8),
30970 => conv_std_logic_vector(117, 8),
30971 => conv_std_logic_vector(117, 8),
30972 => conv_std_logic_vector(118, 8),
30973 => conv_std_logic_vector(118, 8),
30974 => conv_std_logic_vector(119, 8),
30975 => conv_std_logic_vector(119, 8),
30976 => conv_std_logic_vector(0, 8),
30977 => conv_std_logic_vector(0, 8),
30978 => conv_std_logic_vector(0, 8),
30979 => conv_std_logic_vector(1, 8),
30980 => conv_std_logic_vector(1, 8),
30981 => conv_std_logic_vector(2, 8),
30982 => conv_std_logic_vector(2, 8),
30983 => conv_std_logic_vector(3, 8),
30984 => conv_std_logic_vector(3, 8),
30985 => conv_std_logic_vector(4, 8),
30986 => conv_std_logic_vector(4, 8),
30987 => conv_std_logic_vector(5, 8),
30988 => conv_std_logic_vector(5, 8),
30989 => conv_std_logic_vector(6, 8),
30990 => conv_std_logic_vector(6, 8),
30991 => conv_std_logic_vector(7, 8),
30992 => conv_std_logic_vector(7, 8),
30993 => conv_std_logic_vector(8, 8),
30994 => conv_std_logic_vector(8, 8),
30995 => conv_std_logic_vector(8, 8),
30996 => conv_std_logic_vector(9, 8),
30997 => conv_std_logic_vector(9, 8),
30998 => conv_std_logic_vector(10, 8),
30999 => conv_std_logic_vector(10, 8),
31000 => conv_std_logic_vector(11, 8),
31001 => conv_std_logic_vector(11, 8),
31002 => conv_std_logic_vector(12, 8),
31003 => conv_std_logic_vector(12, 8),
31004 => conv_std_logic_vector(13, 8),
31005 => conv_std_logic_vector(13, 8),
31006 => conv_std_logic_vector(14, 8),
31007 => conv_std_logic_vector(14, 8),
31008 => conv_std_logic_vector(15, 8),
31009 => conv_std_logic_vector(15, 8),
31010 => conv_std_logic_vector(16, 8),
31011 => conv_std_logic_vector(16, 8),
31012 => conv_std_logic_vector(17, 8),
31013 => conv_std_logic_vector(17, 8),
31014 => conv_std_logic_vector(17, 8),
31015 => conv_std_logic_vector(18, 8),
31016 => conv_std_logic_vector(18, 8),
31017 => conv_std_logic_vector(19, 8),
31018 => conv_std_logic_vector(19, 8),
31019 => conv_std_logic_vector(20, 8),
31020 => conv_std_logic_vector(20, 8),
31021 => conv_std_logic_vector(21, 8),
31022 => conv_std_logic_vector(21, 8),
31023 => conv_std_logic_vector(22, 8),
31024 => conv_std_logic_vector(22, 8),
31025 => conv_std_logic_vector(23, 8),
31026 => conv_std_logic_vector(23, 8),
31027 => conv_std_logic_vector(24, 8),
31028 => conv_std_logic_vector(24, 8),
31029 => conv_std_logic_vector(25, 8),
31030 => conv_std_logic_vector(25, 8),
31031 => conv_std_logic_vector(25, 8),
31032 => conv_std_logic_vector(26, 8),
31033 => conv_std_logic_vector(26, 8),
31034 => conv_std_logic_vector(27, 8),
31035 => conv_std_logic_vector(27, 8),
31036 => conv_std_logic_vector(28, 8),
31037 => conv_std_logic_vector(28, 8),
31038 => conv_std_logic_vector(29, 8),
31039 => conv_std_logic_vector(29, 8),
31040 => conv_std_logic_vector(30, 8),
31041 => conv_std_logic_vector(30, 8),
31042 => conv_std_logic_vector(31, 8),
31043 => conv_std_logic_vector(31, 8),
31044 => conv_std_logic_vector(32, 8),
31045 => conv_std_logic_vector(32, 8),
31046 => conv_std_logic_vector(33, 8),
31047 => conv_std_logic_vector(33, 8),
31048 => conv_std_logic_vector(34, 8),
31049 => conv_std_logic_vector(34, 8),
31050 => conv_std_logic_vector(34, 8),
31051 => conv_std_logic_vector(35, 8),
31052 => conv_std_logic_vector(35, 8),
31053 => conv_std_logic_vector(36, 8),
31054 => conv_std_logic_vector(36, 8),
31055 => conv_std_logic_vector(37, 8),
31056 => conv_std_logic_vector(37, 8),
31057 => conv_std_logic_vector(38, 8),
31058 => conv_std_logic_vector(38, 8),
31059 => conv_std_logic_vector(39, 8),
31060 => conv_std_logic_vector(39, 8),
31061 => conv_std_logic_vector(40, 8),
31062 => conv_std_logic_vector(40, 8),
31063 => conv_std_logic_vector(41, 8),
31064 => conv_std_logic_vector(41, 8),
31065 => conv_std_logic_vector(42, 8),
31066 => conv_std_logic_vector(42, 8),
31067 => conv_std_logic_vector(43, 8),
31068 => conv_std_logic_vector(43, 8),
31069 => conv_std_logic_vector(43, 8),
31070 => conv_std_logic_vector(44, 8),
31071 => conv_std_logic_vector(44, 8),
31072 => conv_std_logic_vector(45, 8),
31073 => conv_std_logic_vector(45, 8),
31074 => conv_std_logic_vector(46, 8),
31075 => conv_std_logic_vector(46, 8),
31076 => conv_std_logic_vector(47, 8),
31077 => conv_std_logic_vector(47, 8),
31078 => conv_std_logic_vector(48, 8),
31079 => conv_std_logic_vector(48, 8),
31080 => conv_std_logic_vector(49, 8),
31081 => conv_std_logic_vector(49, 8),
31082 => conv_std_logic_vector(50, 8),
31083 => conv_std_logic_vector(50, 8),
31084 => conv_std_logic_vector(51, 8),
31085 => conv_std_logic_vector(51, 8),
31086 => conv_std_logic_vector(51, 8),
31087 => conv_std_logic_vector(52, 8),
31088 => conv_std_logic_vector(52, 8),
31089 => conv_std_logic_vector(53, 8),
31090 => conv_std_logic_vector(53, 8),
31091 => conv_std_logic_vector(54, 8),
31092 => conv_std_logic_vector(54, 8),
31093 => conv_std_logic_vector(55, 8),
31094 => conv_std_logic_vector(55, 8),
31095 => conv_std_logic_vector(56, 8),
31096 => conv_std_logic_vector(56, 8),
31097 => conv_std_logic_vector(57, 8),
31098 => conv_std_logic_vector(57, 8),
31099 => conv_std_logic_vector(58, 8),
31100 => conv_std_logic_vector(58, 8),
31101 => conv_std_logic_vector(59, 8),
31102 => conv_std_logic_vector(59, 8),
31103 => conv_std_logic_vector(60, 8),
31104 => conv_std_logic_vector(60, 8),
31105 => conv_std_logic_vector(60, 8),
31106 => conv_std_logic_vector(61, 8),
31107 => conv_std_logic_vector(61, 8),
31108 => conv_std_logic_vector(62, 8),
31109 => conv_std_logic_vector(62, 8),
31110 => conv_std_logic_vector(63, 8),
31111 => conv_std_logic_vector(63, 8),
31112 => conv_std_logic_vector(64, 8),
31113 => conv_std_logic_vector(64, 8),
31114 => conv_std_logic_vector(65, 8),
31115 => conv_std_logic_vector(65, 8),
31116 => conv_std_logic_vector(66, 8),
31117 => conv_std_logic_vector(66, 8),
31118 => conv_std_logic_vector(67, 8),
31119 => conv_std_logic_vector(67, 8),
31120 => conv_std_logic_vector(68, 8),
31121 => conv_std_logic_vector(68, 8),
31122 => conv_std_logic_vector(69, 8),
31123 => conv_std_logic_vector(69, 8),
31124 => conv_std_logic_vector(69, 8),
31125 => conv_std_logic_vector(70, 8),
31126 => conv_std_logic_vector(70, 8),
31127 => conv_std_logic_vector(71, 8),
31128 => conv_std_logic_vector(71, 8),
31129 => conv_std_logic_vector(72, 8),
31130 => conv_std_logic_vector(72, 8),
31131 => conv_std_logic_vector(73, 8),
31132 => conv_std_logic_vector(73, 8),
31133 => conv_std_logic_vector(74, 8),
31134 => conv_std_logic_vector(74, 8),
31135 => conv_std_logic_vector(75, 8),
31136 => conv_std_logic_vector(75, 8),
31137 => conv_std_logic_vector(76, 8),
31138 => conv_std_logic_vector(76, 8),
31139 => conv_std_logic_vector(77, 8),
31140 => conv_std_logic_vector(77, 8),
31141 => conv_std_logic_vector(77, 8),
31142 => conv_std_logic_vector(78, 8),
31143 => conv_std_logic_vector(78, 8),
31144 => conv_std_logic_vector(79, 8),
31145 => conv_std_logic_vector(79, 8),
31146 => conv_std_logic_vector(80, 8),
31147 => conv_std_logic_vector(80, 8),
31148 => conv_std_logic_vector(81, 8),
31149 => conv_std_logic_vector(81, 8),
31150 => conv_std_logic_vector(82, 8),
31151 => conv_std_logic_vector(82, 8),
31152 => conv_std_logic_vector(83, 8),
31153 => conv_std_logic_vector(83, 8),
31154 => conv_std_logic_vector(84, 8),
31155 => conv_std_logic_vector(84, 8),
31156 => conv_std_logic_vector(85, 8),
31157 => conv_std_logic_vector(85, 8),
31158 => conv_std_logic_vector(86, 8),
31159 => conv_std_logic_vector(86, 8),
31160 => conv_std_logic_vector(86, 8),
31161 => conv_std_logic_vector(87, 8),
31162 => conv_std_logic_vector(87, 8),
31163 => conv_std_logic_vector(88, 8),
31164 => conv_std_logic_vector(88, 8),
31165 => conv_std_logic_vector(89, 8),
31166 => conv_std_logic_vector(89, 8),
31167 => conv_std_logic_vector(90, 8),
31168 => conv_std_logic_vector(90, 8),
31169 => conv_std_logic_vector(91, 8),
31170 => conv_std_logic_vector(91, 8),
31171 => conv_std_logic_vector(92, 8),
31172 => conv_std_logic_vector(92, 8),
31173 => conv_std_logic_vector(93, 8),
31174 => conv_std_logic_vector(93, 8),
31175 => conv_std_logic_vector(94, 8),
31176 => conv_std_logic_vector(94, 8),
31177 => conv_std_logic_vector(95, 8),
31178 => conv_std_logic_vector(95, 8),
31179 => conv_std_logic_vector(95, 8),
31180 => conv_std_logic_vector(96, 8),
31181 => conv_std_logic_vector(96, 8),
31182 => conv_std_logic_vector(97, 8),
31183 => conv_std_logic_vector(97, 8),
31184 => conv_std_logic_vector(98, 8),
31185 => conv_std_logic_vector(98, 8),
31186 => conv_std_logic_vector(99, 8),
31187 => conv_std_logic_vector(99, 8),
31188 => conv_std_logic_vector(100, 8),
31189 => conv_std_logic_vector(100, 8),
31190 => conv_std_logic_vector(101, 8),
31191 => conv_std_logic_vector(101, 8),
31192 => conv_std_logic_vector(102, 8),
31193 => conv_std_logic_vector(102, 8),
31194 => conv_std_logic_vector(103, 8),
31195 => conv_std_logic_vector(103, 8),
31196 => conv_std_logic_vector(103, 8),
31197 => conv_std_logic_vector(104, 8),
31198 => conv_std_logic_vector(104, 8),
31199 => conv_std_logic_vector(105, 8),
31200 => conv_std_logic_vector(105, 8),
31201 => conv_std_logic_vector(106, 8),
31202 => conv_std_logic_vector(106, 8),
31203 => conv_std_logic_vector(107, 8),
31204 => conv_std_logic_vector(107, 8),
31205 => conv_std_logic_vector(108, 8),
31206 => conv_std_logic_vector(108, 8),
31207 => conv_std_logic_vector(109, 8),
31208 => conv_std_logic_vector(109, 8),
31209 => conv_std_logic_vector(110, 8),
31210 => conv_std_logic_vector(110, 8),
31211 => conv_std_logic_vector(111, 8),
31212 => conv_std_logic_vector(111, 8),
31213 => conv_std_logic_vector(112, 8),
31214 => conv_std_logic_vector(112, 8),
31215 => conv_std_logic_vector(112, 8),
31216 => conv_std_logic_vector(113, 8),
31217 => conv_std_logic_vector(113, 8),
31218 => conv_std_logic_vector(114, 8),
31219 => conv_std_logic_vector(114, 8),
31220 => conv_std_logic_vector(115, 8),
31221 => conv_std_logic_vector(115, 8),
31222 => conv_std_logic_vector(116, 8),
31223 => conv_std_logic_vector(116, 8),
31224 => conv_std_logic_vector(117, 8),
31225 => conv_std_logic_vector(117, 8),
31226 => conv_std_logic_vector(118, 8),
31227 => conv_std_logic_vector(118, 8),
31228 => conv_std_logic_vector(119, 8),
31229 => conv_std_logic_vector(119, 8),
31230 => conv_std_logic_vector(120, 8),
31231 => conv_std_logic_vector(120, 8),
31232 => conv_std_logic_vector(0, 8),
31233 => conv_std_logic_vector(0, 8),
31234 => conv_std_logic_vector(0, 8),
31235 => conv_std_logic_vector(1, 8),
31236 => conv_std_logic_vector(1, 8),
31237 => conv_std_logic_vector(2, 8),
31238 => conv_std_logic_vector(2, 8),
31239 => conv_std_logic_vector(3, 8),
31240 => conv_std_logic_vector(3, 8),
31241 => conv_std_logic_vector(4, 8),
31242 => conv_std_logic_vector(4, 8),
31243 => conv_std_logic_vector(5, 8),
31244 => conv_std_logic_vector(5, 8),
31245 => conv_std_logic_vector(6, 8),
31246 => conv_std_logic_vector(6, 8),
31247 => conv_std_logic_vector(7, 8),
31248 => conv_std_logic_vector(7, 8),
31249 => conv_std_logic_vector(8, 8),
31250 => conv_std_logic_vector(8, 8),
31251 => conv_std_logic_vector(9, 8),
31252 => conv_std_logic_vector(9, 8),
31253 => conv_std_logic_vector(10, 8),
31254 => conv_std_logic_vector(10, 8),
31255 => conv_std_logic_vector(10, 8),
31256 => conv_std_logic_vector(11, 8),
31257 => conv_std_logic_vector(11, 8),
31258 => conv_std_logic_vector(12, 8),
31259 => conv_std_logic_vector(12, 8),
31260 => conv_std_logic_vector(13, 8),
31261 => conv_std_logic_vector(13, 8),
31262 => conv_std_logic_vector(14, 8),
31263 => conv_std_logic_vector(14, 8),
31264 => conv_std_logic_vector(15, 8),
31265 => conv_std_logic_vector(15, 8),
31266 => conv_std_logic_vector(16, 8),
31267 => conv_std_logic_vector(16, 8),
31268 => conv_std_logic_vector(17, 8),
31269 => conv_std_logic_vector(17, 8),
31270 => conv_std_logic_vector(18, 8),
31271 => conv_std_logic_vector(18, 8),
31272 => conv_std_logic_vector(19, 8),
31273 => conv_std_logic_vector(19, 8),
31274 => conv_std_logic_vector(20, 8),
31275 => conv_std_logic_vector(20, 8),
31276 => conv_std_logic_vector(20, 8),
31277 => conv_std_logic_vector(21, 8),
31278 => conv_std_logic_vector(21, 8),
31279 => conv_std_logic_vector(22, 8),
31280 => conv_std_logic_vector(22, 8),
31281 => conv_std_logic_vector(23, 8),
31282 => conv_std_logic_vector(23, 8),
31283 => conv_std_logic_vector(24, 8),
31284 => conv_std_logic_vector(24, 8),
31285 => conv_std_logic_vector(25, 8),
31286 => conv_std_logic_vector(25, 8),
31287 => conv_std_logic_vector(26, 8),
31288 => conv_std_logic_vector(26, 8),
31289 => conv_std_logic_vector(27, 8),
31290 => conv_std_logic_vector(27, 8),
31291 => conv_std_logic_vector(28, 8),
31292 => conv_std_logic_vector(28, 8),
31293 => conv_std_logic_vector(29, 8),
31294 => conv_std_logic_vector(29, 8),
31295 => conv_std_logic_vector(30, 8),
31296 => conv_std_logic_vector(30, 8),
31297 => conv_std_logic_vector(30, 8),
31298 => conv_std_logic_vector(31, 8),
31299 => conv_std_logic_vector(31, 8),
31300 => conv_std_logic_vector(32, 8),
31301 => conv_std_logic_vector(32, 8),
31302 => conv_std_logic_vector(33, 8),
31303 => conv_std_logic_vector(33, 8),
31304 => conv_std_logic_vector(34, 8),
31305 => conv_std_logic_vector(34, 8),
31306 => conv_std_logic_vector(35, 8),
31307 => conv_std_logic_vector(35, 8),
31308 => conv_std_logic_vector(36, 8),
31309 => conv_std_logic_vector(36, 8),
31310 => conv_std_logic_vector(37, 8),
31311 => conv_std_logic_vector(37, 8),
31312 => conv_std_logic_vector(38, 8),
31313 => conv_std_logic_vector(38, 8),
31314 => conv_std_logic_vector(39, 8),
31315 => conv_std_logic_vector(39, 8),
31316 => conv_std_logic_vector(40, 8),
31317 => conv_std_logic_vector(40, 8),
31318 => conv_std_logic_vector(40, 8),
31319 => conv_std_logic_vector(41, 8),
31320 => conv_std_logic_vector(41, 8),
31321 => conv_std_logic_vector(42, 8),
31322 => conv_std_logic_vector(42, 8),
31323 => conv_std_logic_vector(43, 8),
31324 => conv_std_logic_vector(43, 8),
31325 => conv_std_logic_vector(44, 8),
31326 => conv_std_logic_vector(44, 8),
31327 => conv_std_logic_vector(45, 8),
31328 => conv_std_logic_vector(45, 8),
31329 => conv_std_logic_vector(46, 8),
31330 => conv_std_logic_vector(46, 8),
31331 => conv_std_logic_vector(47, 8),
31332 => conv_std_logic_vector(47, 8),
31333 => conv_std_logic_vector(48, 8),
31334 => conv_std_logic_vector(48, 8),
31335 => conv_std_logic_vector(49, 8),
31336 => conv_std_logic_vector(49, 8),
31337 => conv_std_logic_vector(50, 8),
31338 => conv_std_logic_vector(50, 8),
31339 => conv_std_logic_vector(50, 8),
31340 => conv_std_logic_vector(51, 8),
31341 => conv_std_logic_vector(51, 8),
31342 => conv_std_logic_vector(52, 8),
31343 => conv_std_logic_vector(52, 8),
31344 => conv_std_logic_vector(53, 8),
31345 => conv_std_logic_vector(53, 8),
31346 => conv_std_logic_vector(54, 8),
31347 => conv_std_logic_vector(54, 8),
31348 => conv_std_logic_vector(55, 8),
31349 => conv_std_logic_vector(55, 8),
31350 => conv_std_logic_vector(56, 8),
31351 => conv_std_logic_vector(56, 8),
31352 => conv_std_logic_vector(57, 8),
31353 => conv_std_logic_vector(57, 8),
31354 => conv_std_logic_vector(58, 8),
31355 => conv_std_logic_vector(58, 8),
31356 => conv_std_logic_vector(59, 8),
31357 => conv_std_logic_vector(59, 8),
31358 => conv_std_logic_vector(60, 8),
31359 => conv_std_logic_vector(60, 8),
31360 => conv_std_logic_vector(61, 8),
31361 => conv_std_logic_vector(61, 8),
31362 => conv_std_logic_vector(61, 8),
31363 => conv_std_logic_vector(62, 8),
31364 => conv_std_logic_vector(62, 8),
31365 => conv_std_logic_vector(63, 8),
31366 => conv_std_logic_vector(63, 8),
31367 => conv_std_logic_vector(64, 8),
31368 => conv_std_logic_vector(64, 8),
31369 => conv_std_logic_vector(65, 8),
31370 => conv_std_logic_vector(65, 8),
31371 => conv_std_logic_vector(66, 8),
31372 => conv_std_logic_vector(66, 8),
31373 => conv_std_logic_vector(67, 8),
31374 => conv_std_logic_vector(67, 8),
31375 => conv_std_logic_vector(68, 8),
31376 => conv_std_logic_vector(68, 8),
31377 => conv_std_logic_vector(69, 8),
31378 => conv_std_logic_vector(69, 8),
31379 => conv_std_logic_vector(70, 8),
31380 => conv_std_logic_vector(70, 8),
31381 => conv_std_logic_vector(71, 8),
31382 => conv_std_logic_vector(71, 8),
31383 => conv_std_logic_vector(71, 8),
31384 => conv_std_logic_vector(72, 8),
31385 => conv_std_logic_vector(72, 8),
31386 => conv_std_logic_vector(73, 8),
31387 => conv_std_logic_vector(73, 8),
31388 => conv_std_logic_vector(74, 8),
31389 => conv_std_logic_vector(74, 8),
31390 => conv_std_logic_vector(75, 8),
31391 => conv_std_logic_vector(75, 8),
31392 => conv_std_logic_vector(76, 8),
31393 => conv_std_logic_vector(76, 8),
31394 => conv_std_logic_vector(77, 8),
31395 => conv_std_logic_vector(77, 8),
31396 => conv_std_logic_vector(78, 8),
31397 => conv_std_logic_vector(78, 8),
31398 => conv_std_logic_vector(79, 8),
31399 => conv_std_logic_vector(79, 8),
31400 => conv_std_logic_vector(80, 8),
31401 => conv_std_logic_vector(80, 8),
31402 => conv_std_logic_vector(81, 8),
31403 => conv_std_logic_vector(81, 8),
31404 => conv_std_logic_vector(81, 8),
31405 => conv_std_logic_vector(82, 8),
31406 => conv_std_logic_vector(82, 8),
31407 => conv_std_logic_vector(83, 8),
31408 => conv_std_logic_vector(83, 8),
31409 => conv_std_logic_vector(84, 8),
31410 => conv_std_logic_vector(84, 8),
31411 => conv_std_logic_vector(85, 8),
31412 => conv_std_logic_vector(85, 8),
31413 => conv_std_logic_vector(86, 8),
31414 => conv_std_logic_vector(86, 8),
31415 => conv_std_logic_vector(87, 8),
31416 => conv_std_logic_vector(87, 8),
31417 => conv_std_logic_vector(88, 8),
31418 => conv_std_logic_vector(88, 8),
31419 => conv_std_logic_vector(89, 8),
31420 => conv_std_logic_vector(89, 8),
31421 => conv_std_logic_vector(90, 8),
31422 => conv_std_logic_vector(90, 8),
31423 => conv_std_logic_vector(91, 8),
31424 => conv_std_logic_vector(91, 8),
31425 => conv_std_logic_vector(91, 8),
31426 => conv_std_logic_vector(92, 8),
31427 => conv_std_logic_vector(92, 8),
31428 => conv_std_logic_vector(93, 8),
31429 => conv_std_logic_vector(93, 8),
31430 => conv_std_logic_vector(94, 8),
31431 => conv_std_logic_vector(94, 8),
31432 => conv_std_logic_vector(95, 8),
31433 => conv_std_logic_vector(95, 8),
31434 => conv_std_logic_vector(96, 8),
31435 => conv_std_logic_vector(96, 8),
31436 => conv_std_logic_vector(97, 8),
31437 => conv_std_logic_vector(97, 8),
31438 => conv_std_logic_vector(98, 8),
31439 => conv_std_logic_vector(98, 8),
31440 => conv_std_logic_vector(99, 8),
31441 => conv_std_logic_vector(99, 8),
31442 => conv_std_logic_vector(100, 8),
31443 => conv_std_logic_vector(100, 8),
31444 => conv_std_logic_vector(101, 8),
31445 => conv_std_logic_vector(101, 8),
31446 => conv_std_logic_vector(101, 8),
31447 => conv_std_logic_vector(102, 8),
31448 => conv_std_logic_vector(102, 8),
31449 => conv_std_logic_vector(103, 8),
31450 => conv_std_logic_vector(103, 8),
31451 => conv_std_logic_vector(104, 8),
31452 => conv_std_logic_vector(104, 8),
31453 => conv_std_logic_vector(105, 8),
31454 => conv_std_logic_vector(105, 8),
31455 => conv_std_logic_vector(106, 8),
31456 => conv_std_logic_vector(106, 8),
31457 => conv_std_logic_vector(107, 8),
31458 => conv_std_logic_vector(107, 8),
31459 => conv_std_logic_vector(108, 8),
31460 => conv_std_logic_vector(108, 8),
31461 => conv_std_logic_vector(109, 8),
31462 => conv_std_logic_vector(109, 8),
31463 => conv_std_logic_vector(110, 8),
31464 => conv_std_logic_vector(110, 8),
31465 => conv_std_logic_vector(111, 8),
31466 => conv_std_logic_vector(111, 8),
31467 => conv_std_logic_vector(111, 8),
31468 => conv_std_logic_vector(112, 8),
31469 => conv_std_logic_vector(112, 8),
31470 => conv_std_logic_vector(113, 8),
31471 => conv_std_logic_vector(113, 8),
31472 => conv_std_logic_vector(114, 8),
31473 => conv_std_logic_vector(114, 8),
31474 => conv_std_logic_vector(115, 8),
31475 => conv_std_logic_vector(115, 8),
31476 => conv_std_logic_vector(116, 8),
31477 => conv_std_logic_vector(116, 8),
31478 => conv_std_logic_vector(117, 8),
31479 => conv_std_logic_vector(117, 8),
31480 => conv_std_logic_vector(118, 8),
31481 => conv_std_logic_vector(118, 8),
31482 => conv_std_logic_vector(119, 8),
31483 => conv_std_logic_vector(119, 8),
31484 => conv_std_logic_vector(120, 8),
31485 => conv_std_logic_vector(120, 8),
31486 => conv_std_logic_vector(121, 8),
31487 => conv_std_logic_vector(121, 8),
31488 => conv_std_logic_vector(0, 8),
31489 => conv_std_logic_vector(0, 8),
31490 => conv_std_logic_vector(0, 8),
31491 => conv_std_logic_vector(1, 8),
31492 => conv_std_logic_vector(1, 8),
31493 => conv_std_logic_vector(2, 8),
31494 => conv_std_logic_vector(2, 8),
31495 => conv_std_logic_vector(3, 8),
31496 => conv_std_logic_vector(3, 8),
31497 => conv_std_logic_vector(4, 8),
31498 => conv_std_logic_vector(4, 8),
31499 => conv_std_logic_vector(5, 8),
31500 => conv_std_logic_vector(5, 8),
31501 => conv_std_logic_vector(6, 8),
31502 => conv_std_logic_vector(6, 8),
31503 => conv_std_logic_vector(7, 8),
31504 => conv_std_logic_vector(7, 8),
31505 => conv_std_logic_vector(8, 8),
31506 => conv_std_logic_vector(8, 8),
31507 => conv_std_logic_vector(9, 8),
31508 => conv_std_logic_vector(9, 8),
31509 => conv_std_logic_vector(10, 8),
31510 => conv_std_logic_vector(10, 8),
31511 => conv_std_logic_vector(11, 8),
31512 => conv_std_logic_vector(11, 8),
31513 => conv_std_logic_vector(12, 8),
31514 => conv_std_logic_vector(12, 8),
31515 => conv_std_logic_vector(12, 8),
31516 => conv_std_logic_vector(13, 8),
31517 => conv_std_logic_vector(13, 8),
31518 => conv_std_logic_vector(14, 8),
31519 => conv_std_logic_vector(14, 8),
31520 => conv_std_logic_vector(15, 8),
31521 => conv_std_logic_vector(15, 8),
31522 => conv_std_logic_vector(16, 8),
31523 => conv_std_logic_vector(16, 8),
31524 => conv_std_logic_vector(17, 8),
31525 => conv_std_logic_vector(17, 8),
31526 => conv_std_logic_vector(18, 8),
31527 => conv_std_logic_vector(18, 8),
31528 => conv_std_logic_vector(19, 8),
31529 => conv_std_logic_vector(19, 8),
31530 => conv_std_logic_vector(20, 8),
31531 => conv_std_logic_vector(20, 8),
31532 => conv_std_logic_vector(21, 8),
31533 => conv_std_logic_vector(21, 8),
31534 => conv_std_logic_vector(22, 8),
31535 => conv_std_logic_vector(22, 8),
31536 => conv_std_logic_vector(23, 8),
31537 => conv_std_logic_vector(23, 8),
31538 => conv_std_logic_vector(24, 8),
31539 => conv_std_logic_vector(24, 8),
31540 => conv_std_logic_vector(24, 8),
31541 => conv_std_logic_vector(25, 8),
31542 => conv_std_logic_vector(25, 8),
31543 => conv_std_logic_vector(26, 8),
31544 => conv_std_logic_vector(26, 8),
31545 => conv_std_logic_vector(27, 8),
31546 => conv_std_logic_vector(27, 8),
31547 => conv_std_logic_vector(28, 8),
31548 => conv_std_logic_vector(28, 8),
31549 => conv_std_logic_vector(29, 8),
31550 => conv_std_logic_vector(29, 8),
31551 => conv_std_logic_vector(30, 8),
31552 => conv_std_logic_vector(30, 8),
31553 => conv_std_logic_vector(31, 8),
31554 => conv_std_logic_vector(31, 8),
31555 => conv_std_logic_vector(32, 8),
31556 => conv_std_logic_vector(32, 8),
31557 => conv_std_logic_vector(33, 8),
31558 => conv_std_logic_vector(33, 8),
31559 => conv_std_logic_vector(34, 8),
31560 => conv_std_logic_vector(34, 8),
31561 => conv_std_logic_vector(35, 8),
31562 => conv_std_logic_vector(35, 8),
31563 => conv_std_logic_vector(36, 8),
31564 => conv_std_logic_vector(36, 8),
31565 => conv_std_logic_vector(36, 8),
31566 => conv_std_logic_vector(37, 8),
31567 => conv_std_logic_vector(37, 8),
31568 => conv_std_logic_vector(38, 8),
31569 => conv_std_logic_vector(38, 8),
31570 => conv_std_logic_vector(39, 8),
31571 => conv_std_logic_vector(39, 8),
31572 => conv_std_logic_vector(40, 8),
31573 => conv_std_logic_vector(40, 8),
31574 => conv_std_logic_vector(41, 8),
31575 => conv_std_logic_vector(41, 8),
31576 => conv_std_logic_vector(42, 8),
31577 => conv_std_logic_vector(42, 8),
31578 => conv_std_logic_vector(43, 8),
31579 => conv_std_logic_vector(43, 8),
31580 => conv_std_logic_vector(44, 8),
31581 => conv_std_logic_vector(44, 8),
31582 => conv_std_logic_vector(45, 8),
31583 => conv_std_logic_vector(45, 8),
31584 => conv_std_logic_vector(46, 8),
31585 => conv_std_logic_vector(46, 8),
31586 => conv_std_logic_vector(47, 8),
31587 => conv_std_logic_vector(47, 8),
31588 => conv_std_logic_vector(48, 8),
31589 => conv_std_logic_vector(48, 8),
31590 => conv_std_logic_vector(49, 8),
31591 => conv_std_logic_vector(49, 8),
31592 => conv_std_logic_vector(49, 8),
31593 => conv_std_logic_vector(50, 8),
31594 => conv_std_logic_vector(50, 8),
31595 => conv_std_logic_vector(51, 8),
31596 => conv_std_logic_vector(51, 8),
31597 => conv_std_logic_vector(52, 8),
31598 => conv_std_logic_vector(52, 8),
31599 => conv_std_logic_vector(53, 8),
31600 => conv_std_logic_vector(53, 8),
31601 => conv_std_logic_vector(54, 8),
31602 => conv_std_logic_vector(54, 8),
31603 => conv_std_logic_vector(55, 8),
31604 => conv_std_logic_vector(55, 8),
31605 => conv_std_logic_vector(56, 8),
31606 => conv_std_logic_vector(56, 8),
31607 => conv_std_logic_vector(57, 8),
31608 => conv_std_logic_vector(57, 8),
31609 => conv_std_logic_vector(58, 8),
31610 => conv_std_logic_vector(58, 8),
31611 => conv_std_logic_vector(59, 8),
31612 => conv_std_logic_vector(59, 8),
31613 => conv_std_logic_vector(60, 8),
31614 => conv_std_logic_vector(60, 8),
31615 => conv_std_logic_vector(61, 8),
31616 => conv_std_logic_vector(61, 8),
31617 => conv_std_logic_vector(61, 8),
31618 => conv_std_logic_vector(62, 8),
31619 => conv_std_logic_vector(62, 8),
31620 => conv_std_logic_vector(63, 8),
31621 => conv_std_logic_vector(63, 8),
31622 => conv_std_logic_vector(64, 8),
31623 => conv_std_logic_vector(64, 8),
31624 => conv_std_logic_vector(65, 8),
31625 => conv_std_logic_vector(65, 8),
31626 => conv_std_logic_vector(66, 8),
31627 => conv_std_logic_vector(66, 8),
31628 => conv_std_logic_vector(67, 8),
31629 => conv_std_logic_vector(67, 8),
31630 => conv_std_logic_vector(68, 8),
31631 => conv_std_logic_vector(68, 8),
31632 => conv_std_logic_vector(69, 8),
31633 => conv_std_logic_vector(69, 8),
31634 => conv_std_logic_vector(70, 8),
31635 => conv_std_logic_vector(70, 8),
31636 => conv_std_logic_vector(71, 8),
31637 => conv_std_logic_vector(71, 8),
31638 => conv_std_logic_vector(72, 8),
31639 => conv_std_logic_vector(72, 8),
31640 => conv_std_logic_vector(73, 8),
31641 => conv_std_logic_vector(73, 8),
31642 => conv_std_logic_vector(73, 8),
31643 => conv_std_logic_vector(74, 8),
31644 => conv_std_logic_vector(74, 8),
31645 => conv_std_logic_vector(75, 8),
31646 => conv_std_logic_vector(75, 8),
31647 => conv_std_logic_vector(76, 8),
31648 => conv_std_logic_vector(76, 8),
31649 => conv_std_logic_vector(77, 8),
31650 => conv_std_logic_vector(77, 8),
31651 => conv_std_logic_vector(78, 8),
31652 => conv_std_logic_vector(78, 8),
31653 => conv_std_logic_vector(79, 8),
31654 => conv_std_logic_vector(79, 8),
31655 => conv_std_logic_vector(80, 8),
31656 => conv_std_logic_vector(80, 8),
31657 => conv_std_logic_vector(81, 8),
31658 => conv_std_logic_vector(81, 8),
31659 => conv_std_logic_vector(82, 8),
31660 => conv_std_logic_vector(82, 8),
31661 => conv_std_logic_vector(83, 8),
31662 => conv_std_logic_vector(83, 8),
31663 => conv_std_logic_vector(84, 8),
31664 => conv_std_logic_vector(84, 8),
31665 => conv_std_logic_vector(85, 8),
31666 => conv_std_logic_vector(85, 8),
31667 => conv_std_logic_vector(86, 8),
31668 => conv_std_logic_vector(86, 8),
31669 => conv_std_logic_vector(86, 8),
31670 => conv_std_logic_vector(87, 8),
31671 => conv_std_logic_vector(87, 8),
31672 => conv_std_logic_vector(88, 8),
31673 => conv_std_logic_vector(88, 8),
31674 => conv_std_logic_vector(89, 8),
31675 => conv_std_logic_vector(89, 8),
31676 => conv_std_logic_vector(90, 8),
31677 => conv_std_logic_vector(90, 8),
31678 => conv_std_logic_vector(91, 8),
31679 => conv_std_logic_vector(91, 8),
31680 => conv_std_logic_vector(92, 8),
31681 => conv_std_logic_vector(92, 8),
31682 => conv_std_logic_vector(93, 8),
31683 => conv_std_logic_vector(93, 8),
31684 => conv_std_logic_vector(94, 8),
31685 => conv_std_logic_vector(94, 8),
31686 => conv_std_logic_vector(95, 8),
31687 => conv_std_logic_vector(95, 8),
31688 => conv_std_logic_vector(96, 8),
31689 => conv_std_logic_vector(96, 8),
31690 => conv_std_logic_vector(97, 8),
31691 => conv_std_logic_vector(97, 8),
31692 => conv_std_logic_vector(98, 8),
31693 => conv_std_logic_vector(98, 8),
31694 => conv_std_logic_vector(98, 8),
31695 => conv_std_logic_vector(99, 8),
31696 => conv_std_logic_vector(99, 8),
31697 => conv_std_logic_vector(100, 8),
31698 => conv_std_logic_vector(100, 8),
31699 => conv_std_logic_vector(101, 8),
31700 => conv_std_logic_vector(101, 8),
31701 => conv_std_logic_vector(102, 8),
31702 => conv_std_logic_vector(102, 8),
31703 => conv_std_logic_vector(103, 8),
31704 => conv_std_logic_vector(103, 8),
31705 => conv_std_logic_vector(104, 8),
31706 => conv_std_logic_vector(104, 8),
31707 => conv_std_logic_vector(105, 8),
31708 => conv_std_logic_vector(105, 8),
31709 => conv_std_logic_vector(106, 8),
31710 => conv_std_logic_vector(106, 8),
31711 => conv_std_logic_vector(107, 8),
31712 => conv_std_logic_vector(107, 8),
31713 => conv_std_logic_vector(108, 8),
31714 => conv_std_logic_vector(108, 8),
31715 => conv_std_logic_vector(109, 8),
31716 => conv_std_logic_vector(109, 8),
31717 => conv_std_logic_vector(110, 8),
31718 => conv_std_logic_vector(110, 8),
31719 => conv_std_logic_vector(110, 8),
31720 => conv_std_logic_vector(111, 8),
31721 => conv_std_logic_vector(111, 8),
31722 => conv_std_logic_vector(112, 8),
31723 => conv_std_logic_vector(112, 8),
31724 => conv_std_logic_vector(113, 8),
31725 => conv_std_logic_vector(113, 8),
31726 => conv_std_logic_vector(114, 8),
31727 => conv_std_logic_vector(114, 8),
31728 => conv_std_logic_vector(115, 8),
31729 => conv_std_logic_vector(115, 8),
31730 => conv_std_logic_vector(116, 8),
31731 => conv_std_logic_vector(116, 8),
31732 => conv_std_logic_vector(117, 8),
31733 => conv_std_logic_vector(117, 8),
31734 => conv_std_logic_vector(118, 8),
31735 => conv_std_logic_vector(118, 8),
31736 => conv_std_logic_vector(119, 8),
31737 => conv_std_logic_vector(119, 8),
31738 => conv_std_logic_vector(120, 8),
31739 => conv_std_logic_vector(120, 8),
31740 => conv_std_logic_vector(121, 8),
31741 => conv_std_logic_vector(121, 8),
31742 => conv_std_logic_vector(122, 8),
31743 => conv_std_logic_vector(122, 8),
31744 => conv_std_logic_vector(0, 8),
31745 => conv_std_logic_vector(0, 8),
31746 => conv_std_logic_vector(0, 8),
31747 => conv_std_logic_vector(1, 8),
31748 => conv_std_logic_vector(1, 8),
31749 => conv_std_logic_vector(2, 8),
31750 => conv_std_logic_vector(2, 8),
31751 => conv_std_logic_vector(3, 8),
31752 => conv_std_logic_vector(3, 8),
31753 => conv_std_logic_vector(4, 8),
31754 => conv_std_logic_vector(4, 8),
31755 => conv_std_logic_vector(5, 8),
31756 => conv_std_logic_vector(5, 8),
31757 => conv_std_logic_vector(6, 8),
31758 => conv_std_logic_vector(6, 8),
31759 => conv_std_logic_vector(7, 8),
31760 => conv_std_logic_vector(7, 8),
31761 => conv_std_logic_vector(8, 8),
31762 => conv_std_logic_vector(8, 8),
31763 => conv_std_logic_vector(9, 8),
31764 => conv_std_logic_vector(9, 8),
31765 => conv_std_logic_vector(10, 8),
31766 => conv_std_logic_vector(10, 8),
31767 => conv_std_logic_vector(11, 8),
31768 => conv_std_logic_vector(11, 8),
31769 => conv_std_logic_vector(12, 8),
31770 => conv_std_logic_vector(12, 8),
31771 => conv_std_logic_vector(13, 8),
31772 => conv_std_logic_vector(13, 8),
31773 => conv_std_logic_vector(14, 8),
31774 => conv_std_logic_vector(14, 8),
31775 => conv_std_logic_vector(15, 8),
31776 => conv_std_logic_vector(15, 8),
31777 => conv_std_logic_vector(15, 8),
31778 => conv_std_logic_vector(16, 8),
31779 => conv_std_logic_vector(16, 8),
31780 => conv_std_logic_vector(17, 8),
31781 => conv_std_logic_vector(17, 8),
31782 => conv_std_logic_vector(18, 8),
31783 => conv_std_logic_vector(18, 8),
31784 => conv_std_logic_vector(19, 8),
31785 => conv_std_logic_vector(19, 8),
31786 => conv_std_logic_vector(20, 8),
31787 => conv_std_logic_vector(20, 8),
31788 => conv_std_logic_vector(21, 8),
31789 => conv_std_logic_vector(21, 8),
31790 => conv_std_logic_vector(22, 8),
31791 => conv_std_logic_vector(22, 8),
31792 => conv_std_logic_vector(23, 8),
31793 => conv_std_logic_vector(23, 8),
31794 => conv_std_logic_vector(24, 8),
31795 => conv_std_logic_vector(24, 8),
31796 => conv_std_logic_vector(25, 8),
31797 => conv_std_logic_vector(25, 8),
31798 => conv_std_logic_vector(26, 8),
31799 => conv_std_logic_vector(26, 8),
31800 => conv_std_logic_vector(27, 8),
31801 => conv_std_logic_vector(27, 8),
31802 => conv_std_logic_vector(28, 8),
31803 => conv_std_logic_vector(28, 8),
31804 => conv_std_logic_vector(29, 8),
31805 => conv_std_logic_vector(29, 8),
31806 => conv_std_logic_vector(30, 8),
31807 => conv_std_logic_vector(30, 8),
31808 => conv_std_logic_vector(31, 8),
31809 => conv_std_logic_vector(31, 8),
31810 => conv_std_logic_vector(31, 8),
31811 => conv_std_logic_vector(32, 8),
31812 => conv_std_logic_vector(32, 8),
31813 => conv_std_logic_vector(33, 8),
31814 => conv_std_logic_vector(33, 8),
31815 => conv_std_logic_vector(34, 8),
31816 => conv_std_logic_vector(34, 8),
31817 => conv_std_logic_vector(35, 8),
31818 => conv_std_logic_vector(35, 8),
31819 => conv_std_logic_vector(36, 8),
31820 => conv_std_logic_vector(36, 8),
31821 => conv_std_logic_vector(37, 8),
31822 => conv_std_logic_vector(37, 8),
31823 => conv_std_logic_vector(38, 8),
31824 => conv_std_logic_vector(38, 8),
31825 => conv_std_logic_vector(39, 8),
31826 => conv_std_logic_vector(39, 8),
31827 => conv_std_logic_vector(40, 8),
31828 => conv_std_logic_vector(40, 8),
31829 => conv_std_logic_vector(41, 8),
31830 => conv_std_logic_vector(41, 8),
31831 => conv_std_logic_vector(42, 8),
31832 => conv_std_logic_vector(42, 8),
31833 => conv_std_logic_vector(43, 8),
31834 => conv_std_logic_vector(43, 8),
31835 => conv_std_logic_vector(44, 8),
31836 => conv_std_logic_vector(44, 8),
31837 => conv_std_logic_vector(45, 8),
31838 => conv_std_logic_vector(45, 8),
31839 => conv_std_logic_vector(46, 8),
31840 => conv_std_logic_vector(46, 8),
31841 => conv_std_logic_vector(46, 8),
31842 => conv_std_logic_vector(47, 8),
31843 => conv_std_logic_vector(47, 8),
31844 => conv_std_logic_vector(48, 8),
31845 => conv_std_logic_vector(48, 8),
31846 => conv_std_logic_vector(49, 8),
31847 => conv_std_logic_vector(49, 8),
31848 => conv_std_logic_vector(50, 8),
31849 => conv_std_logic_vector(50, 8),
31850 => conv_std_logic_vector(51, 8),
31851 => conv_std_logic_vector(51, 8),
31852 => conv_std_logic_vector(52, 8),
31853 => conv_std_logic_vector(52, 8),
31854 => conv_std_logic_vector(53, 8),
31855 => conv_std_logic_vector(53, 8),
31856 => conv_std_logic_vector(54, 8),
31857 => conv_std_logic_vector(54, 8),
31858 => conv_std_logic_vector(55, 8),
31859 => conv_std_logic_vector(55, 8),
31860 => conv_std_logic_vector(56, 8),
31861 => conv_std_logic_vector(56, 8),
31862 => conv_std_logic_vector(57, 8),
31863 => conv_std_logic_vector(57, 8),
31864 => conv_std_logic_vector(58, 8),
31865 => conv_std_logic_vector(58, 8),
31866 => conv_std_logic_vector(59, 8),
31867 => conv_std_logic_vector(59, 8),
31868 => conv_std_logic_vector(60, 8),
31869 => conv_std_logic_vector(60, 8),
31870 => conv_std_logic_vector(61, 8),
31871 => conv_std_logic_vector(61, 8),
31872 => conv_std_logic_vector(62, 8),
31873 => conv_std_logic_vector(62, 8),
31874 => conv_std_logic_vector(62, 8),
31875 => conv_std_logic_vector(63, 8),
31876 => conv_std_logic_vector(63, 8),
31877 => conv_std_logic_vector(64, 8),
31878 => conv_std_logic_vector(64, 8),
31879 => conv_std_logic_vector(65, 8),
31880 => conv_std_logic_vector(65, 8),
31881 => conv_std_logic_vector(66, 8),
31882 => conv_std_logic_vector(66, 8),
31883 => conv_std_logic_vector(67, 8),
31884 => conv_std_logic_vector(67, 8),
31885 => conv_std_logic_vector(68, 8),
31886 => conv_std_logic_vector(68, 8),
31887 => conv_std_logic_vector(69, 8),
31888 => conv_std_logic_vector(69, 8),
31889 => conv_std_logic_vector(70, 8),
31890 => conv_std_logic_vector(70, 8),
31891 => conv_std_logic_vector(71, 8),
31892 => conv_std_logic_vector(71, 8),
31893 => conv_std_logic_vector(72, 8),
31894 => conv_std_logic_vector(72, 8),
31895 => conv_std_logic_vector(73, 8),
31896 => conv_std_logic_vector(73, 8),
31897 => conv_std_logic_vector(74, 8),
31898 => conv_std_logic_vector(74, 8),
31899 => conv_std_logic_vector(75, 8),
31900 => conv_std_logic_vector(75, 8),
31901 => conv_std_logic_vector(76, 8),
31902 => conv_std_logic_vector(76, 8),
31903 => conv_std_logic_vector(77, 8),
31904 => conv_std_logic_vector(77, 8),
31905 => conv_std_logic_vector(77, 8),
31906 => conv_std_logic_vector(78, 8),
31907 => conv_std_logic_vector(78, 8),
31908 => conv_std_logic_vector(79, 8),
31909 => conv_std_logic_vector(79, 8),
31910 => conv_std_logic_vector(80, 8),
31911 => conv_std_logic_vector(80, 8),
31912 => conv_std_logic_vector(81, 8),
31913 => conv_std_logic_vector(81, 8),
31914 => conv_std_logic_vector(82, 8),
31915 => conv_std_logic_vector(82, 8),
31916 => conv_std_logic_vector(83, 8),
31917 => conv_std_logic_vector(83, 8),
31918 => conv_std_logic_vector(84, 8),
31919 => conv_std_logic_vector(84, 8),
31920 => conv_std_logic_vector(85, 8),
31921 => conv_std_logic_vector(85, 8),
31922 => conv_std_logic_vector(86, 8),
31923 => conv_std_logic_vector(86, 8),
31924 => conv_std_logic_vector(87, 8),
31925 => conv_std_logic_vector(87, 8),
31926 => conv_std_logic_vector(88, 8),
31927 => conv_std_logic_vector(88, 8),
31928 => conv_std_logic_vector(89, 8),
31929 => conv_std_logic_vector(89, 8),
31930 => conv_std_logic_vector(90, 8),
31931 => conv_std_logic_vector(90, 8),
31932 => conv_std_logic_vector(91, 8),
31933 => conv_std_logic_vector(91, 8),
31934 => conv_std_logic_vector(92, 8),
31935 => conv_std_logic_vector(92, 8),
31936 => conv_std_logic_vector(93, 8),
31937 => conv_std_logic_vector(93, 8),
31938 => conv_std_logic_vector(93, 8),
31939 => conv_std_logic_vector(94, 8),
31940 => conv_std_logic_vector(94, 8),
31941 => conv_std_logic_vector(95, 8),
31942 => conv_std_logic_vector(95, 8),
31943 => conv_std_logic_vector(96, 8),
31944 => conv_std_logic_vector(96, 8),
31945 => conv_std_logic_vector(97, 8),
31946 => conv_std_logic_vector(97, 8),
31947 => conv_std_logic_vector(98, 8),
31948 => conv_std_logic_vector(98, 8),
31949 => conv_std_logic_vector(99, 8),
31950 => conv_std_logic_vector(99, 8),
31951 => conv_std_logic_vector(100, 8),
31952 => conv_std_logic_vector(100, 8),
31953 => conv_std_logic_vector(101, 8),
31954 => conv_std_logic_vector(101, 8),
31955 => conv_std_logic_vector(102, 8),
31956 => conv_std_logic_vector(102, 8),
31957 => conv_std_logic_vector(103, 8),
31958 => conv_std_logic_vector(103, 8),
31959 => conv_std_logic_vector(104, 8),
31960 => conv_std_logic_vector(104, 8),
31961 => conv_std_logic_vector(105, 8),
31962 => conv_std_logic_vector(105, 8),
31963 => conv_std_logic_vector(106, 8),
31964 => conv_std_logic_vector(106, 8),
31965 => conv_std_logic_vector(107, 8),
31966 => conv_std_logic_vector(107, 8),
31967 => conv_std_logic_vector(108, 8),
31968 => conv_std_logic_vector(108, 8),
31969 => conv_std_logic_vector(108, 8),
31970 => conv_std_logic_vector(109, 8),
31971 => conv_std_logic_vector(109, 8),
31972 => conv_std_logic_vector(110, 8),
31973 => conv_std_logic_vector(110, 8),
31974 => conv_std_logic_vector(111, 8),
31975 => conv_std_logic_vector(111, 8),
31976 => conv_std_logic_vector(112, 8),
31977 => conv_std_logic_vector(112, 8),
31978 => conv_std_logic_vector(113, 8),
31979 => conv_std_logic_vector(113, 8),
31980 => conv_std_logic_vector(114, 8),
31981 => conv_std_logic_vector(114, 8),
31982 => conv_std_logic_vector(115, 8),
31983 => conv_std_logic_vector(115, 8),
31984 => conv_std_logic_vector(116, 8),
31985 => conv_std_logic_vector(116, 8),
31986 => conv_std_logic_vector(117, 8),
31987 => conv_std_logic_vector(117, 8),
31988 => conv_std_logic_vector(118, 8),
31989 => conv_std_logic_vector(118, 8),
31990 => conv_std_logic_vector(119, 8),
31991 => conv_std_logic_vector(119, 8),
31992 => conv_std_logic_vector(120, 8),
31993 => conv_std_logic_vector(120, 8),
31994 => conv_std_logic_vector(121, 8),
31995 => conv_std_logic_vector(121, 8),
31996 => conv_std_logic_vector(122, 8),
31997 => conv_std_logic_vector(122, 8),
31998 => conv_std_logic_vector(123, 8),
31999 => conv_std_logic_vector(123, 8),
32000 => conv_std_logic_vector(0, 8),
32001 => conv_std_logic_vector(0, 8),
32002 => conv_std_logic_vector(0, 8),
32003 => conv_std_logic_vector(1, 8),
32004 => conv_std_logic_vector(1, 8),
32005 => conv_std_logic_vector(2, 8),
32006 => conv_std_logic_vector(2, 8),
32007 => conv_std_logic_vector(3, 8),
32008 => conv_std_logic_vector(3, 8),
32009 => conv_std_logic_vector(4, 8),
32010 => conv_std_logic_vector(4, 8),
32011 => conv_std_logic_vector(5, 8),
32012 => conv_std_logic_vector(5, 8),
32013 => conv_std_logic_vector(6, 8),
32014 => conv_std_logic_vector(6, 8),
32015 => conv_std_logic_vector(7, 8),
32016 => conv_std_logic_vector(7, 8),
32017 => conv_std_logic_vector(8, 8),
32018 => conv_std_logic_vector(8, 8),
32019 => conv_std_logic_vector(9, 8),
32020 => conv_std_logic_vector(9, 8),
32021 => conv_std_logic_vector(10, 8),
32022 => conv_std_logic_vector(10, 8),
32023 => conv_std_logic_vector(11, 8),
32024 => conv_std_logic_vector(11, 8),
32025 => conv_std_logic_vector(12, 8),
32026 => conv_std_logic_vector(12, 8),
32027 => conv_std_logic_vector(13, 8),
32028 => conv_std_logic_vector(13, 8),
32029 => conv_std_logic_vector(14, 8),
32030 => conv_std_logic_vector(14, 8),
32031 => conv_std_logic_vector(15, 8),
32032 => conv_std_logic_vector(15, 8),
32033 => conv_std_logic_vector(16, 8),
32034 => conv_std_logic_vector(16, 8),
32035 => conv_std_logic_vector(17, 8),
32036 => conv_std_logic_vector(17, 8),
32037 => conv_std_logic_vector(18, 8),
32038 => conv_std_logic_vector(18, 8),
32039 => conv_std_logic_vector(19, 8),
32040 => conv_std_logic_vector(19, 8),
32041 => conv_std_logic_vector(20, 8),
32042 => conv_std_logic_vector(20, 8),
32043 => conv_std_logic_vector(20, 8),
32044 => conv_std_logic_vector(21, 8),
32045 => conv_std_logic_vector(21, 8),
32046 => conv_std_logic_vector(22, 8),
32047 => conv_std_logic_vector(22, 8),
32048 => conv_std_logic_vector(23, 8),
32049 => conv_std_logic_vector(23, 8),
32050 => conv_std_logic_vector(24, 8),
32051 => conv_std_logic_vector(24, 8),
32052 => conv_std_logic_vector(25, 8),
32053 => conv_std_logic_vector(25, 8),
32054 => conv_std_logic_vector(26, 8),
32055 => conv_std_logic_vector(26, 8),
32056 => conv_std_logic_vector(27, 8),
32057 => conv_std_logic_vector(27, 8),
32058 => conv_std_logic_vector(28, 8),
32059 => conv_std_logic_vector(28, 8),
32060 => conv_std_logic_vector(29, 8),
32061 => conv_std_logic_vector(29, 8),
32062 => conv_std_logic_vector(30, 8),
32063 => conv_std_logic_vector(30, 8),
32064 => conv_std_logic_vector(31, 8),
32065 => conv_std_logic_vector(31, 8),
32066 => conv_std_logic_vector(32, 8),
32067 => conv_std_logic_vector(32, 8),
32068 => conv_std_logic_vector(33, 8),
32069 => conv_std_logic_vector(33, 8),
32070 => conv_std_logic_vector(34, 8),
32071 => conv_std_logic_vector(34, 8),
32072 => conv_std_logic_vector(35, 8),
32073 => conv_std_logic_vector(35, 8),
32074 => conv_std_logic_vector(36, 8),
32075 => conv_std_logic_vector(36, 8),
32076 => conv_std_logic_vector(37, 8),
32077 => conv_std_logic_vector(37, 8),
32078 => conv_std_logic_vector(38, 8),
32079 => conv_std_logic_vector(38, 8),
32080 => conv_std_logic_vector(39, 8),
32081 => conv_std_logic_vector(39, 8),
32082 => conv_std_logic_vector(40, 8),
32083 => conv_std_logic_vector(40, 8),
32084 => conv_std_logic_vector(41, 8),
32085 => conv_std_logic_vector(41, 8),
32086 => conv_std_logic_vector(41, 8),
32087 => conv_std_logic_vector(42, 8),
32088 => conv_std_logic_vector(42, 8),
32089 => conv_std_logic_vector(43, 8),
32090 => conv_std_logic_vector(43, 8),
32091 => conv_std_logic_vector(44, 8),
32092 => conv_std_logic_vector(44, 8),
32093 => conv_std_logic_vector(45, 8),
32094 => conv_std_logic_vector(45, 8),
32095 => conv_std_logic_vector(46, 8),
32096 => conv_std_logic_vector(46, 8),
32097 => conv_std_logic_vector(47, 8),
32098 => conv_std_logic_vector(47, 8),
32099 => conv_std_logic_vector(48, 8),
32100 => conv_std_logic_vector(48, 8),
32101 => conv_std_logic_vector(49, 8),
32102 => conv_std_logic_vector(49, 8),
32103 => conv_std_logic_vector(50, 8),
32104 => conv_std_logic_vector(50, 8),
32105 => conv_std_logic_vector(51, 8),
32106 => conv_std_logic_vector(51, 8),
32107 => conv_std_logic_vector(52, 8),
32108 => conv_std_logic_vector(52, 8),
32109 => conv_std_logic_vector(53, 8),
32110 => conv_std_logic_vector(53, 8),
32111 => conv_std_logic_vector(54, 8),
32112 => conv_std_logic_vector(54, 8),
32113 => conv_std_logic_vector(55, 8),
32114 => conv_std_logic_vector(55, 8),
32115 => conv_std_logic_vector(56, 8),
32116 => conv_std_logic_vector(56, 8),
32117 => conv_std_logic_vector(57, 8),
32118 => conv_std_logic_vector(57, 8),
32119 => conv_std_logic_vector(58, 8),
32120 => conv_std_logic_vector(58, 8),
32121 => conv_std_logic_vector(59, 8),
32122 => conv_std_logic_vector(59, 8),
32123 => conv_std_logic_vector(60, 8),
32124 => conv_std_logic_vector(60, 8),
32125 => conv_std_logic_vector(61, 8),
32126 => conv_std_logic_vector(61, 8),
32127 => conv_std_logic_vector(62, 8),
32128 => conv_std_logic_vector(62, 8),
32129 => conv_std_logic_vector(62, 8),
32130 => conv_std_logic_vector(63, 8),
32131 => conv_std_logic_vector(63, 8),
32132 => conv_std_logic_vector(64, 8),
32133 => conv_std_logic_vector(64, 8),
32134 => conv_std_logic_vector(65, 8),
32135 => conv_std_logic_vector(65, 8),
32136 => conv_std_logic_vector(66, 8),
32137 => conv_std_logic_vector(66, 8),
32138 => conv_std_logic_vector(67, 8),
32139 => conv_std_logic_vector(67, 8),
32140 => conv_std_logic_vector(68, 8),
32141 => conv_std_logic_vector(68, 8),
32142 => conv_std_logic_vector(69, 8),
32143 => conv_std_logic_vector(69, 8),
32144 => conv_std_logic_vector(70, 8),
32145 => conv_std_logic_vector(70, 8),
32146 => conv_std_logic_vector(71, 8),
32147 => conv_std_logic_vector(71, 8),
32148 => conv_std_logic_vector(72, 8),
32149 => conv_std_logic_vector(72, 8),
32150 => conv_std_logic_vector(73, 8),
32151 => conv_std_logic_vector(73, 8),
32152 => conv_std_logic_vector(74, 8),
32153 => conv_std_logic_vector(74, 8),
32154 => conv_std_logic_vector(75, 8),
32155 => conv_std_logic_vector(75, 8),
32156 => conv_std_logic_vector(76, 8),
32157 => conv_std_logic_vector(76, 8),
32158 => conv_std_logic_vector(77, 8),
32159 => conv_std_logic_vector(77, 8),
32160 => conv_std_logic_vector(78, 8),
32161 => conv_std_logic_vector(78, 8),
32162 => conv_std_logic_vector(79, 8),
32163 => conv_std_logic_vector(79, 8),
32164 => conv_std_logic_vector(80, 8),
32165 => conv_std_logic_vector(80, 8),
32166 => conv_std_logic_vector(81, 8),
32167 => conv_std_logic_vector(81, 8),
32168 => conv_std_logic_vector(82, 8),
32169 => conv_std_logic_vector(82, 8),
32170 => conv_std_logic_vector(83, 8),
32171 => conv_std_logic_vector(83, 8),
32172 => conv_std_logic_vector(83, 8),
32173 => conv_std_logic_vector(84, 8),
32174 => conv_std_logic_vector(84, 8),
32175 => conv_std_logic_vector(85, 8),
32176 => conv_std_logic_vector(85, 8),
32177 => conv_std_logic_vector(86, 8),
32178 => conv_std_logic_vector(86, 8),
32179 => conv_std_logic_vector(87, 8),
32180 => conv_std_logic_vector(87, 8),
32181 => conv_std_logic_vector(88, 8),
32182 => conv_std_logic_vector(88, 8),
32183 => conv_std_logic_vector(89, 8),
32184 => conv_std_logic_vector(89, 8),
32185 => conv_std_logic_vector(90, 8),
32186 => conv_std_logic_vector(90, 8),
32187 => conv_std_logic_vector(91, 8),
32188 => conv_std_logic_vector(91, 8),
32189 => conv_std_logic_vector(92, 8),
32190 => conv_std_logic_vector(92, 8),
32191 => conv_std_logic_vector(93, 8),
32192 => conv_std_logic_vector(93, 8),
32193 => conv_std_logic_vector(94, 8),
32194 => conv_std_logic_vector(94, 8),
32195 => conv_std_logic_vector(95, 8),
32196 => conv_std_logic_vector(95, 8),
32197 => conv_std_logic_vector(96, 8),
32198 => conv_std_logic_vector(96, 8),
32199 => conv_std_logic_vector(97, 8),
32200 => conv_std_logic_vector(97, 8),
32201 => conv_std_logic_vector(98, 8),
32202 => conv_std_logic_vector(98, 8),
32203 => conv_std_logic_vector(99, 8),
32204 => conv_std_logic_vector(99, 8),
32205 => conv_std_logic_vector(100, 8),
32206 => conv_std_logic_vector(100, 8),
32207 => conv_std_logic_vector(101, 8),
32208 => conv_std_logic_vector(101, 8),
32209 => conv_std_logic_vector(102, 8),
32210 => conv_std_logic_vector(102, 8),
32211 => conv_std_logic_vector(103, 8),
32212 => conv_std_logic_vector(103, 8),
32213 => conv_std_logic_vector(104, 8),
32214 => conv_std_logic_vector(104, 8),
32215 => conv_std_logic_vector(104, 8),
32216 => conv_std_logic_vector(105, 8),
32217 => conv_std_logic_vector(105, 8),
32218 => conv_std_logic_vector(106, 8),
32219 => conv_std_logic_vector(106, 8),
32220 => conv_std_logic_vector(107, 8),
32221 => conv_std_logic_vector(107, 8),
32222 => conv_std_logic_vector(108, 8),
32223 => conv_std_logic_vector(108, 8),
32224 => conv_std_logic_vector(109, 8),
32225 => conv_std_logic_vector(109, 8),
32226 => conv_std_logic_vector(110, 8),
32227 => conv_std_logic_vector(110, 8),
32228 => conv_std_logic_vector(111, 8),
32229 => conv_std_logic_vector(111, 8),
32230 => conv_std_logic_vector(112, 8),
32231 => conv_std_logic_vector(112, 8),
32232 => conv_std_logic_vector(113, 8),
32233 => conv_std_logic_vector(113, 8),
32234 => conv_std_logic_vector(114, 8),
32235 => conv_std_logic_vector(114, 8),
32236 => conv_std_logic_vector(115, 8),
32237 => conv_std_logic_vector(115, 8),
32238 => conv_std_logic_vector(116, 8),
32239 => conv_std_logic_vector(116, 8),
32240 => conv_std_logic_vector(117, 8),
32241 => conv_std_logic_vector(117, 8),
32242 => conv_std_logic_vector(118, 8),
32243 => conv_std_logic_vector(118, 8),
32244 => conv_std_logic_vector(119, 8),
32245 => conv_std_logic_vector(119, 8),
32246 => conv_std_logic_vector(120, 8),
32247 => conv_std_logic_vector(120, 8),
32248 => conv_std_logic_vector(121, 8),
32249 => conv_std_logic_vector(121, 8),
32250 => conv_std_logic_vector(122, 8),
32251 => conv_std_logic_vector(122, 8),
32252 => conv_std_logic_vector(123, 8),
32253 => conv_std_logic_vector(123, 8),
32254 => conv_std_logic_vector(124, 8),
32255 => conv_std_logic_vector(124, 8),
32256 => conv_std_logic_vector(0, 8),
32257 => conv_std_logic_vector(0, 8),
32258 => conv_std_logic_vector(0, 8),
32259 => conv_std_logic_vector(1, 8),
32260 => conv_std_logic_vector(1, 8),
32261 => conv_std_logic_vector(2, 8),
32262 => conv_std_logic_vector(2, 8),
32263 => conv_std_logic_vector(3, 8),
32264 => conv_std_logic_vector(3, 8),
32265 => conv_std_logic_vector(4, 8),
32266 => conv_std_logic_vector(4, 8),
32267 => conv_std_logic_vector(5, 8),
32268 => conv_std_logic_vector(5, 8),
32269 => conv_std_logic_vector(6, 8),
32270 => conv_std_logic_vector(6, 8),
32271 => conv_std_logic_vector(7, 8),
32272 => conv_std_logic_vector(7, 8),
32273 => conv_std_logic_vector(8, 8),
32274 => conv_std_logic_vector(8, 8),
32275 => conv_std_logic_vector(9, 8),
32276 => conv_std_logic_vector(9, 8),
32277 => conv_std_logic_vector(10, 8),
32278 => conv_std_logic_vector(10, 8),
32279 => conv_std_logic_vector(11, 8),
32280 => conv_std_logic_vector(11, 8),
32281 => conv_std_logic_vector(12, 8),
32282 => conv_std_logic_vector(12, 8),
32283 => conv_std_logic_vector(13, 8),
32284 => conv_std_logic_vector(13, 8),
32285 => conv_std_logic_vector(14, 8),
32286 => conv_std_logic_vector(14, 8),
32287 => conv_std_logic_vector(15, 8),
32288 => conv_std_logic_vector(15, 8),
32289 => conv_std_logic_vector(16, 8),
32290 => conv_std_logic_vector(16, 8),
32291 => conv_std_logic_vector(17, 8),
32292 => conv_std_logic_vector(17, 8),
32293 => conv_std_logic_vector(18, 8),
32294 => conv_std_logic_vector(18, 8),
32295 => conv_std_logic_vector(19, 8),
32296 => conv_std_logic_vector(19, 8),
32297 => conv_std_logic_vector(20, 8),
32298 => conv_std_logic_vector(20, 8),
32299 => conv_std_logic_vector(21, 8),
32300 => conv_std_logic_vector(21, 8),
32301 => conv_std_logic_vector(22, 8),
32302 => conv_std_logic_vector(22, 8),
32303 => conv_std_logic_vector(23, 8),
32304 => conv_std_logic_vector(23, 8),
32305 => conv_std_logic_vector(24, 8),
32306 => conv_std_logic_vector(24, 8),
32307 => conv_std_logic_vector(25, 8),
32308 => conv_std_logic_vector(25, 8),
32309 => conv_std_logic_vector(26, 8),
32310 => conv_std_logic_vector(26, 8),
32311 => conv_std_logic_vector(27, 8),
32312 => conv_std_logic_vector(27, 8),
32313 => conv_std_logic_vector(28, 8),
32314 => conv_std_logic_vector(28, 8),
32315 => conv_std_logic_vector(29, 8),
32316 => conv_std_logic_vector(29, 8),
32317 => conv_std_logic_vector(30, 8),
32318 => conv_std_logic_vector(30, 8),
32319 => conv_std_logic_vector(31, 8),
32320 => conv_std_logic_vector(31, 8),
32321 => conv_std_logic_vector(31, 8),
32322 => conv_std_logic_vector(32, 8),
32323 => conv_std_logic_vector(32, 8),
32324 => conv_std_logic_vector(33, 8),
32325 => conv_std_logic_vector(33, 8),
32326 => conv_std_logic_vector(34, 8),
32327 => conv_std_logic_vector(34, 8),
32328 => conv_std_logic_vector(35, 8),
32329 => conv_std_logic_vector(35, 8),
32330 => conv_std_logic_vector(36, 8),
32331 => conv_std_logic_vector(36, 8),
32332 => conv_std_logic_vector(37, 8),
32333 => conv_std_logic_vector(37, 8),
32334 => conv_std_logic_vector(38, 8),
32335 => conv_std_logic_vector(38, 8),
32336 => conv_std_logic_vector(39, 8),
32337 => conv_std_logic_vector(39, 8),
32338 => conv_std_logic_vector(40, 8),
32339 => conv_std_logic_vector(40, 8),
32340 => conv_std_logic_vector(41, 8),
32341 => conv_std_logic_vector(41, 8),
32342 => conv_std_logic_vector(42, 8),
32343 => conv_std_logic_vector(42, 8),
32344 => conv_std_logic_vector(43, 8),
32345 => conv_std_logic_vector(43, 8),
32346 => conv_std_logic_vector(44, 8),
32347 => conv_std_logic_vector(44, 8),
32348 => conv_std_logic_vector(45, 8),
32349 => conv_std_logic_vector(45, 8),
32350 => conv_std_logic_vector(46, 8),
32351 => conv_std_logic_vector(46, 8),
32352 => conv_std_logic_vector(47, 8),
32353 => conv_std_logic_vector(47, 8),
32354 => conv_std_logic_vector(48, 8),
32355 => conv_std_logic_vector(48, 8),
32356 => conv_std_logic_vector(49, 8),
32357 => conv_std_logic_vector(49, 8),
32358 => conv_std_logic_vector(50, 8),
32359 => conv_std_logic_vector(50, 8),
32360 => conv_std_logic_vector(51, 8),
32361 => conv_std_logic_vector(51, 8),
32362 => conv_std_logic_vector(52, 8),
32363 => conv_std_logic_vector(52, 8),
32364 => conv_std_logic_vector(53, 8),
32365 => conv_std_logic_vector(53, 8),
32366 => conv_std_logic_vector(54, 8),
32367 => conv_std_logic_vector(54, 8),
32368 => conv_std_logic_vector(55, 8),
32369 => conv_std_logic_vector(55, 8),
32370 => conv_std_logic_vector(56, 8),
32371 => conv_std_logic_vector(56, 8),
32372 => conv_std_logic_vector(57, 8),
32373 => conv_std_logic_vector(57, 8),
32374 => conv_std_logic_vector(58, 8),
32375 => conv_std_logic_vector(58, 8),
32376 => conv_std_logic_vector(59, 8),
32377 => conv_std_logic_vector(59, 8),
32378 => conv_std_logic_vector(60, 8),
32379 => conv_std_logic_vector(60, 8),
32380 => conv_std_logic_vector(61, 8),
32381 => conv_std_logic_vector(61, 8),
32382 => conv_std_logic_vector(62, 8),
32383 => conv_std_logic_vector(62, 8),
32384 => conv_std_logic_vector(63, 8),
32385 => conv_std_logic_vector(63, 8),
32386 => conv_std_logic_vector(63, 8),
32387 => conv_std_logic_vector(64, 8),
32388 => conv_std_logic_vector(64, 8),
32389 => conv_std_logic_vector(65, 8),
32390 => conv_std_logic_vector(65, 8),
32391 => conv_std_logic_vector(66, 8),
32392 => conv_std_logic_vector(66, 8),
32393 => conv_std_logic_vector(67, 8),
32394 => conv_std_logic_vector(67, 8),
32395 => conv_std_logic_vector(68, 8),
32396 => conv_std_logic_vector(68, 8),
32397 => conv_std_logic_vector(69, 8),
32398 => conv_std_logic_vector(69, 8),
32399 => conv_std_logic_vector(70, 8),
32400 => conv_std_logic_vector(70, 8),
32401 => conv_std_logic_vector(71, 8),
32402 => conv_std_logic_vector(71, 8),
32403 => conv_std_logic_vector(72, 8),
32404 => conv_std_logic_vector(72, 8),
32405 => conv_std_logic_vector(73, 8),
32406 => conv_std_logic_vector(73, 8),
32407 => conv_std_logic_vector(74, 8),
32408 => conv_std_logic_vector(74, 8),
32409 => conv_std_logic_vector(75, 8),
32410 => conv_std_logic_vector(75, 8),
32411 => conv_std_logic_vector(76, 8),
32412 => conv_std_logic_vector(76, 8),
32413 => conv_std_logic_vector(77, 8),
32414 => conv_std_logic_vector(77, 8),
32415 => conv_std_logic_vector(78, 8),
32416 => conv_std_logic_vector(78, 8),
32417 => conv_std_logic_vector(79, 8),
32418 => conv_std_logic_vector(79, 8),
32419 => conv_std_logic_vector(80, 8),
32420 => conv_std_logic_vector(80, 8),
32421 => conv_std_logic_vector(81, 8),
32422 => conv_std_logic_vector(81, 8),
32423 => conv_std_logic_vector(82, 8),
32424 => conv_std_logic_vector(82, 8),
32425 => conv_std_logic_vector(83, 8),
32426 => conv_std_logic_vector(83, 8),
32427 => conv_std_logic_vector(84, 8),
32428 => conv_std_logic_vector(84, 8),
32429 => conv_std_logic_vector(85, 8),
32430 => conv_std_logic_vector(85, 8),
32431 => conv_std_logic_vector(86, 8),
32432 => conv_std_logic_vector(86, 8),
32433 => conv_std_logic_vector(87, 8),
32434 => conv_std_logic_vector(87, 8),
32435 => conv_std_logic_vector(88, 8),
32436 => conv_std_logic_vector(88, 8),
32437 => conv_std_logic_vector(89, 8),
32438 => conv_std_logic_vector(89, 8),
32439 => conv_std_logic_vector(90, 8),
32440 => conv_std_logic_vector(90, 8),
32441 => conv_std_logic_vector(91, 8),
32442 => conv_std_logic_vector(91, 8),
32443 => conv_std_logic_vector(92, 8),
32444 => conv_std_logic_vector(92, 8),
32445 => conv_std_logic_vector(93, 8),
32446 => conv_std_logic_vector(93, 8),
32447 => conv_std_logic_vector(94, 8),
32448 => conv_std_logic_vector(94, 8),
32449 => conv_std_logic_vector(94, 8),
32450 => conv_std_logic_vector(95, 8),
32451 => conv_std_logic_vector(95, 8),
32452 => conv_std_logic_vector(96, 8),
32453 => conv_std_logic_vector(96, 8),
32454 => conv_std_logic_vector(97, 8),
32455 => conv_std_logic_vector(97, 8),
32456 => conv_std_logic_vector(98, 8),
32457 => conv_std_logic_vector(98, 8),
32458 => conv_std_logic_vector(99, 8),
32459 => conv_std_logic_vector(99, 8),
32460 => conv_std_logic_vector(100, 8),
32461 => conv_std_logic_vector(100, 8),
32462 => conv_std_logic_vector(101, 8),
32463 => conv_std_logic_vector(101, 8),
32464 => conv_std_logic_vector(102, 8),
32465 => conv_std_logic_vector(102, 8),
32466 => conv_std_logic_vector(103, 8),
32467 => conv_std_logic_vector(103, 8),
32468 => conv_std_logic_vector(104, 8),
32469 => conv_std_logic_vector(104, 8),
32470 => conv_std_logic_vector(105, 8),
32471 => conv_std_logic_vector(105, 8),
32472 => conv_std_logic_vector(106, 8),
32473 => conv_std_logic_vector(106, 8),
32474 => conv_std_logic_vector(107, 8),
32475 => conv_std_logic_vector(107, 8),
32476 => conv_std_logic_vector(108, 8),
32477 => conv_std_logic_vector(108, 8),
32478 => conv_std_logic_vector(109, 8),
32479 => conv_std_logic_vector(109, 8),
32480 => conv_std_logic_vector(110, 8),
32481 => conv_std_logic_vector(110, 8),
32482 => conv_std_logic_vector(111, 8),
32483 => conv_std_logic_vector(111, 8),
32484 => conv_std_logic_vector(112, 8),
32485 => conv_std_logic_vector(112, 8),
32486 => conv_std_logic_vector(113, 8),
32487 => conv_std_logic_vector(113, 8),
32488 => conv_std_logic_vector(114, 8),
32489 => conv_std_logic_vector(114, 8),
32490 => conv_std_logic_vector(115, 8),
32491 => conv_std_logic_vector(115, 8),
32492 => conv_std_logic_vector(116, 8),
32493 => conv_std_logic_vector(116, 8),
32494 => conv_std_logic_vector(117, 8),
32495 => conv_std_logic_vector(117, 8),
32496 => conv_std_logic_vector(118, 8),
32497 => conv_std_logic_vector(118, 8),
32498 => conv_std_logic_vector(119, 8),
32499 => conv_std_logic_vector(119, 8),
32500 => conv_std_logic_vector(120, 8),
32501 => conv_std_logic_vector(120, 8),
32502 => conv_std_logic_vector(121, 8),
32503 => conv_std_logic_vector(121, 8),
32504 => conv_std_logic_vector(122, 8),
32505 => conv_std_logic_vector(122, 8),
32506 => conv_std_logic_vector(123, 8),
32507 => conv_std_logic_vector(123, 8),
32508 => conv_std_logic_vector(124, 8),
32509 => conv_std_logic_vector(124, 8),
32510 => conv_std_logic_vector(125, 8),
32511 => conv_std_logic_vector(125, 8),
32512 => conv_std_logic_vector(0, 8),
32513 => conv_std_logic_vector(0, 8),
32514 => conv_std_logic_vector(0, 8),
32515 => conv_std_logic_vector(1, 8),
32516 => conv_std_logic_vector(1, 8),
32517 => conv_std_logic_vector(2, 8),
32518 => conv_std_logic_vector(2, 8),
32519 => conv_std_logic_vector(3, 8),
32520 => conv_std_logic_vector(3, 8),
32521 => conv_std_logic_vector(4, 8),
32522 => conv_std_logic_vector(4, 8),
32523 => conv_std_logic_vector(5, 8),
32524 => conv_std_logic_vector(5, 8),
32525 => conv_std_logic_vector(6, 8),
32526 => conv_std_logic_vector(6, 8),
32527 => conv_std_logic_vector(7, 8),
32528 => conv_std_logic_vector(7, 8),
32529 => conv_std_logic_vector(8, 8),
32530 => conv_std_logic_vector(8, 8),
32531 => conv_std_logic_vector(9, 8),
32532 => conv_std_logic_vector(9, 8),
32533 => conv_std_logic_vector(10, 8),
32534 => conv_std_logic_vector(10, 8),
32535 => conv_std_logic_vector(11, 8),
32536 => conv_std_logic_vector(11, 8),
32537 => conv_std_logic_vector(12, 8),
32538 => conv_std_logic_vector(12, 8),
32539 => conv_std_logic_vector(13, 8),
32540 => conv_std_logic_vector(13, 8),
32541 => conv_std_logic_vector(14, 8),
32542 => conv_std_logic_vector(14, 8),
32543 => conv_std_logic_vector(15, 8),
32544 => conv_std_logic_vector(15, 8),
32545 => conv_std_logic_vector(16, 8),
32546 => conv_std_logic_vector(16, 8),
32547 => conv_std_logic_vector(17, 8),
32548 => conv_std_logic_vector(17, 8),
32549 => conv_std_logic_vector(18, 8),
32550 => conv_std_logic_vector(18, 8),
32551 => conv_std_logic_vector(19, 8),
32552 => conv_std_logic_vector(19, 8),
32553 => conv_std_logic_vector(20, 8),
32554 => conv_std_logic_vector(20, 8),
32555 => conv_std_logic_vector(21, 8),
32556 => conv_std_logic_vector(21, 8),
32557 => conv_std_logic_vector(22, 8),
32558 => conv_std_logic_vector(22, 8),
32559 => conv_std_logic_vector(23, 8),
32560 => conv_std_logic_vector(23, 8),
32561 => conv_std_logic_vector(24, 8),
32562 => conv_std_logic_vector(24, 8),
32563 => conv_std_logic_vector(25, 8),
32564 => conv_std_logic_vector(25, 8),
32565 => conv_std_logic_vector(26, 8),
32566 => conv_std_logic_vector(26, 8),
32567 => conv_std_logic_vector(27, 8),
32568 => conv_std_logic_vector(27, 8),
32569 => conv_std_logic_vector(28, 8),
32570 => conv_std_logic_vector(28, 8),
32571 => conv_std_logic_vector(29, 8),
32572 => conv_std_logic_vector(29, 8),
32573 => conv_std_logic_vector(30, 8),
32574 => conv_std_logic_vector(30, 8),
32575 => conv_std_logic_vector(31, 8),
32576 => conv_std_logic_vector(31, 8),
32577 => conv_std_logic_vector(32, 8),
32578 => conv_std_logic_vector(32, 8),
32579 => conv_std_logic_vector(33, 8),
32580 => conv_std_logic_vector(33, 8),
32581 => conv_std_logic_vector(34, 8),
32582 => conv_std_logic_vector(34, 8),
32583 => conv_std_logic_vector(35, 8),
32584 => conv_std_logic_vector(35, 8),
32585 => conv_std_logic_vector(36, 8),
32586 => conv_std_logic_vector(36, 8),
32587 => conv_std_logic_vector(37, 8),
32588 => conv_std_logic_vector(37, 8),
32589 => conv_std_logic_vector(38, 8),
32590 => conv_std_logic_vector(38, 8),
32591 => conv_std_logic_vector(39, 8),
32592 => conv_std_logic_vector(39, 8),
32593 => conv_std_logic_vector(40, 8),
32594 => conv_std_logic_vector(40, 8),
32595 => conv_std_logic_vector(41, 8),
32596 => conv_std_logic_vector(41, 8),
32597 => conv_std_logic_vector(42, 8),
32598 => conv_std_logic_vector(42, 8),
32599 => conv_std_logic_vector(43, 8),
32600 => conv_std_logic_vector(43, 8),
32601 => conv_std_logic_vector(44, 8),
32602 => conv_std_logic_vector(44, 8),
32603 => conv_std_logic_vector(45, 8),
32604 => conv_std_logic_vector(45, 8),
32605 => conv_std_logic_vector(46, 8),
32606 => conv_std_logic_vector(46, 8),
32607 => conv_std_logic_vector(47, 8),
32608 => conv_std_logic_vector(47, 8),
32609 => conv_std_logic_vector(48, 8),
32610 => conv_std_logic_vector(48, 8),
32611 => conv_std_logic_vector(49, 8),
32612 => conv_std_logic_vector(49, 8),
32613 => conv_std_logic_vector(50, 8),
32614 => conv_std_logic_vector(50, 8),
32615 => conv_std_logic_vector(51, 8),
32616 => conv_std_logic_vector(51, 8),
32617 => conv_std_logic_vector(52, 8),
32618 => conv_std_logic_vector(52, 8),
32619 => conv_std_logic_vector(53, 8),
32620 => conv_std_logic_vector(53, 8),
32621 => conv_std_logic_vector(54, 8),
32622 => conv_std_logic_vector(54, 8),
32623 => conv_std_logic_vector(55, 8),
32624 => conv_std_logic_vector(55, 8),
32625 => conv_std_logic_vector(56, 8),
32626 => conv_std_logic_vector(56, 8),
32627 => conv_std_logic_vector(57, 8),
32628 => conv_std_logic_vector(57, 8),
32629 => conv_std_logic_vector(58, 8),
32630 => conv_std_logic_vector(58, 8),
32631 => conv_std_logic_vector(59, 8),
32632 => conv_std_logic_vector(59, 8),
32633 => conv_std_logic_vector(60, 8),
32634 => conv_std_logic_vector(60, 8),
32635 => conv_std_logic_vector(61, 8),
32636 => conv_std_logic_vector(61, 8),
32637 => conv_std_logic_vector(62, 8),
32638 => conv_std_logic_vector(62, 8),
32639 => conv_std_logic_vector(63, 8),
32640 => conv_std_logic_vector(63, 8),
32641 => conv_std_logic_vector(63, 8),
32642 => conv_std_logic_vector(64, 8),
32643 => conv_std_logic_vector(64, 8),
32644 => conv_std_logic_vector(65, 8),
32645 => conv_std_logic_vector(65, 8),
32646 => conv_std_logic_vector(66, 8),
32647 => conv_std_logic_vector(66, 8),
32648 => conv_std_logic_vector(67, 8),
32649 => conv_std_logic_vector(67, 8),
32650 => conv_std_logic_vector(68, 8),
32651 => conv_std_logic_vector(68, 8),
32652 => conv_std_logic_vector(69, 8),
32653 => conv_std_logic_vector(69, 8),
32654 => conv_std_logic_vector(70, 8),
32655 => conv_std_logic_vector(70, 8),
32656 => conv_std_logic_vector(71, 8),
32657 => conv_std_logic_vector(71, 8),
32658 => conv_std_logic_vector(72, 8),
32659 => conv_std_logic_vector(72, 8),
32660 => conv_std_logic_vector(73, 8),
32661 => conv_std_logic_vector(73, 8),
32662 => conv_std_logic_vector(74, 8),
32663 => conv_std_logic_vector(74, 8),
32664 => conv_std_logic_vector(75, 8),
32665 => conv_std_logic_vector(75, 8),
32666 => conv_std_logic_vector(76, 8),
32667 => conv_std_logic_vector(76, 8),
32668 => conv_std_logic_vector(77, 8),
32669 => conv_std_logic_vector(77, 8),
32670 => conv_std_logic_vector(78, 8),
32671 => conv_std_logic_vector(78, 8),
32672 => conv_std_logic_vector(79, 8),
32673 => conv_std_logic_vector(79, 8),
32674 => conv_std_logic_vector(80, 8),
32675 => conv_std_logic_vector(80, 8),
32676 => conv_std_logic_vector(81, 8),
32677 => conv_std_logic_vector(81, 8),
32678 => conv_std_logic_vector(82, 8),
32679 => conv_std_logic_vector(82, 8),
32680 => conv_std_logic_vector(83, 8),
32681 => conv_std_logic_vector(83, 8),
32682 => conv_std_logic_vector(84, 8),
32683 => conv_std_logic_vector(84, 8),
32684 => conv_std_logic_vector(85, 8),
32685 => conv_std_logic_vector(85, 8),
32686 => conv_std_logic_vector(86, 8),
32687 => conv_std_logic_vector(86, 8),
32688 => conv_std_logic_vector(87, 8),
32689 => conv_std_logic_vector(87, 8),
32690 => conv_std_logic_vector(88, 8),
32691 => conv_std_logic_vector(88, 8),
32692 => conv_std_logic_vector(89, 8),
32693 => conv_std_logic_vector(89, 8),
32694 => conv_std_logic_vector(90, 8),
32695 => conv_std_logic_vector(90, 8),
32696 => conv_std_logic_vector(91, 8),
32697 => conv_std_logic_vector(91, 8),
32698 => conv_std_logic_vector(92, 8),
32699 => conv_std_logic_vector(92, 8),
32700 => conv_std_logic_vector(93, 8),
32701 => conv_std_logic_vector(93, 8),
32702 => conv_std_logic_vector(94, 8),
32703 => conv_std_logic_vector(94, 8),
32704 => conv_std_logic_vector(95, 8),
32705 => conv_std_logic_vector(95, 8),
32706 => conv_std_logic_vector(96, 8),
32707 => conv_std_logic_vector(96, 8),
32708 => conv_std_logic_vector(97, 8),
32709 => conv_std_logic_vector(97, 8),
32710 => conv_std_logic_vector(98, 8),
32711 => conv_std_logic_vector(98, 8),
32712 => conv_std_logic_vector(99, 8),
32713 => conv_std_logic_vector(99, 8),
32714 => conv_std_logic_vector(100, 8),
32715 => conv_std_logic_vector(100, 8),
32716 => conv_std_logic_vector(101, 8),
32717 => conv_std_logic_vector(101, 8),
32718 => conv_std_logic_vector(102, 8),
32719 => conv_std_logic_vector(102, 8),
32720 => conv_std_logic_vector(103, 8),
32721 => conv_std_logic_vector(103, 8),
32722 => conv_std_logic_vector(104, 8),
32723 => conv_std_logic_vector(104, 8),
32724 => conv_std_logic_vector(105, 8),
32725 => conv_std_logic_vector(105, 8),
32726 => conv_std_logic_vector(106, 8),
32727 => conv_std_logic_vector(106, 8),
32728 => conv_std_logic_vector(107, 8),
32729 => conv_std_logic_vector(107, 8),
32730 => conv_std_logic_vector(108, 8),
32731 => conv_std_logic_vector(108, 8),
32732 => conv_std_logic_vector(109, 8),
32733 => conv_std_logic_vector(109, 8),
32734 => conv_std_logic_vector(110, 8),
32735 => conv_std_logic_vector(110, 8),
32736 => conv_std_logic_vector(111, 8),
32737 => conv_std_logic_vector(111, 8),
32738 => conv_std_logic_vector(112, 8),
32739 => conv_std_logic_vector(112, 8),
32740 => conv_std_logic_vector(113, 8),
32741 => conv_std_logic_vector(113, 8),
32742 => conv_std_logic_vector(114, 8),
32743 => conv_std_logic_vector(114, 8),
32744 => conv_std_logic_vector(115, 8),
32745 => conv_std_logic_vector(115, 8),
32746 => conv_std_logic_vector(116, 8),
32747 => conv_std_logic_vector(116, 8),
32748 => conv_std_logic_vector(117, 8),
32749 => conv_std_logic_vector(117, 8),
32750 => conv_std_logic_vector(118, 8),
32751 => conv_std_logic_vector(118, 8),
32752 => conv_std_logic_vector(119, 8),
32753 => conv_std_logic_vector(119, 8),
32754 => conv_std_logic_vector(120, 8),
32755 => conv_std_logic_vector(120, 8),
32756 => conv_std_logic_vector(121, 8),
32757 => conv_std_logic_vector(121, 8),
32758 => conv_std_logic_vector(122, 8),
32759 => conv_std_logic_vector(122, 8),
32760 => conv_std_logic_vector(123, 8),
32761 => conv_std_logic_vector(123, 8),
32762 => conv_std_logic_vector(124, 8),
32763 => conv_std_logic_vector(124, 8),
32764 => conv_std_logic_vector(125, 8),
32765 => conv_std_logic_vector(125, 8),
32766 => conv_std_logic_vector(126, 8),
32767 => conv_std_logic_vector(126, 8),
32768 => conv_std_logic_vector(0, 8),
32769 => conv_std_logic_vector(0, 8),
32770 => conv_std_logic_vector(1, 8),
32771 => conv_std_logic_vector(1, 8),
32772 => conv_std_logic_vector(2, 8),
32773 => conv_std_logic_vector(2, 8),
32774 => conv_std_logic_vector(3, 8),
32775 => conv_std_logic_vector(3, 8),
32776 => conv_std_logic_vector(4, 8),
32777 => conv_std_logic_vector(4, 8),
32778 => conv_std_logic_vector(5, 8),
32779 => conv_std_logic_vector(5, 8),
32780 => conv_std_logic_vector(6, 8),
32781 => conv_std_logic_vector(6, 8),
32782 => conv_std_logic_vector(7, 8),
32783 => conv_std_logic_vector(7, 8),
32784 => conv_std_logic_vector(8, 8),
32785 => conv_std_logic_vector(8, 8),
32786 => conv_std_logic_vector(9, 8),
32787 => conv_std_logic_vector(9, 8),
32788 => conv_std_logic_vector(10, 8),
32789 => conv_std_logic_vector(10, 8),
32790 => conv_std_logic_vector(11, 8),
32791 => conv_std_logic_vector(11, 8),
32792 => conv_std_logic_vector(12, 8),
32793 => conv_std_logic_vector(12, 8),
32794 => conv_std_logic_vector(13, 8),
32795 => conv_std_logic_vector(13, 8),
32796 => conv_std_logic_vector(14, 8),
32797 => conv_std_logic_vector(14, 8),
32798 => conv_std_logic_vector(15, 8),
32799 => conv_std_logic_vector(15, 8),
32800 => conv_std_logic_vector(16, 8),
32801 => conv_std_logic_vector(16, 8),
32802 => conv_std_logic_vector(17, 8),
32803 => conv_std_logic_vector(17, 8),
32804 => conv_std_logic_vector(18, 8),
32805 => conv_std_logic_vector(18, 8),
32806 => conv_std_logic_vector(19, 8),
32807 => conv_std_logic_vector(19, 8),
32808 => conv_std_logic_vector(20, 8),
32809 => conv_std_logic_vector(20, 8),
32810 => conv_std_logic_vector(21, 8),
32811 => conv_std_logic_vector(21, 8),
32812 => conv_std_logic_vector(22, 8),
32813 => conv_std_logic_vector(22, 8),
32814 => conv_std_logic_vector(23, 8),
32815 => conv_std_logic_vector(23, 8),
32816 => conv_std_logic_vector(24, 8),
32817 => conv_std_logic_vector(24, 8),
32818 => conv_std_logic_vector(25, 8),
32819 => conv_std_logic_vector(25, 8),
32820 => conv_std_logic_vector(26, 8),
32821 => conv_std_logic_vector(26, 8),
32822 => conv_std_logic_vector(27, 8),
32823 => conv_std_logic_vector(27, 8),
32824 => conv_std_logic_vector(28, 8),
32825 => conv_std_logic_vector(28, 8),
32826 => conv_std_logic_vector(29, 8),
32827 => conv_std_logic_vector(29, 8),
32828 => conv_std_logic_vector(30, 8),
32829 => conv_std_logic_vector(30, 8),
32830 => conv_std_logic_vector(31, 8),
32831 => conv_std_logic_vector(31, 8),
32832 => conv_std_logic_vector(32, 8),
32833 => conv_std_logic_vector(32, 8),
32834 => conv_std_logic_vector(33, 8),
32835 => conv_std_logic_vector(33, 8),
32836 => conv_std_logic_vector(34, 8),
32837 => conv_std_logic_vector(34, 8),
32838 => conv_std_logic_vector(35, 8),
32839 => conv_std_logic_vector(35, 8),
32840 => conv_std_logic_vector(36, 8),
32841 => conv_std_logic_vector(36, 8),
32842 => conv_std_logic_vector(37, 8),
32843 => conv_std_logic_vector(37, 8),
32844 => conv_std_logic_vector(38, 8),
32845 => conv_std_logic_vector(38, 8),
32846 => conv_std_logic_vector(39, 8),
32847 => conv_std_logic_vector(39, 8),
32848 => conv_std_logic_vector(40, 8),
32849 => conv_std_logic_vector(40, 8),
32850 => conv_std_logic_vector(41, 8),
32851 => conv_std_logic_vector(41, 8),
32852 => conv_std_logic_vector(42, 8),
32853 => conv_std_logic_vector(42, 8),
32854 => conv_std_logic_vector(43, 8),
32855 => conv_std_logic_vector(43, 8),
32856 => conv_std_logic_vector(44, 8),
32857 => conv_std_logic_vector(44, 8),
32858 => conv_std_logic_vector(45, 8),
32859 => conv_std_logic_vector(45, 8),
32860 => conv_std_logic_vector(46, 8),
32861 => conv_std_logic_vector(46, 8),
32862 => conv_std_logic_vector(47, 8),
32863 => conv_std_logic_vector(47, 8),
32864 => conv_std_logic_vector(48, 8),
32865 => conv_std_logic_vector(48, 8),
32866 => conv_std_logic_vector(49, 8),
32867 => conv_std_logic_vector(49, 8),
32868 => conv_std_logic_vector(50, 8),
32869 => conv_std_logic_vector(50, 8),
32870 => conv_std_logic_vector(51, 8),
32871 => conv_std_logic_vector(51, 8),
32872 => conv_std_logic_vector(52, 8),
32873 => conv_std_logic_vector(52, 8),
32874 => conv_std_logic_vector(53, 8),
32875 => conv_std_logic_vector(53, 8),
32876 => conv_std_logic_vector(54, 8),
32877 => conv_std_logic_vector(54, 8),
32878 => conv_std_logic_vector(55, 8),
32879 => conv_std_logic_vector(55, 8),
32880 => conv_std_logic_vector(56, 8),
32881 => conv_std_logic_vector(56, 8),
32882 => conv_std_logic_vector(57, 8),
32883 => conv_std_logic_vector(57, 8),
32884 => conv_std_logic_vector(58, 8),
32885 => conv_std_logic_vector(58, 8),
32886 => conv_std_logic_vector(59, 8),
32887 => conv_std_logic_vector(59, 8),
32888 => conv_std_logic_vector(60, 8),
32889 => conv_std_logic_vector(60, 8),
32890 => conv_std_logic_vector(61, 8),
32891 => conv_std_logic_vector(61, 8),
32892 => conv_std_logic_vector(62, 8),
32893 => conv_std_logic_vector(62, 8),
32894 => conv_std_logic_vector(63, 8),
32895 => conv_std_logic_vector(63, 8),
32896 => conv_std_logic_vector(64, 8),
32897 => conv_std_logic_vector(64, 8),
32898 => conv_std_logic_vector(65, 8),
32899 => conv_std_logic_vector(65, 8),
32900 => conv_std_logic_vector(66, 8),
32901 => conv_std_logic_vector(66, 8),
32902 => conv_std_logic_vector(67, 8),
32903 => conv_std_logic_vector(67, 8),
32904 => conv_std_logic_vector(68, 8),
32905 => conv_std_logic_vector(68, 8),
32906 => conv_std_logic_vector(69, 8),
32907 => conv_std_logic_vector(69, 8),
32908 => conv_std_logic_vector(70, 8),
32909 => conv_std_logic_vector(70, 8),
32910 => conv_std_logic_vector(71, 8),
32911 => conv_std_logic_vector(71, 8),
32912 => conv_std_logic_vector(72, 8),
32913 => conv_std_logic_vector(72, 8),
32914 => conv_std_logic_vector(73, 8),
32915 => conv_std_logic_vector(73, 8),
32916 => conv_std_logic_vector(74, 8),
32917 => conv_std_logic_vector(74, 8),
32918 => conv_std_logic_vector(75, 8),
32919 => conv_std_logic_vector(75, 8),
32920 => conv_std_logic_vector(76, 8),
32921 => conv_std_logic_vector(76, 8),
32922 => conv_std_logic_vector(77, 8),
32923 => conv_std_logic_vector(77, 8),
32924 => conv_std_logic_vector(78, 8),
32925 => conv_std_logic_vector(78, 8),
32926 => conv_std_logic_vector(79, 8),
32927 => conv_std_logic_vector(79, 8),
32928 => conv_std_logic_vector(80, 8),
32929 => conv_std_logic_vector(80, 8),
32930 => conv_std_logic_vector(81, 8),
32931 => conv_std_logic_vector(81, 8),
32932 => conv_std_logic_vector(82, 8),
32933 => conv_std_logic_vector(82, 8),
32934 => conv_std_logic_vector(83, 8),
32935 => conv_std_logic_vector(83, 8),
32936 => conv_std_logic_vector(84, 8),
32937 => conv_std_logic_vector(84, 8),
32938 => conv_std_logic_vector(85, 8),
32939 => conv_std_logic_vector(85, 8),
32940 => conv_std_logic_vector(86, 8),
32941 => conv_std_logic_vector(86, 8),
32942 => conv_std_logic_vector(87, 8),
32943 => conv_std_logic_vector(87, 8),
32944 => conv_std_logic_vector(88, 8),
32945 => conv_std_logic_vector(88, 8),
32946 => conv_std_logic_vector(89, 8),
32947 => conv_std_logic_vector(89, 8),
32948 => conv_std_logic_vector(90, 8),
32949 => conv_std_logic_vector(90, 8),
32950 => conv_std_logic_vector(91, 8),
32951 => conv_std_logic_vector(91, 8),
32952 => conv_std_logic_vector(92, 8),
32953 => conv_std_logic_vector(92, 8),
32954 => conv_std_logic_vector(93, 8),
32955 => conv_std_logic_vector(93, 8),
32956 => conv_std_logic_vector(94, 8),
32957 => conv_std_logic_vector(94, 8),
32958 => conv_std_logic_vector(95, 8),
32959 => conv_std_logic_vector(95, 8),
32960 => conv_std_logic_vector(96, 8),
32961 => conv_std_logic_vector(96, 8),
32962 => conv_std_logic_vector(97, 8),
32963 => conv_std_logic_vector(97, 8),
32964 => conv_std_logic_vector(98, 8),
32965 => conv_std_logic_vector(98, 8),
32966 => conv_std_logic_vector(99, 8),
32967 => conv_std_logic_vector(99, 8),
32968 => conv_std_logic_vector(100, 8),
32969 => conv_std_logic_vector(100, 8),
32970 => conv_std_logic_vector(101, 8),
32971 => conv_std_logic_vector(101, 8),
32972 => conv_std_logic_vector(102, 8),
32973 => conv_std_logic_vector(102, 8),
32974 => conv_std_logic_vector(103, 8),
32975 => conv_std_logic_vector(103, 8),
32976 => conv_std_logic_vector(104, 8),
32977 => conv_std_logic_vector(104, 8),
32978 => conv_std_logic_vector(105, 8),
32979 => conv_std_logic_vector(105, 8),
32980 => conv_std_logic_vector(106, 8),
32981 => conv_std_logic_vector(106, 8),
32982 => conv_std_logic_vector(107, 8),
32983 => conv_std_logic_vector(107, 8),
32984 => conv_std_logic_vector(108, 8),
32985 => conv_std_logic_vector(108, 8),
32986 => conv_std_logic_vector(109, 8),
32987 => conv_std_logic_vector(109, 8),
32988 => conv_std_logic_vector(110, 8),
32989 => conv_std_logic_vector(110, 8),
32990 => conv_std_logic_vector(111, 8),
32991 => conv_std_logic_vector(111, 8),
32992 => conv_std_logic_vector(112, 8),
32993 => conv_std_logic_vector(112, 8),
32994 => conv_std_logic_vector(113, 8),
32995 => conv_std_logic_vector(113, 8),
32996 => conv_std_logic_vector(114, 8),
32997 => conv_std_logic_vector(114, 8),
32998 => conv_std_logic_vector(115, 8),
32999 => conv_std_logic_vector(115, 8),
33000 => conv_std_logic_vector(116, 8),
33001 => conv_std_logic_vector(116, 8),
33002 => conv_std_logic_vector(117, 8),
33003 => conv_std_logic_vector(117, 8),
33004 => conv_std_logic_vector(118, 8),
33005 => conv_std_logic_vector(118, 8),
33006 => conv_std_logic_vector(119, 8),
33007 => conv_std_logic_vector(119, 8),
33008 => conv_std_logic_vector(120, 8),
33009 => conv_std_logic_vector(120, 8),
33010 => conv_std_logic_vector(121, 8),
33011 => conv_std_logic_vector(121, 8),
33012 => conv_std_logic_vector(122, 8),
33013 => conv_std_logic_vector(122, 8),
33014 => conv_std_logic_vector(123, 8),
33015 => conv_std_logic_vector(123, 8),
33016 => conv_std_logic_vector(124, 8),
33017 => conv_std_logic_vector(124, 8),
33018 => conv_std_logic_vector(125, 8),
33019 => conv_std_logic_vector(125, 8),
33020 => conv_std_logic_vector(126, 8),
33021 => conv_std_logic_vector(126, 8),
33022 => conv_std_logic_vector(127, 8),
33023 => conv_std_logic_vector(127, 8),
33024 => conv_std_logic_vector(0, 8),
33025 => conv_std_logic_vector(0, 8),
33026 => conv_std_logic_vector(1, 8),
33027 => conv_std_logic_vector(1, 8),
33028 => conv_std_logic_vector(2, 8),
33029 => conv_std_logic_vector(2, 8),
33030 => conv_std_logic_vector(3, 8),
33031 => conv_std_logic_vector(3, 8),
33032 => conv_std_logic_vector(4, 8),
33033 => conv_std_logic_vector(4, 8),
33034 => conv_std_logic_vector(5, 8),
33035 => conv_std_logic_vector(5, 8),
33036 => conv_std_logic_vector(6, 8),
33037 => conv_std_logic_vector(6, 8),
33038 => conv_std_logic_vector(7, 8),
33039 => conv_std_logic_vector(7, 8),
33040 => conv_std_logic_vector(8, 8),
33041 => conv_std_logic_vector(8, 8),
33042 => conv_std_logic_vector(9, 8),
33043 => conv_std_logic_vector(9, 8),
33044 => conv_std_logic_vector(10, 8),
33045 => conv_std_logic_vector(10, 8),
33046 => conv_std_logic_vector(11, 8),
33047 => conv_std_logic_vector(11, 8),
33048 => conv_std_logic_vector(12, 8),
33049 => conv_std_logic_vector(12, 8),
33050 => conv_std_logic_vector(13, 8),
33051 => conv_std_logic_vector(13, 8),
33052 => conv_std_logic_vector(14, 8),
33053 => conv_std_logic_vector(14, 8),
33054 => conv_std_logic_vector(15, 8),
33055 => conv_std_logic_vector(15, 8),
33056 => conv_std_logic_vector(16, 8),
33057 => conv_std_logic_vector(16, 8),
33058 => conv_std_logic_vector(17, 8),
33059 => conv_std_logic_vector(17, 8),
33060 => conv_std_logic_vector(18, 8),
33061 => conv_std_logic_vector(18, 8),
33062 => conv_std_logic_vector(19, 8),
33063 => conv_std_logic_vector(19, 8),
33064 => conv_std_logic_vector(20, 8),
33065 => conv_std_logic_vector(20, 8),
33066 => conv_std_logic_vector(21, 8),
33067 => conv_std_logic_vector(21, 8),
33068 => conv_std_logic_vector(22, 8),
33069 => conv_std_logic_vector(22, 8),
33070 => conv_std_logic_vector(23, 8),
33071 => conv_std_logic_vector(23, 8),
33072 => conv_std_logic_vector(24, 8),
33073 => conv_std_logic_vector(24, 8),
33074 => conv_std_logic_vector(25, 8),
33075 => conv_std_logic_vector(25, 8),
33076 => conv_std_logic_vector(26, 8),
33077 => conv_std_logic_vector(26, 8),
33078 => conv_std_logic_vector(27, 8),
33079 => conv_std_logic_vector(27, 8),
33080 => conv_std_logic_vector(28, 8),
33081 => conv_std_logic_vector(28, 8),
33082 => conv_std_logic_vector(29, 8),
33083 => conv_std_logic_vector(29, 8),
33084 => conv_std_logic_vector(30, 8),
33085 => conv_std_logic_vector(30, 8),
33086 => conv_std_logic_vector(31, 8),
33087 => conv_std_logic_vector(31, 8),
33088 => conv_std_logic_vector(32, 8),
33089 => conv_std_logic_vector(32, 8),
33090 => conv_std_logic_vector(33, 8),
33091 => conv_std_logic_vector(33, 8),
33092 => conv_std_logic_vector(34, 8),
33093 => conv_std_logic_vector(34, 8),
33094 => conv_std_logic_vector(35, 8),
33095 => conv_std_logic_vector(35, 8),
33096 => conv_std_logic_vector(36, 8),
33097 => conv_std_logic_vector(36, 8),
33098 => conv_std_logic_vector(37, 8),
33099 => conv_std_logic_vector(37, 8),
33100 => conv_std_logic_vector(38, 8),
33101 => conv_std_logic_vector(38, 8),
33102 => conv_std_logic_vector(39, 8),
33103 => conv_std_logic_vector(39, 8),
33104 => conv_std_logic_vector(40, 8),
33105 => conv_std_logic_vector(40, 8),
33106 => conv_std_logic_vector(41, 8),
33107 => conv_std_logic_vector(41, 8),
33108 => conv_std_logic_vector(42, 8),
33109 => conv_std_logic_vector(42, 8),
33110 => conv_std_logic_vector(43, 8),
33111 => conv_std_logic_vector(43, 8),
33112 => conv_std_logic_vector(44, 8),
33113 => conv_std_logic_vector(44, 8),
33114 => conv_std_logic_vector(45, 8),
33115 => conv_std_logic_vector(45, 8),
33116 => conv_std_logic_vector(46, 8),
33117 => conv_std_logic_vector(46, 8),
33118 => conv_std_logic_vector(47, 8),
33119 => conv_std_logic_vector(47, 8),
33120 => conv_std_logic_vector(48, 8),
33121 => conv_std_logic_vector(48, 8),
33122 => conv_std_logic_vector(49, 8),
33123 => conv_std_logic_vector(49, 8),
33124 => conv_std_logic_vector(50, 8),
33125 => conv_std_logic_vector(50, 8),
33126 => conv_std_logic_vector(51, 8),
33127 => conv_std_logic_vector(51, 8),
33128 => conv_std_logic_vector(52, 8),
33129 => conv_std_logic_vector(52, 8),
33130 => conv_std_logic_vector(53, 8),
33131 => conv_std_logic_vector(53, 8),
33132 => conv_std_logic_vector(54, 8),
33133 => conv_std_logic_vector(54, 8),
33134 => conv_std_logic_vector(55, 8),
33135 => conv_std_logic_vector(55, 8),
33136 => conv_std_logic_vector(56, 8),
33137 => conv_std_logic_vector(56, 8),
33138 => conv_std_logic_vector(57, 8),
33139 => conv_std_logic_vector(57, 8),
33140 => conv_std_logic_vector(58, 8),
33141 => conv_std_logic_vector(58, 8),
33142 => conv_std_logic_vector(59, 8),
33143 => conv_std_logic_vector(59, 8),
33144 => conv_std_logic_vector(60, 8),
33145 => conv_std_logic_vector(60, 8),
33146 => conv_std_logic_vector(61, 8),
33147 => conv_std_logic_vector(61, 8),
33148 => conv_std_logic_vector(62, 8),
33149 => conv_std_logic_vector(62, 8),
33150 => conv_std_logic_vector(63, 8),
33151 => conv_std_logic_vector(63, 8),
33152 => conv_std_logic_vector(64, 8),
33153 => conv_std_logic_vector(65, 8),
33154 => conv_std_logic_vector(65, 8),
33155 => conv_std_logic_vector(66, 8),
33156 => conv_std_logic_vector(66, 8),
33157 => conv_std_logic_vector(67, 8),
33158 => conv_std_logic_vector(67, 8),
33159 => conv_std_logic_vector(68, 8),
33160 => conv_std_logic_vector(68, 8),
33161 => conv_std_logic_vector(69, 8),
33162 => conv_std_logic_vector(69, 8),
33163 => conv_std_logic_vector(70, 8),
33164 => conv_std_logic_vector(70, 8),
33165 => conv_std_logic_vector(71, 8),
33166 => conv_std_logic_vector(71, 8),
33167 => conv_std_logic_vector(72, 8),
33168 => conv_std_logic_vector(72, 8),
33169 => conv_std_logic_vector(73, 8),
33170 => conv_std_logic_vector(73, 8),
33171 => conv_std_logic_vector(74, 8),
33172 => conv_std_logic_vector(74, 8),
33173 => conv_std_logic_vector(75, 8),
33174 => conv_std_logic_vector(75, 8),
33175 => conv_std_logic_vector(76, 8),
33176 => conv_std_logic_vector(76, 8),
33177 => conv_std_logic_vector(77, 8),
33178 => conv_std_logic_vector(77, 8),
33179 => conv_std_logic_vector(78, 8),
33180 => conv_std_logic_vector(78, 8),
33181 => conv_std_logic_vector(79, 8),
33182 => conv_std_logic_vector(79, 8),
33183 => conv_std_logic_vector(80, 8),
33184 => conv_std_logic_vector(80, 8),
33185 => conv_std_logic_vector(81, 8),
33186 => conv_std_logic_vector(81, 8),
33187 => conv_std_logic_vector(82, 8),
33188 => conv_std_logic_vector(82, 8),
33189 => conv_std_logic_vector(83, 8),
33190 => conv_std_logic_vector(83, 8),
33191 => conv_std_logic_vector(84, 8),
33192 => conv_std_logic_vector(84, 8),
33193 => conv_std_logic_vector(85, 8),
33194 => conv_std_logic_vector(85, 8),
33195 => conv_std_logic_vector(86, 8),
33196 => conv_std_logic_vector(86, 8),
33197 => conv_std_logic_vector(87, 8),
33198 => conv_std_logic_vector(87, 8),
33199 => conv_std_logic_vector(88, 8),
33200 => conv_std_logic_vector(88, 8),
33201 => conv_std_logic_vector(89, 8),
33202 => conv_std_logic_vector(89, 8),
33203 => conv_std_logic_vector(90, 8),
33204 => conv_std_logic_vector(90, 8),
33205 => conv_std_logic_vector(91, 8),
33206 => conv_std_logic_vector(91, 8),
33207 => conv_std_logic_vector(92, 8),
33208 => conv_std_logic_vector(92, 8),
33209 => conv_std_logic_vector(93, 8),
33210 => conv_std_logic_vector(93, 8),
33211 => conv_std_logic_vector(94, 8),
33212 => conv_std_logic_vector(94, 8),
33213 => conv_std_logic_vector(95, 8),
33214 => conv_std_logic_vector(95, 8),
33215 => conv_std_logic_vector(96, 8),
33216 => conv_std_logic_vector(96, 8),
33217 => conv_std_logic_vector(97, 8),
33218 => conv_std_logic_vector(97, 8),
33219 => conv_std_logic_vector(98, 8),
33220 => conv_std_logic_vector(98, 8),
33221 => conv_std_logic_vector(99, 8),
33222 => conv_std_logic_vector(99, 8),
33223 => conv_std_logic_vector(100, 8),
33224 => conv_std_logic_vector(100, 8),
33225 => conv_std_logic_vector(101, 8),
33226 => conv_std_logic_vector(101, 8),
33227 => conv_std_logic_vector(102, 8),
33228 => conv_std_logic_vector(102, 8),
33229 => conv_std_logic_vector(103, 8),
33230 => conv_std_logic_vector(103, 8),
33231 => conv_std_logic_vector(104, 8),
33232 => conv_std_logic_vector(104, 8),
33233 => conv_std_logic_vector(105, 8),
33234 => conv_std_logic_vector(105, 8),
33235 => conv_std_logic_vector(106, 8),
33236 => conv_std_logic_vector(106, 8),
33237 => conv_std_logic_vector(107, 8),
33238 => conv_std_logic_vector(107, 8),
33239 => conv_std_logic_vector(108, 8),
33240 => conv_std_logic_vector(108, 8),
33241 => conv_std_logic_vector(109, 8),
33242 => conv_std_logic_vector(109, 8),
33243 => conv_std_logic_vector(110, 8),
33244 => conv_std_logic_vector(110, 8),
33245 => conv_std_logic_vector(111, 8),
33246 => conv_std_logic_vector(111, 8),
33247 => conv_std_logic_vector(112, 8),
33248 => conv_std_logic_vector(112, 8),
33249 => conv_std_logic_vector(113, 8),
33250 => conv_std_logic_vector(113, 8),
33251 => conv_std_logic_vector(114, 8),
33252 => conv_std_logic_vector(114, 8),
33253 => conv_std_logic_vector(115, 8),
33254 => conv_std_logic_vector(115, 8),
33255 => conv_std_logic_vector(116, 8),
33256 => conv_std_logic_vector(116, 8),
33257 => conv_std_logic_vector(117, 8),
33258 => conv_std_logic_vector(117, 8),
33259 => conv_std_logic_vector(118, 8),
33260 => conv_std_logic_vector(118, 8),
33261 => conv_std_logic_vector(119, 8),
33262 => conv_std_logic_vector(119, 8),
33263 => conv_std_logic_vector(120, 8),
33264 => conv_std_logic_vector(120, 8),
33265 => conv_std_logic_vector(121, 8),
33266 => conv_std_logic_vector(121, 8),
33267 => conv_std_logic_vector(122, 8),
33268 => conv_std_logic_vector(122, 8),
33269 => conv_std_logic_vector(123, 8),
33270 => conv_std_logic_vector(123, 8),
33271 => conv_std_logic_vector(124, 8),
33272 => conv_std_logic_vector(124, 8),
33273 => conv_std_logic_vector(125, 8),
33274 => conv_std_logic_vector(125, 8),
33275 => conv_std_logic_vector(126, 8),
33276 => conv_std_logic_vector(126, 8),
33277 => conv_std_logic_vector(127, 8),
33278 => conv_std_logic_vector(127, 8),
33279 => conv_std_logic_vector(128, 8),
33280 => conv_std_logic_vector(0, 8),
33281 => conv_std_logic_vector(0, 8),
33282 => conv_std_logic_vector(1, 8),
33283 => conv_std_logic_vector(1, 8),
33284 => conv_std_logic_vector(2, 8),
33285 => conv_std_logic_vector(2, 8),
33286 => conv_std_logic_vector(3, 8),
33287 => conv_std_logic_vector(3, 8),
33288 => conv_std_logic_vector(4, 8),
33289 => conv_std_logic_vector(4, 8),
33290 => conv_std_logic_vector(5, 8),
33291 => conv_std_logic_vector(5, 8),
33292 => conv_std_logic_vector(6, 8),
33293 => conv_std_logic_vector(6, 8),
33294 => conv_std_logic_vector(7, 8),
33295 => conv_std_logic_vector(7, 8),
33296 => conv_std_logic_vector(8, 8),
33297 => conv_std_logic_vector(8, 8),
33298 => conv_std_logic_vector(9, 8),
33299 => conv_std_logic_vector(9, 8),
33300 => conv_std_logic_vector(10, 8),
33301 => conv_std_logic_vector(10, 8),
33302 => conv_std_logic_vector(11, 8),
33303 => conv_std_logic_vector(11, 8),
33304 => conv_std_logic_vector(12, 8),
33305 => conv_std_logic_vector(12, 8),
33306 => conv_std_logic_vector(13, 8),
33307 => conv_std_logic_vector(13, 8),
33308 => conv_std_logic_vector(14, 8),
33309 => conv_std_logic_vector(14, 8),
33310 => conv_std_logic_vector(15, 8),
33311 => conv_std_logic_vector(15, 8),
33312 => conv_std_logic_vector(16, 8),
33313 => conv_std_logic_vector(16, 8),
33314 => conv_std_logic_vector(17, 8),
33315 => conv_std_logic_vector(17, 8),
33316 => conv_std_logic_vector(18, 8),
33317 => conv_std_logic_vector(18, 8),
33318 => conv_std_logic_vector(19, 8),
33319 => conv_std_logic_vector(19, 8),
33320 => conv_std_logic_vector(20, 8),
33321 => conv_std_logic_vector(20, 8),
33322 => conv_std_logic_vector(21, 8),
33323 => conv_std_logic_vector(21, 8),
33324 => conv_std_logic_vector(22, 8),
33325 => conv_std_logic_vector(22, 8),
33326 => conv_std_logic_vector(23, 8),
33327 => conv_std_logic_vector(23, 8),
33328 => conv_std_logic_vector(24, 8),
33329 => conv_std_logic_vector(24, 8),
33330 => conv_std_logic_vector(25, 8),
33331 => conv_std_logic_vector(25, 8),
33332 => conv_std_logic_vector(26, 8),
33333 => conv_std_logic_vector(26, 8),
33334 => conv_std_logic_vector(27, 8),
33335 => conv_std_logic_vector(27, 8),
33336 => conv_std_logic_vector(28, 8),
33337 => conv_std_logic_vector(28, 8),
33338 => conv_std_logic_vector(29, 8),
33339 => conv_std_logic_vector(29, 8),
33340 => conv_std_logic_vector(30, 8),
33341 => conv_std_logic_vector(30, 8),
33342 => conv_std_logic_vector(31, 8),
33343 => conv_std_logic_vector(31, 8),
33344 => conv_std_logic_vector(32, 8),
33345 => conv_std_logic_vector(33, 8),
33346 => conv_std_logic_vector(33, 8),
33347 => conv_std_logic_vector(34, 8),
33348 => conv_std_logic_vector(34, 8),
33349 => conv_std_logic_vector(35, 8),
33350 => conv_std_logic_vector(35, 8),
33351 => conv_std_logic_vector(36, 8),
33352 => conv_std_logic_vector(36, 8),
33353 => conv_std_logic_vector(37, 8),
33354 => conv_std_logic_vector(37, 8),
33355 => conv_std_logic_vector(38, 8),
33356 => conv_std_logic_vector(38, 8),
33357 => conv_std_logic_vector(39, 8),
33358 => conv_std_logic_vector(39, 8),
33359 => conv_std_logic_vector(40, 8),
33360 => conv_std_logic_vector(40, 8),
33361 => conv_std_logic_vector(41, 8),
33362 => conv_std_logic_vector(41, 8),
33363 => conv_std_logic_vector(42, 8),
33364 => conv_std_logic_vector(42, 8),
33365 => conv_std_logic_vector(43, 8),
33366 => conv_std_logic_vector(43, 8),
33367 => conv_std_logic_vector(44, 8),
33368 => conv_std_logic_vector(44, 8),
33369 => conv_std_logic_vector(45, 8),
33370 => conv_std_logic_vector(45, 8),
33371 => conv_std_logic_vector(46, 8),
33372 => conv_std_logic_vector(46, 8),
33373 => conv_std_logic_vector(47, 8),
33374 => conv_std_logic_vector(47, 8),
33375 => conv_std_logic_vector(48, 8),
33376 => conv_std_logic_vector(48, 8),
33377 => conv_std_logic_vector(49, 8),
33378 => conv_std_logic_vector(49, 8),
33379 => conv_std_logic_vector(50, 8),
33380 => conv_std_logic_vector(50, 8),
33381 => conv_std_logic_vector(51, 8),
33382 => conv_std_logic_vector(51, 8),
33383 => conv_std_logic_vector(52, 8),
33384 => conv_std_logic_vector(52, 8),
33385 => conv_std_logic_vector(53, 8),
33386 => conv_std_logic_vector(53, 8),
33387 => conv_std_logic_vector(54, 8),
33388 => conv_std_logic_vector(54, 8),
33389 => conv_std_logic_vector(55, 8),
33390 => conv_std_logic_vector(55, 8),
33391 => conv_std_logic_vector(56, 8),
33392 => conv_std_logic_vector(56, 8),
33393 => conv_std_logic_vector(57, 8),
33394 => conv_std_logic_vector(57, 8),
33395 => conv_std_logic_vector(58, 8),
33396 => conv_std_logic_vector(58, 8),
33397 => conv_std_logic_vector(59, 8),
33398 => conv_std_logic_vector(59, 8),
33399 => conv_std_logic_vector(60, 8),
33400 => conv_std_logic_vector(60, 8),
33401 => conv_std_logic_vector(61, 8),
33402 => conv_std_logic_vector(61, 8),
33403 => conv_std_logic_vector(62, 8),
33404 => conv_std_logic_vector(62, 8),
33405 => conv_std_logic_vector(63, 8),
33406 => conv_std_logic_vector(63, 8),
33407 => conv_std_logic_vector(64, 8),
33408 => conv_std_logic_vector(65, 8),
33409 => conv_std_logic_vector(65, 8),
33410 => conv_std_logic_vector(66, 8),
33411 => conv_std_logic_vector(66, 8),
33412 => conv_std_logic_vector(67, 8),
33413 => conv_std_logic_vector(67, 8),
33414 => conv_std_logic_vector(68, 8),
33415 => conv_std_logic_vector(68, 8),
33416 => conv_std_logic_vector(69, 8),
33417 => conv_std_logic_vector(69, 8),
33418 => conv_std_logic_vector(70, 8),
33419 => conv_std_logic_vector(70, 8),
33420 => conv_std_logic_vector(71, 8),
33421 => conv_std_logic_vector(71, 8),
33422 => conv_std_logic_vector(72, 8),
33423 => conv_std_logic_vector(72, 8),
33424 => conv_std_logic_vector(73, 8),
33425 => conv_std_logic_vector(73, 8),
33426 => conv_std_logic_vector(74, 8),
33427 => conv_std_logic_vector(74, 8),
33428 => conv_std_logic_vector(75, 8),
33429 => conv_std_logic_vector(75, 8),
33430 => conv_std_logic_vector(76, 8),
33431 => conv_std_logic_vector(76, 8),
33432 => conv_std_logic_vector(77, 8),
33433 => conv_std_logic_vector(77, 8),
33434 => conv_std_logic_vector(78, 8),
33435 => conv_std_logic_vector(78, 8),
33436 => conv_std_logic_vector(79, 8),
33437 => conv_std_logic_vector(79, 8),
33438 => conv_std_logic_vector(80, 8),
33439 => conv_std_logic_vector(80, 8),
33440 => conv_std_logic_vector(81, 8),
33441 => conv_std_logic_vector(81, 8),
33442 => conv_std_logic_vector(82, 8),
33443 => conv_std_logic_vector(82, 8),
33444 => conv_std_logic_vector(83, 8),
33445 => conv_std_logic_vector(83, 8),
33446 => conv_std_logic_vector(84, 8),
33447 => conv_std_logic_vector(84, 8),
33448 => conv_std_logic_vector(85, 8),
33449 => conv_std_logic_vector(85, 8),
33450 => conv_std_logic_vector(86, 8),
33451 => conv_std_logic_vector(86, 8),
33452 => conv_std_logic_vector(87, 8),
33453 => conv_std_logic_vector(87, 8),
33454 => conv_std_logic_vector(88, 8),
33455 => conv_std_logic_vector(88, 8),
33456 => conv_std_logic_vector(89, 8),
33457 => conv_std_logic_vector(89, 8),
33458 => conv_std_logic_vector(90, 8),
33459 => conv_std_logic_vector(90, 8),
33460 => conv_std_logic_vector(91, 8),
33461 => conv_std_logic_vector(91, 8),
33462 => conv_std_logic_vector(92, 8),
33463 => conv_std_logic_vector(92, 8),
33464 => conv_std_logic_vector(93, 8),
33465 => conv_std_logic_vector(93, 8),
33466 => conv_std_logic_vector(94, 8),
33467 => conv_std_logic_vector(94, 8),
33468 => conv_std_logic_vector(95, 8),
33469 => conv_std_logic_vector(95, 8),
33470 => conv_std_logic_vector(96, 8),
33471 => conv_std_logic_vector(96, 8),
33472 => conv_std_logic_vector(97, 8),
33473 => conv_std_logic_vector(98, 8),
33474 => conv_std_logic_vector(98, 8),
33475 => conv_std_logic_vector(99, 8),
33476 => conv_std_logic_vector(99, 8),
33477 => conv_std_logic_vector(100, 8),
33478 => conv_std_logic_vector(100, 8),
33479 => conv_std_logic_vector(101, 8),
33480 => conv_std_logic_vector(101, 8),
33481 => conv_std_logic_vector(102, 8),
33482 => conv_std_logic_vector(102, 8),
33483 => conv_std_logic_vector(103, 8),
33484 => conv_std_logic_vector(103, 8),
33485 => conv_std_logic_vector(104, 8),
33486 => conv_std_logic_vector(104, 8),
33487 => conv_std_logic_vector(105, 8),
33488 => conv_std_logic_vector(105, 8),
33489 => conv_std_logic_vector(106, 8),
33490 => conv_std_logic_vector(106, 8),
33491 => conv_std_logic_vector(107, 8),
33492 => conv_std_logic_vector(107, 8),
33493 => conv_std_logic_vector(108, 8),
33494 => conv_std_logic_vector(108, 8),
33495 => conv_std_logic_vector(109, 8),
33496 => conv_std_logic_vector(109, 8),
33497 => conv_std_logic_vector(110, 8),
33498 => conv_std_logic_vector(110, 8),
33499 => conv_std_logic_vector(111, 8),
33500 => conv_std_logic_vector(111, 8),
33501 => conv_std_logic_vector(112, 8),
33502 => conv_std_logic_vector(112, 8),
33503 => conv_std_logic_vector(113, 8),
33504 => conv_std_logic_vector(113, 8),
33505 => conv_std_logic_vector(114, 8),
33506 => conv_std_logic_vector(114, 8),
33507 => conv_std_logic_vector(115, 8),
33508 => conv_std_logic_vector(115, 8),
33509 => conv_std_logic_vector(116, 8),
33510 => conv_std_logic_vector(116, 8),
33511 => conv_std_logic_vector(117, 8),
33512 => conv_std_logic_vector(117, 8),
33513 => conv_std_logic_vector(118, 8),
33514 => conv_std_logic_vector(118, 8),
33515 => conv_std_logic_vector(119, 8),
33516 => conv_std_logic_vector(119, 8),
33517 => conv_std_logic_vector(120, 8),
33518 => conv_std_logic_vector(120, 8),
33519 => conv_std_logic_vector(121, 8),
33520 => conv_std_logic_vector(121, 8),
33521 => conv_std_logic_vector(122, 8),
33522 => conv_std_logic_vector(122, 8),
33523 => conv_std_logic_vector(123, 8),
33524 => conv_std_logic_vector(123, 8),
33525 => conv_std_logic_vector(124, 8),
33526 => conv_std_logic_vector(124, 8),
33527 => conv_std_logic_vector(125, 8),
33528 => conv_std_logic_vector(125, 8),
33529 => conv_std_logic_vector(126, 8),
33530 => conv_std_logic_vector(126, 8),
33531 => conv_std_logic_vector(127, 8),
33532 => conv_std_logic_vector(127, 8),
33533 => conv_std_logic_vector(128, 8),
33534 => conv_std_logic_vector(128, 8),
33535 => conv_std_logic_vector(129, 8),
33536 => conv_std_logic_vector(0, 8),
33537 => conv_std_logic_vector(0, 8),
33538 => conv_std_logic_vector(1, 8),
33539 => conv_std_logic_vector(1, 8),
33540 => conv_std_logic_vector(2, 8),
33541 => conv_std_logic_vector(2, 8),
33542 => conv_std_logic_vector(3, 8),
33543 => conv_std_logic_vector(3, 8),
33544 => conv_std_logic_vector(4, 8),
33545 => conv_std_logic_vector(4, 8),
33546 => conv_std_logic_vector(5, 8),
33547 => conv_std_logic_vector(5, 8),
33548 => conv_std_logic_vector(6, 8),
33549 => conv_std_logic_vector(6, 8),
33550 => conv_std_logic_vector(7, 8),
33551 => conv_std_logic_vector(7, 8),
33552 => conv_std_logic_vector(8, 8),
33553 => conv_std_logic_vector(8, 8),
33554 => conv_std_logic_vector(9, 8),
33555 => conv_std_logic_vector(9, 8),
33556 => conv_std_logic_vector(10, 8),
33557 => conv_std_logic_vector(10, 8),
33558 => conv_std_logic_vector(11, 8),
33559 => conv_std_logic_vector(11, 8),
33560 => conv_std_logic_vector(12, 8),
33561 => conv_std_logic_vector(12, 8),
33562 => conv_std_logic_vector(13, 8),
33563 => conv_std_logic_vector(13, 8),
33564 => conv_std_logic_vector(14, 8),
33565 => conv_std_logic_vector(14, 8),
33566 => conv_std_logic_vector(15, 8),
33567 => conv_std_logic_vector(15, 8),
33568 => conv_std_logic_vector(16, 8),
33569 => conv_std_logic_vector(16, 8),
33570 => conv_std_logic_vector(17, 8),
33571 => conv_std_logic_vector(17, 8),
33572 => conv_std_logic_vector(18, 8),
33573 => conv_std_logic_vector(18, 8),
33574 => conv_std_logic_vector(19, 8),
33575 => conv_std_logic_vector(19, 8),
33576 => conv_std_logic_vector(20, 8),
33577 => conv_std_logic_vector(20, 8),
33578 => conv_std_logic_vector(21, 8),
33579 => conv_std_logic_vector(22, 8),
33580 => conv_std_logic_vector(22, 8),
33581 => conv_std_logic_vector(23, 8),
33582 => conv_std_logic_vector(23, 8),
33583 => conv_std_logic_vector(24, 8),
33584 => conv_std_logic_vector(24, 8),
33585 => conv_std_logic_vector(25, 8),
33586 => conv_std_logic_vector(25, 8),
33587 => conv_std_logic_vector(26, 8),
33588 => conv_std_logic_vector(26, 8),
33589 => conv_std_logic_vector(27, 8),
33590 => conv_std_logic_vector(27, 8),
33591 => conv_std_logic_vector(28, 8),
33592 => conv_std_logic_vector(28, 8),
33593 => conv_std_logic_vector(29, 8),
33594 => conv_std_logic_vector(29, 8),
33595 => conv_std_logic_vector(30, 8),
33596 => conv_std_logic_vector(30, 8),
33597 => conv_std_logic_vector(31, 8),
33598 => conv_std_logic_vector(31, 8),
33599 => conv_std_logic_vector(32, 8),
33600 => conv_std_logic_vector(32, 8),
33601 => conv_std_logic_vector(33, 8),
33602 => conv_std_logic_vector(33, 8),
33603 => conv_std_logic_vector(34, 8),
33604 => conv_std_logic_vector(34, 8),
33605 => conv_std_logic_vector(35, 8),
33606 => conv_std_logic_vector(35, 8),
33607 => conv_std_logic_vector(36, 8),
33608 => conv_std_logic_vector(36, 8),
33609 => conv_std_logic_vector(37, 8),
33610 => conv_std_logic_vector(37, 8),
33611 => conv_std_logic_vector(38, 8),
33612 => conv_std_logic_vector(38, 8),
33613 => conv_std_logic_vector(39, 8),
33614 => conv_std_logic_vector(39, 8),
33615 => conv_std_logic_vector(40, 8),
33616 => conv_std_logic_vector(40, 8),
33617 => conv_std_logic_vector(41, 8),
33618 => conv_std_logic_vector(41, 8),
33619 => conv_std_logic_vector(42, 8),
33620 => conv_std_logic_vector(42, 8),
33621 => conv_std_logic_vector(43, 8),
33622 => conv_std_logic_vector(44, 8),
33623 => conv_std_logic_vector(44, 8),
33624 => conv_std_logic_vector(45, 8),
33625 => conv_std_logic_vector(45, 8),
33626 => conv_std_logic_vector(46, 8),
33627 => conv_std_logic_vector(46, 8),
33628 => conv_std_logic_vector(47, 8),
33629 => conv_std_logic_vector(47, 8),
33630 => conv_std_logic_vector(48, 8),
33631 => conv_std_logic_vector(48, 8),
33632 => conv_std_logic_vector(49, 8),
33633 => conv_std_logic_vector(49, 8),
33634 => conv_std_logic_vector(50, 8),
33635 => conv_std_logic_vector(50, 8),
33636 => conv_std_logic_vector(51, 8),
33637 => conv_std_logic_vector(51, 8),
33638 => conv_std_logic_vector(52, 8),
33639 => conv_std_logic_vector(52, 8),
33640 => conv_std_logic_vector(53, 8),
33641 => conv_std_logic_vector(53, 8),
33642 => conv_std_logic_vector(54, 8),
33643 => conv_std_logic_vector(54, 8),
33644 => conv_std_logic_vector(55, 8),
33645 => conv_std_logic_vector(55, 8),
33646 => conv_std_logic_vector(56, 8),
33647 => conv_std_logic_vector(56, 8),
33648 => conv_std_logic_vector(57, 8),
33649 => conv_std_logic_vector(57, 8),
33650 => conv_std_logic_vector(58, 8),
33651 => conv_std_logic_vector(58, 8),
33652 => conv_std_logic_vector(59, 8),
33653 => conv_std_logic_vector(59, 8),
33654 => conv_std_logic_vector(60, 8),
33655 => conv_std_logic_vector(60, 8),
33656 => conv_std_logic_vector(61, 8),
33657 => conv_std_logic_vector(61, 8),
33658 => conv_std_logic_vector(62, 8),
33659 => conv_std_logic_vector(62, 8),
33660 => conv_std_logic_vector(63, 8),
33661 => conv_std_logic_vector(63, 8),
33662 => conv_std_logic_vector(64, 8),
33663 => conv_std_logic_vector(64, 8),
33664 => conv_std_logic_vector(65, 8),
33665 => conv_std_logic_vector(66, 8),
33666 => conv_std_logic_vector(66, 8),
33667 => conv_std_logic_vector(67, 8),
33668 => conv_std_logic_vector(67, 8),
33669 => conv_std_logic_vector(68, 8),
33670 => conv_std_logic_vector(68, 8),
33671 => conv_std_logic_vector(69, 8),
33672 => conv_std_logic_vector(69, 8),
33673 => conv_std_logic_vector(70, 8),
33674 => conv_std_logic_vector(70, 8),
33675 => conv_std_logic_vector(71, 8),
33676 => conv_std_logic_vector(71, 8),
33677 => conv_std_logic_vector(72, 8),
33678 => conv_std_logic_vector(72, 8),
33679 => conv_std_logic_vector(73, 8),
33680 => conv_std_logic_vector(73, 8),
33681 => conv_std_logic_vector(74, 8),
33682 => conv_std_logic_vector(74, 8),
33683 => conv_std_logic_vector(75, 8),
33684 => conv_std_logic_vector(75, 8),
33685 => conv_std_logic_vector(76, 8),
33686 => conv_std_logic_vector(76, 8),
33687 => conv_std_logic_vector(77, 8),
33688 => conv_std_logic_vector(77, 8),
33689 => conv_std_logic_vector(78, 8),
33690 => conv_std_logic_vector(78, 8),
33691 => conv_std_logic_vector(79, 8),
33692 => conv_std_logic_vector(79, 8),
33693 => conv_std_logic_vector(80, 8),
33694 => conv_std_logic_vector(80, 8),
33695 => conv_std_logic_vector(81, 8),
33696 => conv_std_logic_vector(81, 8),
33697 => conv_std_logic_vector(82, 8),
33698 => conv_std_logic_vector(82, 8),
33699 => conv_std_logic_vector(83, 8),
33700 => conv_std_logic_vector(83, 8),
33701 => conv_std_logic_vector(84, 8),
33702 => conv_std_logic_vector(84, 8),
33703 => conv_std_logic_vector(85, 8),
33704 => conv_std_logic_vector(85, 8),
33705 => conv_std_logic_vector(86, 8),
33706 => conv_std_logic_vector(86, 8),
33707 => conv_std_logic_vector(87, 8),
33708 => conv_std_logic_vector(88, 8),
33709 => conv_std_logic_vector(88, 8),
33710 => conv_std_logic_vector(89, 8),
33711 => conv_std_logic_vector(89, 8),
33712 => conv_std_logic_vector(90, 8),
33713 => conv_std_logic_vector(90, 8),
33714 => conv_std_logic_vector(91, 8),
33715 => conv_std_logic_vector(91, 8),
33716 => conv_std_logic_vector(92, 8),
33717 => conv_std_logic_vector(92, 8),
33718 => conv_std_logic_vector(93, 8),
33719 => conv_std_logic_vector(93, 8),
33720 => conv_std_logic_vector(94, 8),
33721 => conv_std_logic_vector(94, 8),
33722 => conv_std_logic_vector(95, 8),
33723 => conv_std_logic_vector(95, 8),
33724 => conv_std_logic_vector(96, 8),
33725 => conv_std_logic_vector(96, 8),
33726 => conv_std_logic_vector(97, 8),
33727 => conv_std_logic_vector(97, 8),
33728 => conv_std_logic_vector(98, 8),
33729 => conv_std_logic_vector(98, 8),
33730 => conv_std_logic_vector(99, 8),
33731 => conv_std_logic_vector(99, 8),
33732 => conv_std_logic_vector(100, 8),
33733 => conv_std_logic_vector(100, 8),
33734 => conv_std_logic_vector(101, 8),
33735 => conv_std_logic_vector(101, 8),
33736 => conv_std_logic_vector(102, 8),
33737 => conv_std_logic_vector(102, 8),
33738 => conv_std_logic_vector(103, 8),
33739 => conv_std_logic_vector(103, 8),
33740 => conv_std_logic_vector(104, 8),
33741 => conv_std_logic_vector(104, 8),
33742 => conv_std_logic_vector(105, 8),
33743 => conv_std_logic_vector(105, 8),
33744 => conv_std_logic_vector(106, 8),
33745 => conv_std_logic_vector(106, 8),
33746 => conv_std_logic_vector(107, 8),
33747 => conv_std_logic_vector(107, 8),
33748 => conv_std_logic_vector(108, 8),
33749 => conv_std_logic_vector(108, 8),
33750 => conv_std_logic_vector(109, 8),
33751 => conv_std_logic_vector(110, 8),
33752 => conv_std_logic_vector(110, 8),
33753 => conv_std_logic_vector(111, 8),
33754 => conv_std_logic_vector(111, 8),
33755 => conv_std_logic_vector(112, 8),
33756 => conv_std_logic_vector(112, 8),
33757 => conv_std_logic_vector(113, 8),
33758 => conv_std_logic_vector(113, 8),
33759 => conv_std_logic_vector(114, 8),
33760 => conv_std_logic_vector(114, 8),
33761 => conv_std_logic_vector(115, 8),
33762 => conv_std_logic_vector(115, 8),
33763 => conv_std_logic_vector(116, 8),
33764 => conv_std_logic_vector(116, 8),
33765 => conv_std_logic_vector(117, 8),
33766 => conv_std_logic_vector(117, 8),
33767 => conv_std_logic_vector(118, 8),
33768 => conv_std_logic_vector(118, 8),
33769 => conv_std_logic_vector(119, 8),
33770 => conv_std_logic_vector(119, 8),
33771 => conv_std_logic_vector(120, 8),
33772 => conv_std_logic_vector(120, 8),
33773 => conv_std_logic_vector(121, 8),
33774 => conv_std_logic_vector(121, 8),
33775 => conv_std_logic_vector(122, 8),
33776 => conv_std_logic_vector(122, 8),
33777 => conv_std_logic_vector(123, 8),
33778 => conv_std_logic_vector(123, 8),
33779 => conv_std_logic_vector(124, 8),
33780 => conv_std_logic_vector(124, 8),
33781 => conv_std_logic_vector(125, 8),
33782 => conv_std_logic_vector(125, 8),
33783 => conv_std_logic_vector(126, 8),
33784 => conv_std_logic_vector(126, 8),
33785 => conv_std_logic_vector(127, 8),
33786 => conv_std_logic_vector(127, 8),
33787 => conv_std_logic_vector(128, 8),
33788 => conv_std_logic_vector(128, 8),
33789 => conv_std_logic_vector(129, 8),
33790 => conv_std_logic_vector(129, 8),
33791 => conv_std_logic_vector(130, 8),
33792 => conv_std_logic_vector(0, 8),
33793 => conv_std_logic_vector(0, 8),
33794 => conv_std_logic_vector(1, 8),
33795 => conv_std_logic_vector(1, 8),
33796 => conv_std_logic_vector(2, 8),
33797 => conv_std_logic_vector(2, 8),
33798 => conv_std_logic_vector(3, 8),
33799 => conv_std_logic_vector(3, 8),
33800 => conv_std_logic_vector(4, 8),
33801 => conv_std_logic_vector(4, 8),
33802 => conv_std_logic_vector(5, 8),
33803 => conv_std_logic_vector(5, 8),
33804 => conv_std_logic_vector(6, 8),
33805 => conv_std_logic_vector(6, 8),
33806 => conv_std_logic_vector(7, 8),
33807 => conv_std_logic_vector(7, 8),
33808 => conv_std_logic_vector(8, 8),
33809 => conv_std_logic_vector(8, 8),
33810 => conv_std_logic_vector(9, 8),
33811 => conv_std_logic_vector(9, 8),
33812 => conv_std_logic_vector(10, 8),
33813 => conv_std_logic_vector(10, 8),
33814 => conv_std_logic_vector(11, 8),
33815 => conv_std_logic_vector(11, 8),
33816 => conv_std_logic_vector(12, 8),
33817 => conv_std_logic_vector(12, 8),
33818 => conv_std_logic_vector(13, 8),
33819 => conv_std_logic_vector(13, 8),
33820 => conv_std_logic_vector(14, 8),
33821 => conv_std_logic_vector(14, 8),
33822 => conv_std_logic_vector(15, 8),
33823 => conv_std_logic_vector(15, 8),
33824 => conv_std_logic_vector(16, 8),
33825 => conv_std_logic_vector(17, 8),
33826 => conv_std_logic_vector(17, 8),
33827 => conv_std_logic_vector(18, 8),
33828 => conv_std_logic_vector(18, 8),
33829 => conv_std_logic_vector(19, 8),
33830 => conv_std_logic_vector(19, 8),
33831 => conv_std_logic_vector(20, 8),
33832 => conv_std_logic_vector(20, 8),
33833 => conv_std_logic_vector(21, 8),
33834 => conv_std_logic_vector(21, 8),
33835 => conv_std_logic_vector(22, 8),
33836 => conv_std_logic_vector(22, 8),
33837 => conv_std_logic_vector(23, 8),
33838 => conv_std_logic_vector(23, 8),
33839 => conv_std_logic_vector(24, 8),
33840 => conv_std_logic_vector(24, 8),
33841 => conv_std_logic_vector(25, 8),
33842 => conv_std_logic_vector(25, 8),
33843 => conv_std_logic_vector(26, 8),
33844 => conv_std_logic_vector(26, 8),
33845 => conv_std_logic_vector(27, 8),
33846 => conv_std_logic_vector(27, 8),
33847 => conv_std_logic_vector(28, 8),
33848 => conv_std_logic_vector(28, 8),
33849 => conv_std_logic_vector(29, 8),
33850 => conv_std_logic_vector(29, 8),
33851 => conv_std_logic_vector(30, 8),
33852 => conv_std_logic_vector(30, 8),
33853 => conv_std_logic_vector(31, 8),
33854 => conv_std_logic_vector(31, 8),
33855 => conv_std_logic_vector(32, 8),
33856 => conv_std_logic_vector(33, 8),
33857 => conv_std_logic_vector(33, 8),
33858 => conv_std_logic_vector(34, 8),
33859 => conv_std_logic_vector(34, 8),
33860 => conv_std_logic_vector(35, 8),
33861 => conv_std_logic_vector(35, 8),
33862 => conv_std_logic_vector(36, 8),
33863 => conv_std_logic_vector(36, 8),
33864 => conv_std_logic_vector(37, 8),
33865 => conv_std_logic_vector(37, 8),
33866 => conv_std_logic_vector(38, 8),
33867 => conv_std_logic_vector(38, 8),
33868 => conv_std_logic_vector(39, 8),
33869 => conv_std_logic_vector(39, 8),
33870 => conv_std_logic_vector(40, 8),
33871 => conv_std_logic_vector(40, 8),
33872 => conv_std_logic_vector(41, 8),
33873 => conv_std_logic_vector(41, 8),
33874 => conv_std_logic_vector(42, 8),
33875 => conv_std_logic_vector(42, 8),
33876 => conv_std_logic_vector(43, 8),
33877 => conv_std_logic_vector(43, 8),
33878 => conv_std_logic_vector(44, 8),
33879 => conv_std_logic_vector(44, 8),
33880 => conv_std_logic_vector(45, 8),
33881 => conv_std_logic_vector(45, 8),
33882 => conv_std_logic_vector(46, 8),
33883 => conv_std_logic_vector(46, 8),
33884 => conv_std_logic_vector(47, 8),
33885 => conv_std_logic_vector(47, 8),
33886 => conv_std_logic_vector(48, 8),
33887 => conv_std_logic_vector(48, 8),
33888 => conv_std_logic_vector(49, 8),
33889 => conv_std_logic_vector(50, 8),
33890 => conv_std_logic_vector(50, 8),
33891 => conv_std_logic_vector(51, 8),
33892 => conv_std_logic_vector(51, 8),
33893 => conv_std_logic_vector(52, 8),
33894 => conv_std_logic_vector(52, 8),
33895 => conv_std_logic_vector(53, 8),
33896 => conv_std_logic_vector(53, 8),
33897 => conv_std_logic_vector(54, 8),
33898 => conv_std_logic_vector(54, 8),
33899 => conv_std_logic_vector(55, 8),
33900 => conv_std_logic_vector(55, 8),
33901 => conv_std_logic_vector(56, 8),
33902 => conv_std_logic_vector(56, 8),
33903 => conv_std_logic_vector(57, 8),
33904 => conv_std_logic_vector(57, 8),
33905 => conv_std_logic_vector(58, 8),
33906 => conv_std_logic_vector(58, 8),
33907 => conv_std_logic_vector(59, 8),
33908 => conv_std_logic_vector(59, 8),
33909 => conv_std_logic_vector(60, 8),
33910 => conv_std_logic_vector(60, 8),
33911 => conv_std_logic_vector(61, 8),
33912 => conv_std_logic_vector(61, 8),
33913 => conv_std_logic_vector(62, 8),
33914 => conv_std_logic_vector(62, 8),
33915 => conv_std_logic_vector(63, 8),
33916 => conv_std_logic_vector(63, 8),
33917 => conv_std_logic_vector(64, 8),
33918 => conv_std_logic_vector(64, 8),
33919 => conv_std_logic_vector(65, 8),
33920 => conv_std_logic_vector(66, 8),
33921 => conv_std_logic_vector(66, 8),
33922 => conv_std_logic_vector(67, 8),
33923 => conv_std_logic_vector(67, 8),
33924 => conv_std_logic_vector(68, 8),
33925 => conv_std_logic_vector(68, 8),
33926 => conv_std_logic_vector(69, 8),
33927 => conv_std_logic_vector(69, 8),
33928 => conv_std_logic_vector(70, 8),
33929 => conv_std_logic_vector(70, 8),
33930 => conv_std_logic_vector(71, 8),
33931 => conv_std_logic_vector(71, 8),
33932 => conv_std_logic_vector(72, 8),
33933 => conv_std_logic_vector(72, 8),
33934 => conv_std_logic_vector(73, 8),
33935 => conv_std_logic_vector(73, 8),
33936 => conv_std_logic_vector(74, 8),
33937 => conv_std_logic_vector(74, 8),
33938 => conv_std_logic_vector(75, 8),
33939 => conv_std_logic_vector(75, 8),
33940 => conv_std_logic_vector(76, 8),
33941 => conv_std_logic_vector(76, 8),
33942 => conv_std_logic_vector(77, 8),
33943 => conv_std_logic_vector(77, 8),
33944 => conv_std_logic_vector(78, 8),
33945 => conv_std_logic_vector(78, 8),
33946 => conv_std_logic_vector(79, 8),
33947 => conv_std_logic_vector(79, 8),
33948 => conv_std_logic_vector(80, 8),
33949 => conv_std_logic_vector(80, 8),
33950 => conv_std_logic_vector(81, 8),
33951 => conv_std_logic_vector(81, 8),
33952 => conv_std_logic_vector(82, 8),
33953 => conv_std_logic_vector(83, 8),
33954 => conv_std_logic_vector(83, 8),
33955 => conv_std_logic_vector(84, 8),
33956 => conv_std_logic_vector(84, 8),
33957 => conv_std_logic_vector(85, 8),
33958 => conv_std_logic_vector(85, 8),
33959 => conv_std_logic_vector(86, 8),
33960 => conv_std_logic_vector(86, 8),
33961 => conv_std_logic_vector(87, 8),
33962 => conv_std_logic_vector(87, 8),
33963 => conv_std_logic_vector(88, 8),
33964 => conv_std_logic_vector(88, 8),
33965 => conv_std_logic_vector(89, 8),
33966 => conv_std_logic_vector(89, 8),
33967 => conv_std_logic_vector(90, 8),
33968 => conv_std_logic_vector(90, 8),
33969 => conv_std_logic_vector(91, 8),
33970 => conv_std_logic_vector(91, 8),
33971 => conv_std_logic_vector(92, 8),
33972 => conv_std_logic_vector(92, 8),
33973 => conv_std_logic_vector(93, 8),
33974 => conv_std_logic_vector(93, 8),
33975 => conv_std_logic_vector(94, 8),
33976 => conv_std_logic_vector(94, 8),
33977 => conv_std_logic_vector(95, 8),
33978 => conv_std_logic_vector(95, 8),
33979 => conv_std_logic_vector(96, 8),
33980 => conv_std_logic_vector(96, 8),
33981 => conv_std_logic_vector(97, 8),
33982 => conv_std_logic_vector(97, 8),
33983 => conv_std_logic_vector(98, 8),
33984 => conv_std_logic_vector(99, 8),
33985 => conv_std_logic_vector(99, 8),
33986 => conv_std_logic_vector(100, 8),
33987 => conv_std_logic_vector(100, 8),
33988 => conv_std_logic_vector(101, 8),
33989 => conv_std_logic_vector(101, 8),
33990 => conv_std_logic_vector(102, 8),
33991 => conv_std_logic_vector(102, 8),
33992 => conv_std_logic_vector(103, 8),
33993 => conv_std_logic_vector(103, 8),
33994 => conv_std_logic_vector(104, 8),
33995 => conv_std_logic_vector(104, 8),
33996 => conv_std_logic_vector(105, 8),
33997 => conv_std_logic_vector(105, 8),
33998 => conv_std_logic_vector(106, 8),
33999 => conv_std_logic_vector(106, 8),
34000 => conv_std_logic_vector(107, 8),
34001 => conv_std_logic_vector(107, 8),
34002 => conv_std_logic_vector(108, 8),
34003 => conv_std_logic_vector(108, 8),
34004 => conv_std_logic_vector(109, 8),
34005 => conv_std_logic_vector(109, 8),
34006 => conv_std_logic_vector(110, 8),
34007 => conv_std_logic_vector(110, 8),
34008 => conv_std_logic_vector(111, 8),
34009 => conv_std_logic_vector(111, 8),
34010 => conv_std_logic_vector(112, 8),
34011 => conv_std_logic_vector(112, 8),
34012 => conv_std_logic_vector(113, 8),
34013 => conv_std_logic_vector(113, 8),
34014 => conv_std_logic_vector(114, 8),
34015 => conv_std_logic_vector(114, 8),
34016 => conv_std_logic_vector(115, 8),
34017 => conv_std_logic_vector(116, 8),
34018 => conv_std_logic_vector(116, 8),
34019 => conv_std_logic_vector(117, 8),
34020 => conv_std_logic_vector(117, 8),
34021 => conv_std_logic_vector(118, 8),
34022 => conv_std_logic_vector(118, 8),
34023 => conv_std_logic_vector(119, 8),
34024 => conv_std_logic_vector(119, 8),
34025 => conv_std_logic_vector(120, 8),
34026 => conv_std_logic_vector(120, 8),
34027 => conv_std_logic_vector(121, 8),
34028 => conv_std_logic_vector(121, 8),
34029 => conv_std_logic_vector(122, 8),
34030 => conv_std_logic_vector(122, 8),
34031 => conv_std_logic_vector(123, 8),
34032 => conv_std_logic_vector(123, 8),
34033 => conv_std_logic_vector(124, 8),
34034 => conv_std_logic_vector(124, 8),
34035 => conv_std_logic_vector(125, 8),
34036 => conv_std_logic_vector(125, 8),
34037 => conv_std_logic_vector(126, 8),
34038 => conv_std_logic_vector(126, 8),
34039 => conv_std_logic_vector(127, 8),
34040 => conv_std_logic_vector(127, 8),
34041 => conv_std_logic_vector(128, 8),
34042 => conv_std_logic_vector(128, 8),
34043 => conv_std_logic_vector(129, 8),
34044 => conv_std_logic_vector(129, 8),
34045 => conv_std_logic_vector(130, 8),
34046 => conv_std_logic_vector(130, 8),
34047 => conv_std_logic_vector(131, 8),
34048 => conv_std_logic_vector(0, 8),
34049 => conv_std_logic_vector(0, 8),
34050 => conv_std_logic_vector(1, 8),
34051 => conv_std_logic_vector(1, 8),
34052 => conv_std_logic_vector(2, 8),
34053 => conv_std_logic_vector(2, 8),
34054 => conv_std_logic_vector(3, 8),
34055 => conv_std_logic_vector(3, 8),
34056 => conv_std_logic_vector(4, 8),
34057 => conv_std_logic_vector(4, 8),
34058 => conv_std_logic_vector(5, 8),
34059 => conv_std_logic_vector(5, 8),
34060 => conv_std_logic_vector(6, 8),
34061 => conv_std_logic_vector(6, 8),
34062 => conv_std_logic_vector(7, 8),
34063 => conv_std_logic_vector(7, 8),
34064 => conv_std_logic_vector(8, 8),
34065 => conv_std_logic_vector(8, 8),
34066 => conv_std_logic_vector(9, 8),
34067 => conv_std_logic_vector(9, 8),
34068 => conv_std_logic_vector(10, 8),
34069 => conv_std_logic_vector(10, 8),
34070 => conv_std_logic_vector(11, 8),
34071 => conv_std_logic_vector(11, 8),
34072 => conv_std_logic_vector(12, 8),
34073 => conv_std_logic_vector(12, 8),
34074 => conv_std_logic_vector(13, 8),
34075 => conv_std_logic_vector(14, 8),
34076 => conv_std_logic_vector(14, 8),
34077 => conv_std_logic_vector(15, 8),
34078 => conv_std_logic_vector(15, 8),
34079 => conv_std_logic_vector(16, 8),
34080 => conv_std_logic_vector(16, 8),
34081 => conv_std_logic_vector(17, 8),
34082 => conv_std_logic_vector(17, 8),
34083 => conv_std_logic_vector(18, 8),
34084 => conv_std_logic_vector(18, 8),
34085 => conv_std_logic_vector(19, 8),
34086 => conv_std_logic_vector(19, 8),
34087 => conv_std_logic_vector(20, 8),
34088 => conv_std_logic_vector(20, 8),
34089 => conv_std_logic_vector(21, 8),
34090 => conv_std_logic_vector(21, 8),
34091 => conv_std_logic_vector(22, 8),
34092 => conv_std_logic_vector(22, 8),
34093 => conv_std_logic_vector(23, 8),
34094 => conv_std_logic_vector(23, 8),
34095 => conv_std_logic_vector(24, 8),
34096 => conv_std_logic_vector(24, 8),
34097 => conv_std_logic_vector(25, 8),
34098 => conv_std_logic_vector(25, 8),
34099 => conv_std_logic_vector(26, 8),
34100 => conv_std_logic_vector(27, 8),
34101 => conv_std_logic_vector(27, 8),
34102 => conv_std_logic_vector(28, 8),
34103 => conv_std_logic_vector(28, 8),
34104 => conv_std_logic_vector(29, 8),
34105 => conv_std_logic_vector(29, 8),
34106 => conv_std_logic_vector(30, 8),
34107 => conv_std_logic_vector(30, 8),
34108 => conv_std_logic_vector(31, 8),
34109 => conv_std_logic_vector(31, 8),
34110 => conv_std_logic_vector(32, 8),
34111 => conv_std_logic_vector(32, 8),
34112 => conv_std_logic_vector(33, 8),
34113 => conv_std_logic_vector(33, 8),
34114 => conv_std_logic_vector(34, 8),
34115 => conv_std_logic_vector(34, 8),
34116 => conv_std_logic_vector(35, 8),
34117 => conv_std_logic_vector(35, 8),
34118 => conv_std_logic_vector(36, 8),
34119 => conv_std_logic_vector(36, 8),
34120 => conv_std_logic_vector(37, 8),
34121 => conv_std_logic_vector(37, 8),
34122 => conv_std_logic_vector(38, 8),
34123 => conv_std_logic_vector(38, 8),
34124 => conv_std_logic_vector(39, 8),
34125 => conv_std_logic_vector(40, 8),
34126 => conv_std_logic_vector(40, 8),
34127 => conv_std_logic_vector(41, 8),
34128 => conv_std_logic_vector(41, 8),
34129 => conv_std_logic_vector(42, 8),
34130 => conv_std_logic_vector(42, 8),
34131 => conv_std_logic_vector(43, 8),
34132 => conv_std_logic_vector(43, 8),
34133 => conv_std_logic_vector(44, 8),
34134 => conv_std_logic_vector(44, 8),
34135 => conv_std_logic_vector(45, 8),
34136 => conv_std_logic_vector(45, 8),
34137 => conv_std_logic_vector(46, 8),
34138 => conv_std_logic_vector(46, 8),
34139 => conv_std_logic_vector(47, 8),
34140 => conv_std_logic_vector(47, 8),
34141 => conv_std_logic_vector(48, 8),
34142 => conv_std_logic_vector(48, 8),
34143 => conv_std_logic_vector(49, 8),
34144 => conv_std_logic_vector(49, 8),
34145 => conv_std_logic_vector(50, 8),
34146 => conv_std_logic_vector(50, 8),
34147 => conv_std_logic_vector(51, 8),
34148 => conv_std_logic_vector(51, 8),
34149 => conv_std_logic_vector(52, 8),
34150 => conv_std_logic_vector(52, 8),
34151 => conv_std_logic_vector(53, 8),
34152 => conv_std_logic_vector(54, 8),
34153 => conv_std_logic_vector(54, 8),
34154 => conv_std_logic_vector(55, 8),
34155 => conv_std_logic_vector(55, 8),
34156 => conv_std_logic_vector(56, 8),
34157 => conv_std_logic_vector(56, 8),
34158 => conv_std_logic_vector(57, 8),
34159 => conv_std_logic_vector(57, 8),
34160 => conv_std_logic_vector(58, 8),
34161 => conv_std_logic_vector(58, 8),
34162 => conv_std_logic_vector(59, 8),
34163 => conv_std_logic_vector(59, 8),
34164 => conv_std_logic_vector(60, 8),
34165 => conv_std_logic_vector(60, 8),
34166 => conv_std_logic_vector(61, 8),
34167 => conv_std_logic_vector(61, 8),
34168 => conv_std_logic_vector(62, 8),
34169 => conv_std_logic_vector(62, 8),
34170 => conv_std_logic_vector(63, 8),
34171 => conv_std_logic_vector(63, 8),
34172 => conv_std_logic_vector(64, 8),
34173 => conv_std_logic_vector(64, 8),
34174 => conv_std_logic_vector(65, 8),
34175 => conv_std_logic_vector(65, 8),
34176 => conv_std_logic_vector(66, 8),
34177 => conv_std_logic_vector(67, 8),
34178 => conv_std_logic_vector(67, 8),
34179 => conv_std_logic_vector(68, 8),
34180 => conv_std_logic_vector(68, 8),
34181 => conv_std_logic_vector(69, 8),
34182 => conv_std_logic_vector(69, 8),
34183 => conv_std_logic_vector(70, 8),
34184 => conv_std_logic_vector(70, 8),
34185 => conv_std_logic_vector(71, 8),
34186 => conv_std_logic_vector(71, 8),
34187 => conv_std_logic_vector(72, 8),
34188 => conv_std_logic_vector(72, 8),
34189 => conv_std_logic_vector(73, 8),
34190 => conv_std_logic_vector(73, 8),
34191 => conv_std_logic_vector(74, 8),
34192 => conv_std_logic_vector(74, 8),
34193 => conv_std_logic_vector(75, 8),
34194 => conv_std_logic_vector(75, 8),
34195 => conv_std_logic_vector(76, 8),
34196 => conv_std_logic_vector(76, 8),
34197 => conv_std_logic_vector(77, 8),
34198 => conv_std_logic_vector(77, 8),
34199 => conv_std_logic_vector(78, 8),
34200 => conv_std_logic_vector(78, 8),
34201 => conv_std_logic_vector(79, 8),
34202 => conv_std_logic_vector(80, 8),
34203 => conv_std_logic_vector(80, 8),
34204 => conv_std_logic_vector(81, 8),
34205 => conv_std_logic_vector(81, 8),
34206 => conv_std_logic_vector(82, 8),
34207 => conv_std_logic_vector(82, 8),
34208 => conv_std_logic_vector(83, 8),
34209 => conv_std_logic_vector(83, 8),
34210 => conv_std_logic_vector(84, 8),
34211 => conv_std_logic_vector(84, 8),
34212 => conv_std_logic_vector(85, 8),
34213 => conv_std_logic_vector(85, 8),
34214 => conv_std_logic_vector(86, 8),
34215 => conv_std_logic_vector(86, 8),
34216 => conv_std_logic_vector(87, 8),
34217 => conv_std_logic_vector(87, 8),
34218 => conv_std_logic_vector(88, 8),
34219 => conv_std_logic_vector(88, 8),
34220 => conv_std_logic_vector(89, 8),
34221 => conv_std_logic_vector(89, 8),
34222 => conv_std_logic_vector(90, 8),
34223 => conv_std_logic_vector(90, 8),
34224 => conv_std_logic_vector(91, 8),
34225 => conv_std_logic_vector(91, 8),
34226 => conv_std_logic_vector(92, 8),
34227 => conv_std_logic_vector(92, 8),
34228 => conv_std_logic_vector(93, 8),
34229 => conv_std_logic_vector(94, 8),
34230 => conv_std_logic_vector(94, 8),
34231 => conv_std_logic_vector(95, 8),
34232 => conv_std_logic_vector(95, 8),
34233 => conv_std_logic_vector(96, 8),
34234 => conv_std_logic_vector(96, 8),
34235 => conv_std_logic_vector(97, 8),
34236 => conv_std_logic_vector(97, 8),
34237 => conv_std_logic_vector(98, 8),
34238 => conv_std_logic_vector(98, 8),
34239 => conv_std_logic_vector(99, 8),
34240 => conv_std_logic_vector(99, 8),
34241 => conv_std_logic_vector(100, 8),
34242 => conv_std_logic_vector(100, 8),
34243 => conv_std_logic_vector(101, 8),
34244 => conv_std_logic_vector(101, 8),
34245 => conv_std_logic_vector(102, 8),
34246 => conv_std_logic_vector(102, 8),
34247 => conv_std_logic_vector(103, 8),
34248 => conv_std_logic_vector(103, 8),
34249 => conv_std_logic_vector(104, 8),
34250 => conv_std_logic_vector(104, 8),
34251 => conv_std_logic_vector(105, 8),
34252 => conv_std_logic_vector(105, 8),
34253 => conv_std_logic_vector(106, 8),
34254 => conv_std_logic_vector(107, 8),
34255 => conv_std_logic_vector(107, 8),
34256 => conv_std_logic_vector(108, 8),
34257 => conv_std_logic_vector(108, 8),
34258 => conv_std_logic_vector(109, 8),
34259 => conv_std_logic_vector(109, 8),
34260 => conv_std_logic_vector(110, 8),
34261 => conv_std_logic_vector(110, 8),
34262 => conv_std_logic_vector(111, 8),
34263 => conv_std_logic_vector(111, 8),
34264 => conv_std_logic_vector(112, 8),
34265 => conv_std_logic_vector(112, 8),
34266 => conv_std_logic_vector(113, 8),
34267 => conv_std_logic_vector(113, 8),
34268 => conv_std_logic_vector(114, 8),
34269 => conv_std_logic_vector(114, 8),
34270 => conv_std_logic_vector(115, 8),
34271 => conv_std_logic_vector(115, 8),
34272 => conv_std_logic_vector(116, 8),
34273 => conv_std_logic_vector(116, 8),
34274 => conv_std_logic_vector(117, 8),
34275 => conv_std_logic_vector(117, 8),
34276 => conv_std_logic_vector(118, 8),
34277 => conv_std_logic_vector(118, 8),
34278 => conv_std_logic_vector(119, 8),
34279 => conv_std_logic_vector(120, 8),
34280 => conv_std_logic_vector(120, 8),
34281 => conv_std_logic_vector(121, 8),
34282 => conv_std_logic_vector(121, 8),
34283 => conv_std_logic_vector(122, 8),
34284 => conv_std_logic_vector(122, 8),
34285 => conv_std_logic_vector(123, 8),
34286 => conv_std_logic_vector(123, 8),
34287 => conv_std_logic_vector(124, 8),
34288 => conv_std_logic_vector(124, 8),
34289 => conv_std_logic_vector(125, 8),
34290 => conv_std_logic_vector(125, 8),
34291 => conv_std_logic_vector(126, 8),
34292 => conv_std_logic_vector(126, 8),
34293 => conv_std_logic_vector(127, 8),
34294 => conv_std_logic_vector(127, 8),
34295 => conv_std_logic_vector(128, 8),
34296 => conv_std_logic_vector(128, 8),
34297 => conv_std_logic_vector(129, 8),
34298 => conv_std_logic_vector(129, 8),
34299 => conv_std_logic_vector(130, 8),
34300 => conv_std_logic_vector(130, 8),
34301 => conv_std_logic_vector(131, 8),
34302 => conv_std_logic_vector(131, 8),
34303 => conv_std_logic_vector(132, 8),
34304 => conv_std_logic_vector(0, 8),
34305 => conv_std_logic_vector(0, 8),
34306 => conv_std_logic_vector(1, 8),
34307 => conv_std_logic_vector(1, 8),
34308 => conv_std_logic_vector(2, 8),
34309 => conv_std_logic_vector(2, 8),
34310 => conv_std_logic_vector(3, 8),
34311 => conv_std_logic_vector(3, 8),
34312 => conv_std_logic_vector(4, 8),
34313 => conv_std_logic_vector(4, 8),
34314 => conv_std_logic_vector(5, 8),
34315 => conv_std_logic_vector(5, 8),
34316 => conv_std_logic_vector(6, 8),
34317 => conv_std_logic_vector(6, 8),
34318 => conv_std_logic_vector(7, 8),
34319 => conv_std_logic_vector(7, 8),
34320 => conv_std_logic_vector(8, 8),
34321 => conv_std_logic_vector(8, 8),
34322 => conv_std_logic_vector(9, 8),
34323 => conv_std_logic_vector(9, 8),
34324 => conv_std_logic_vector(10, 8),
34325 => conv_std_logic_vector(10, 8),
34326 => conv_std_logic_vector(11, 8),
34327 => conv_std_logic_vector(12, 8),
34328 => conv_std_logic_vector(12, 8),
34329 => conv_std_logic_vector(13, 8),
34330 => conv_std_logic_vector(13, 8),
34331 => conv_std_logic_vector(14, 8),
34332 => conv_std_logic_vector(14, 8),
34333 => conv_std_logic_vector(15, 8),
34334 => conv_std_logic_vector(15, 8),
34335 => conv_std_logic_vector(16, 8),
34336 => conv_std_logic_vector(16, 8),
34337 => conv_std_logic_vector(17, 8),
34338 => conv_std_logic_vector(17, 8),
34339 => conv_std_logic_vector(18, 8),
34340 => conv_std_logic_vector(18, 8),
34341 => conv_std_logic_vector(19, 8),
34342 => conv_std_logic_vector(19, 8),
34343 => conv_std_logic_vector(20, 8),
34344 => conv_std_logic_vector(20, 8),
34345 => conv_std_logic_vector(21, 8),
34346 => conv_std_logic_vector(21, 8),
34347 => conv_std_logic_vector(22, 8),
34348 => conv_std_logic_vector(23, 8),
34349 => conv_std_logic_vector(23, 8),
34350 => conv_std_logic_vector(24, 8),
34351 => conv_std_logic_vector(24, 8),
34352 => conv_std_logic_vector(25, 8),
34353 => conv_std_logic_vector(25, 8),
34354 => conv_std_logic_vector(26, 8),
34355 => conv_std_logic_vector(26, 8),
34356 => conv_std_logic_vector(27, 8),
34357 => conv_std_logic_vector(27, 8),
34358 => conv_std_logic_vector(28, 8),
34359 => conv_std_logic_vector(28, 8),
34360 => conv_std_logic_vector(29, 8),
34361 => conv_std_logic_vector(29, 8),
34362 => conv_std_logic_vector(30, 8),
34363 => conv_std_logic_vector(30, 8),
34364 => conv_std_logic_vector(31, 8),
34365 => conv_std_logic_vector(31, 8),
34366 => conv_std_logic_vector(32, 8),
34367 => conv_std_logic_vector(32, 8),
34368 => conv_std_logic_vector(33, 8),
34369 => conv_std_logic_vector(34, 8),
34370 => conv_std_logic_vector(34, 8),
34371 => conv_std_logic_vector(35, 8),
34372 => conv_std_logic_vector(35, 8),
34373 => conv_std_logic_vector(36, 8),
34374 => conv_std_logic_vector(36, 8),
34375 => conv_std_logic_vector(37, 8),
34376 => conv_std_logic_vector(37, 8),
34377 => conv_std_logic_vector(38, 8),
34378 => conv_std_logic_vector(38, 8),
34379 => conv_std_logic_vector(39, 8),
34380 => conv_std_logic_vector(39, 8),
34381 => conv_std_logic_vector(40, 8),
34382 => conv_std_logic_vector(40, 8),
34383 => conv_std_logic_vector(41, 8),
34384 => conv_std_logic_vector(41, 8),
34385 => conv_std_logic_vector(42, 8),
34386 => conv_std_logic_vector(42, 8),
34387 => conv_std_logic_vector(43, 8),
34388 => conv_std_logic_vector(43, 8),
34389 => conv_std_logic_vector(44, 8),
34390 => conv_std_logic_vector(45, 8),
34391 => conv_std_logic_vector(45, 8),
34392 => conv_std_logic_vector(46, 8),
34393 => conv_std_logic_vector(46, 8),
34394 => conv_std_logic_vector(47, 8),
34395 => conv_std_logic_vector(47, 8),
34396 => conv_std_logic_vector(48, 8),
34397 => conv_std_logic_vector(48, 8),
34398 => conv_std_logic_vector(49, 8),
34399 => conv_std_logic_vector(49, 8),
34400 => conv_std_logic_vector(50, 8),
34401 => conv_std_logic_vector(50, 8),
34402 => conv_std_logic_vector(51, 8),
34403 => conv_std_logic_vector(51, 8),
34404 => conv_std_logic_vector(52, 8),
34405 => conv_std_logic_vector(52, 8),
34406 => conv_std_logic_vector(53, 8),
34407 => conv_std_logic_vector(53, 8),
34408 => conv_std_logic_vector(54, 8),
34409 => conv_std_logic_vector(54, 8),
34410 => conv_std_logic_vector(55, 8),
34411 => conv_std_logic_vector(56, 8),
34412 => conv_std_logic_vector(56, 8),
34413 => conv_std_logic_vector(57, 8),
34414 => conv_std_logic_vector(57, 8),
34415 => conv_std_logic_vector(58, 8),
34416 => conv_std_logic_vector(58, 8),
34417 => conv_std_logic_vector(59, 8),
34418 => conv_std_logic_vector(59, 8),
34419 => conv_std_logic_vector(60, 8),
34420 => conv_std_logic_vector(60, 8),
34421 => conv_std_logic_vector(61, 8),
34422 => conv_std_logic_vector(61, 8),
34423 => conv_std_logic_vector(62, 8),
34424 => conv_std_logic_vector(62, 8),
34425 => conv_std_logic_vector(63, 8),
34426 => conv_std_logic_vector(63, 8),
34427 => conv_std_logic_vector(64, 8),
34428 => conv_std_logic_vector(64, 8),
34429 => conv_std_logic_vector(65, 8),
34430 => conv_std_logic_vector(65, 8),
34431 => conv_std_logic_vector(66, 8),
34432 => conv_std_logic_vector(67, 8),
34433 => conv_std_logic_vector(67, 8),
34434 => conv_std_logic_vector(68, 8),
34435 => conv_std_logic_vector(68, 8),
34436 => conv_std_logic_vector(69, 8),
34437 => conv_std_logic_vector(69, 8),
34438 => conv_std_logic_vector(70, 8),
34439 => conv_std_logic_vector(70, 8),
34440 => conv_std_logic_vector(71, 8),
34441 => conv_std_logic_vector(71, 8),
34442 => conv_std_logic_vector(72, 8),
34443 => conv_std_logic_vector(72, 8),
34444 => conv_std_logic_vector(73, 8),
34445 => conv_std_logic_vector(73, 8),
34446 => conv_std_logic_vector(74, 8),
34447 => conv_std_logic_vector(74, 8),
34448 => conv_std_logic_vector(75, 8),
34449 => conv_std_logic_vector(75, 8),
34450 => conv_std_logic_vector(76, 8),
34451 => conv_std_logic_vector(76, 8),
34452 => conv_std_logic_vector(77, 8),
34453 => conv_std_logic_vector(77, 8),
34454 => conv_std_logic_vector(78, 8),
34455 => conv_std_logic_vector(79, 8),
34456 => conv_std_logic_vector(79, 8),
34457 => conv_std_logic_vector(80, 8),
34458 => conv_std_logic_vector(80, 8),
34459 => conv_std_logic_vector(81, 8),
34460 => conv_std_logic_vector(81, 8),
34461 => conv_std_logic_vector(82, 8),
34462 => conv_std_logic_vector(82, 8),
34463 => conv_std_logic_vector(83, 8),
34464 => conv_std_logic_vector(83, 8),
34465 => conv_std_logic_vector(84, 8),
34466 => conv_std_logic_vector(84, 8),
34467 => conv_std_logic_vector(85, 8),
34468 => conv_std_logic_vector(85, 8),
34469 => conv_std_logic_vector(86, 8),
34470 => conv_std_logic_vector(86, 8),
34471 => conv_std_logic_vector(87, 8),
34472 => conv_std_logic_vector(87, 8),
34473 => conv_std_logic_vector(88, 8),
34474 => conv_std_logic_vector(88, 8),
34475 => conv_std_logic_vector(89, 8),
34476 => conv_std_logic_vector(90, 8),
34477 => conv_std_logic_vector(90, 8),
34478 => conv_std_logic_vector(91, 8),
34479 => conv_std_logic_vector(91, 8),
34480 => conv_std_logic_vector(92, 8),
34481 => conv_std_logic_vector(92, 8),
34482 => conv_std_logic_vector(93, 8),
34483 => conv_std_logic_vector(93, 8),
34484 => conv_std_logic_vector(94, 8),
34485 => conv_std_logic_vector(94, 8),
34486 => conv_std_logic_vector(95, 8),
34487 => conv_std_logic_vector(95, 8),
34488 => conv_std_logic_vector(96, 8),
34489 => conv_std_logic_vector(96, 8),
34490 => conv_std_logic_vector(97, 8),
34491 => conv_std_logic_vector(97, 8),
34492 => conv_std_logic_vector(98, 8),
34493 => conv_std_logic_vector(98, 8),
34494 => conv_std_logic_vector(99, 8),
34495 => conv_std_logic_vector(99, 8),
34496 => conv_std_logic_vector(100, 8),
34497 => conv_std_logic_vector(101, 8),
34498 => conv_std_logic_vector(101, 8),
34499 => conv_std_logic_vector(102, 8),
34500 => conv_std_logic_vector(102, 8),
34501 => conv_std_logic_vector(103, 8),
34502 => conv_std_logic_vector(103, 8),
34503 => conv_std_logic_vector(104, 8),
34504 => conv_std_logic_vector(104, 8),
34505 => conv_std_logic_vector(105, 8),
34506 => conv_std_logic_vector(105, 8),
34507 => conv_std_logic_vector(106, 8),
34508 => conv_std_logic_vector(106, 8),
34509 => conv_std_logic_vector(107, 8),
34510 => conv_std_logic_vector(107, 8),
34511 => conv_std_logic_vector(108, 8),
34512 => conv_std_logic_vector(108, 8),
34513 => conv_std_logic_vector(109, 8),
34514 => conv_std_logic_vector(109, 8),
34515 => conv_std_logic_vector(110, 8),
34516 => conv_std_logic_vector(110, 8),
34517 => conv_std_logic_vector(111, 8),
34518 => conv_std_logic_vector(112, 8),
34519 => conv_std_logic_vector(112, 8),
34520 => conv_std_logic_vector(113, 8),
34521 => conv_std_logic_vector(113, 8),
34522 => conv_std_logic_vector(114, 8),
34523 => conv_std_logic_vector(114, 8),
34524 => conv_std_logic_vector(115, 8),
34525 => conv_std_logic_vector(115, 8),
34526 => conv_std_logic_vector(116, 8),
34527 => conv_std_logic_vector(116, 8),
34528 => conv_std_logic_vector(117, 8),
34529 => conv_std_logic_vector(117, 8),
34530 => conv_std_logic_vector(118, 8),
34531 => conv_std_logic_vector(118, 8),
34532 => conv_std_logic_vector(119, 8),
34533 => conv_std_logic_vector(119, 8),
34534 => conv_std_logic_vector(120, 8),
34535 => conv_std_logic_vector(120, 8),
34536 => conv_std_logic_vector(121, 8),
34537 => conv_std_logic_vector(121, 8),
34538 => conv_std_logic_vector(122, 8),
34539 => conv_std_logic_vector(123, 8),
34540 => conv_std_logic_vector(123, 8),
34541 => conv_std_logic_vector(124, 8),
34542 => conv_std_logic_vector(124, 8),
34543 => conv_std_logic_vector(125, 8),
34544 => conv_std_logic_vector(125, 8),
34545 => conv_std_logic_vector(126, 8),
34546 => conv_std_logic_vector(126, 8),
34547 => conv_std_logic_vector(127, 8),
34548 => conv_std_logic_vector(127, 8),
34549 => conv_std_logic_vector(128, 8),
34550 => conv_std_logic_vector(128, 8),
34551 => conv_std_logic_vector(129, 8),
34552 => conv_std_logic_vector(129, 8),
34553 => conv_std_logic_vector(130, 8),
34554 => conv_std_logic_vector(130, 8),
34555 => conv_std_logic_vector(131, 8),
34556 => conv_std_logic_vector(131, 8),
34557 => conv_std_logic_vector(132, 8),
34558 => conv_std_logic_vector(132, 8),
34559 => conv_std_logic_vector(133, 8),
34560 => conv_std_logic_vector(0, 8),
34561 => conv_std_logic_vector(0, 8),
34562 => conv_std_logic_vector(1, 8),
34563 => conv_std_logic_vector(1, 8),
34564 => conv_std_logic_vector(2, 8),
34565 => conv_std_logic_vector(2, 8),
34566 => conv_std_logic_vector(3, 8),
34567 => conv_std_logic_vector(3, 8),
34568 => conv_std_logic_vector(4, 8),
34569 => conv_std_logic_vector(4, 8),
34570 => conv_std_logic_vector(5, 8),
34571 => conv_std_logic_vector(5, 8),
34572 => conv_std_logic_vector(6, 8),
34573 => conv_std_logic_vector(6, 8),
34574 => conv_std_logic_vector(7, 8),
34575 => conv_std_logic_vector(7, 8),
34576 => conv_std_logic_vector(8, 8),
34577 => conv_std_logic_vector(8, 8),
34578 => conv_std_logic_vector(9, 8),
34579 => conv_std_logic_vector(10, 8),
34580 => conv_std_logic_vector(10, 8),
34581 => conv_std_logic_vector(11, 8),
34582 => conv_std_logic_vector(11, 8),
34583 => conv_std_logic_vector(12, 8),
34584 => conv_std_logic_vector(12, 8),
34585 => conv_std_logic_vector(13, 8),
34586 => conv_std_logic_vector(13, 8),
34587 => conv_std_logic_vector(14, 8),
34588 => conv_std_logic_vector(14, 8),
34589 => conv_std_logic_vector(15, 8),
34590 => conv_std_logic_vector(15, 8),
34591 => conv_std_logic_vector(16, 8),
34592 => conv_std_logic_vector(16, 8),
34593 => conv_std_logic_vector(17, 8),
34594 => conv_std_logic_vector(17, 8),
34595 => conv_std_logic_vector(18, 8),
34596 => conv_std_logic_vector(18, 8),
34597 => conv_std_logic_vector(19, 8),
34598 => conv_std_logic_vector(20, 8),
34599 => conv_std_logic_vector(20, 8),
34600 => conv_std_logic_vector(21, 8),
34601 => conv_std_logic_vector(21, 8),
34602 => conv_std_logic_vector(22, 8),
34603 => conv_std_logic_vector(22, 8),
34604 => conv_std_logic_vector(23, 8),
34605 => conv_std_logic_vector(23, 8),
34606 => conv_std_logic_vector(24, 8),
34607 => conv_std_logic_vector(24, 8),
34608 => conv_std_logic_vector(25, 8),
34609 => conv_std_logic_vector(25, 8),
34610 => conv_std_logic_vector(26, 8),
34611 => conv_std_logic_vector(26, 8),
34612 => conv_std_logic_vector(27, 8),
34613 => conv_std_logic_vector(27, 8),
34614 => conv_std_logic_vector(28, 8),
34615 => conv_std_logic_vector(29, 8),
34616 => conv_std_logic_vector(29, 8),
34617 => conv_std_logic_vector(30, 8),
34618 => conv_std_logic_vector(30, 8),
34619 => conv_std_logic_vector(31, 8),
34620 => conv_std_logic_vector(31, 8),
34621 => conv_std_logic_vector(32, 8),
34622 => conv_std_logic_vector(32, 8),
34623 => conv_std_logic_vector(33, 8),
34624 => conv_std_logic_vector(33, 8),
34625 => conv_std_logic_vector(34, 8),
34626 => conv_std_logic_vector(34, 8),
34627 => conv_std_logic_vector(35, 8),
34628 => conv_std_logic_vector(35, 8),
34629 => conv_std_logic_vector(36, 8),
34630 => conv_std_logic_vector(36, 8),
34631 => conv_std_logic_vector(37, 8),
34632 => conv_std_logic_vector(37, 8),
34633 => conv_std_logic_vector(38, 8),
34634 => conv_std_logic_vector(39, 8),
34635 => conv_std_logic_vector(39, 8),
34636 => conv_std_logic_vector(40, 8),
34637 => conv_std_logic_vector(40, 8),
34638 => conv_std_logic_vector(41, 8),
34639 => conv_std_logic_vector(41, 8),
34640 => conv_std_logic_vector(42, 8),
34641 => conv_std_logic_vector(42, 8),
34642 => conv_std_logic_vector(43, 8),
34643 => conv_std_logic_vector(43, 8),
34644 => conv_std_logic_vector(44, 8),
34645 => conv_std_logic_vector(44, 8),
34646 => conv_std_logic_vector(45, 8),
34647 => conv_std_logic_vector(45, 8),
34648 => conv_std_logic_vector(46, 8),
34649 => conv_std_logic_vector(46, 8),
34650 => conv_std_logic_vector(47, 8),
34651 => conv_std_logic_vector(47, 8),
34652 => conv_std_logic_vector(48, 8),
34653 => conv_std_logic_vector(49, 8),
34654 => conv_std_logic_vector(49, 8),
34655 => conv_std_logic_vector(50, 8),
34656 => conv_std_logic_vector(50, 8),
34657 => conv_std_logic_vector(51, 8),
34658 => conv_std_logic_vector(51, 8),
34659 => conv_std_logic_vector(52, 8),
34660 => conv_std_logic_vector(52, 8),
34661 => conv_std_logic_vector(53, 8),
34662 => conv_std_logic_vector(53, 8),
34663 => conv_std_logic_vector(54, 8),
34664 => conv_std_logic_vector(54, 8),
34665 => conv_std_logic_vector(55, 8),
34666 => conv_std_logic_vector(55, 8),
34667 => conv_std_logic_vector(56, 8),
34668 => conv_std_logic_vector(56, 8),
34669 => conv_std_logic_vector(57, 8),
34670 => conv_std_logic_vector(58, 8),
34671 => conv_std_logic_vector(58, 8),
34672 => conv_std_logic_vector(59, 8),
34673 => conv_std_logic_vector(59, 8),
34674 => conv_std_logic_vector(60, 8),
34675 => conv_std_logic_vector(60, 8),
34676 => conv_std_logic_vector(61, 8),
34677 => conv_std_logic_vector(61, 8),
34678 => conv_std_logic_vector(62, 8),
34679 => conv_std_logic_vector(62, 8),
34680 => conv_std_logic_vector(63, 8),
34681 => conv_std_logic_vector(63, 8),
34682 => conv_std_logic_vector(64, 8),
34683 => conv_std_logic_vector(64, 8),
34684 => conv_std_logic_vector(65, 8),
34685 => conv_std_logic_vector(65, 8),
34686 => conv_std_logic_vector(66, 8),
34687 => conv_std_logic_vector(66, 8),
34688 => conv_std_logic_vector(67, 8),
34689 => conv_std_logic_vector(68, 8),
34690 => conv_std_logic_vector(68, 8),
34691 => conv_std_logic_vector(69, 8),
34692 => conv_std_logic_vector(69, 8),
34693 => conv_std_logic_vector(70, 8),
34694 => conv_std_logic_vector(70, 8),
34695 => conv_std_logic_vector(71, 8),
34696 => conv_std_logic_vector(71, 8),
34697 => conv_std_logic_vector(72, 8),
34698 => conv_std_logic_vector(72, 8),
34699 => conv_std_logic_vector(73, 8),
34700 => conv_std_logic_vector(73, 8),
34701 => conv_std_logic_vector(74, 8),
34702 => conv_std_logic_vector(74, 8),
34703 => conv_std_logic_vector(75, 8),
34704 => conv_std_logic_vector(75, 8),
34705 => conv_std_logic_vector(76, 8),
34706 => conv_std_logic_vector(76, 8),
34707 => conv_std_logic_vector(77, 8),
34708 => conv_std_logic_vector(78, 8),
34709 => conv_std_logic_vector(78, 8),
34710 => conv_std_logic_vector(79, 8),
34711 => conv_std_logic_vector(79, 8),
34712 => conv_std_logic_vector(80, 8),
34713 => conv_std_logic_vector(80, 8),
34714 => conv_std_logic_vector(81, 8),
34715 => conv_std_logic_vector(81, 8),
34716 => conv_std_logic_vector(82, 8),
34717 => conv_std_logic_vector(82, 8),
34718 => conv_std_logic_vector(83, 8),
34719 => conv_std_logic_vector(83, 8),
34720 => conv_std_logic_vector(84, 8),
34721 => conv_std_logic_vector(84, 8),
34722 => conv_std_logic_vector(85, 8),
34723 => conv_std_logic_vector(85, 8),
34724 => conv_std_logic_vector(86, 8),
34725 => conv_std_logic_vector(87, 8),
34726 => conv_std_logic_vector(87, 8),
34727 => conv_std_logic_vector(88, 8),
34728 => conv_std_logic_vector(88, 8),
34729 => conv_std_logic_vector(89, 8),
34730 => conv_std_logic_vector(89, 8),
34731 => conv_std_logic_vector(90, 8),
34732 => conv_std_logic_vector(90, 8),
34733 => conv_std_logic_vector(91, 8),
34734 => conv_std_logic_vector(91, 8),
34735 => conv_std_logic_vector(92, 8),
34736 => conv_std_logic_vector(92, 8),
34737 => conv_std_logic_vector(93, 8),
34738 => conv_std_logic_vector(93, 8),
34739 => conv_std_logic_vector(94, 8),
34740 => conv_std_logic_vector(94, 8),
34741 => conv_std_logic_vector(95, 8),
34742 => conv_std_logic_vector(95, 8),
34743 => conv_std_logic_vector(96, 8),
34744 => conv_std_logic_vector(97, 8),
34745 => conv_std_logic_vector(97, 8),
34746 => conv_std_logic_vector(98, 8),
34747 => conv_std_logic_vector(98, 8),
34748 => conv_std_logic_vector(99, 8),
34749 => conv_std_logic_vector(99, 8),
34750 => conv_std_logic_vector(100, 8),
34751 => conv_std_logic_vector(100, 8),
34752 => conv_std_logic_vector(101, 8),
34753 => conv_std_logic_vector(101, 8),
34754 => conv_std_logic_vector(102, 8),
34755 => conv_std_logic_vector(102, 8),
34756 => conv_std_logic_vector(103, 8),
34757 => conv_std_logic_vector(103, 8),
34758 => conv_std_logic_vector(104, 8),
34759 => conv_std_logic_vector(104, 8),
34760 => conv_std_logic_vector(105, 8),
34761 => conv_std_logic_vector(105, 8),
34762 => conv_std_logic_vector(106, 8),
34763 => conv_std_logic_vector(107, 8),
34764 => conv_std_logic_vector(107, 8),
34765 => conv_std_logic_vector(108, 8),
34766 => conv_std_logic_vector(108, 8),
34767 => conv_std_logic_vector(109, 8),
34768 => conv_std_logic_vector(109, 8),
34769 => conv_std_logic_vector(110, 8),
34770 => conv_std_logic_vector(110, 8),
34771 => conv_std_logic_vector(111, 8),
34772 => conv_std_logic_vector(111, 8),
34773 => conv_std_logic_vector(112, 8),
34774 => conv_std_logic_vector(112, 8),
34775 => conv_std_logic_vector(113, 8),
34776 => conv_std_logic_vector(113, 8),
34777 => conv_std_logic_vector(114, 8),
34778 => conv_std_logic_vector(114, 8),
34779 => conv_std_logic_vector(115, 8),
34780 => conv_std_logic_vector(116, 8),
34781 => conv_std_logic_vector(116, 8),
34782 => conv_std_logic_vector(117, 8),
34783 => conv_std_logic_vector(117, 8),
34784 => conv_std_logic_vector(118, 8),
34785 => conv_std_logic_vector(118, 8),
34786 => conv_std_logic_vector(119, 8),
34787 => conv_std_logic_vector(119, 8),
34788 => conv_std_logic_vector(120, 8),
34789 => conv_std_logic_vector(120, 8),
34790 => conv_std_logic_vector(121, 8),
34791 => conv_std_logic_vector(121, 8),
34792 => conv_std_logic_vector(122, 8),
34793 => conv_std_logic_vector(122, 8),
34794 => conv_std_logic_vector(123, 8),
34795 => conv_std_logic_vector(123, 8),
34796 => conv_std_logic_vector(124, 8),
34797 => conv_std_logic_vector(124, 8),
34798 => conv_std_logic_vector(125, 8),
34799 => conv_std_logic_vector(126, 8),
34800 => conv_std_logic_vector(126, 8),
34801 => conv_std_logic_vector(127, 8),
34802 => conv_std_logic_vector(127, 8),
34803 => conv_std_logic_vector(128, 8),
34804 => conv_std_logic_vector(128, 8),
34805 => conv_std_logic_vector(129, 8),
34806 => conv_std_logic_vector(129, 8),
34807 => conv_std_logic_vector(130, 8),
34808 => conv_std_logic_vector(130, 8),
34809 => conv_std_logic_vector(131, 8),
34810 => conv_std_logic_vector(131, 8),
34811 => conv_std_logic_vector(132, 8),
34812 => conv_std_logic_vector(132, 8),
34813 => conv_std_logic_vector(133, 8),
34814 => conv_std_logic_vector(133, 8),
34815 => conv_std_logic_vector(134, 8),
34816 => conv_std_logic_vector(0, 8),
34817 => conv_std_logic_vector(0, 8),
34818 => conv_std_logic_vector(1, 8),
34819 => conv_std_logic_vector(1, 8),
34820 => conv_std_logic_vector(2, 8),
34821 => conv_std_logic_vector(2, 8),
34822 => conv_std_logic_vector(3, 8),
34823 => conv_std_logic_vector(3, 8),
34824 => conv_std_logic_vector(4, 8),
34825 => conv_std_logic_vector(4, 8),
34826 => conv_std_logic_vector(5, 8),
34827 => conv_std_logic_vector(5, 8),
34828 => conv_std_logic_vector(6, 8),
34829 => conv_std_logic_vector(6, 8),
34830 => conv_std_logic_vector(7, 8),
34831 => conv_std_logic_vector(7, 8),
34832 => conv_std_logic_vector(8, 8),
34833 => conv_std_logic_vector(9, 8),
34834 => conv_std_logic_vector(9, 8),
34835 => conv_std_logic_vector(10, 8),
34836 => conv_std_logic_vector(10, 8),
34837 => conv_std_logic_vector(11, 8),
34838 => conv_std_logic_vector(11, 8),
34839 => conv_std_logic_vector(12, 8),
34840 => conv_std_logic_vector(12, 8),
34841 => conv_std_logic_vector(13, 8),
34842 => conv_std_logic_vector(13, 8),
34843 => conv_std_logic_vector(14, 8),
34844 => conv_std_logic_vector(14, 8),
34845 => conv_std_logic_vector(15, 8),
34846 => conv_std_logic_vector(15, 8),
34847 => conv_std_logic_vector(16, 8),
34848 => conv_std_logic_vector(17, 8),
34849 => conv_std_logic_vector(17, 8),
34850 => conv_std_logic_vector(18, 8),
34851 => conv_std_logic_vector(18, 8),
34852 => conv_std_logic_vector(19, 8),
34853 => conv_std_logic_vector(19, 8),
34854 => conv_std_logic_vector(20, 8),
34855 => conv_std_logic_vector(20, 8),
34856 => conv_std_logic_vector(21, 8),
34857 => conv_std_logic_vector(21, 8),
34858 => conv_std_logic_vector(22, 8),
34859 => conv_std_logic_vector(22, 8),
34860 => conv_std_logic_vector(23, 8),
34861 => conv_std_logic_vector(23, 8),
34862 => conv_std_logic_vector(24, 8),
34863 => conv_std_logic_vector(24, 8),
34864 => conv_std_logic_vector(25, 8),
34865 => conv_std_logic_vector(26, 8),
34866 => conv_std_logic_vector(26, 8),
34867 => conv_std_logic_vector(27, 8),
34868 => conv_std_logic_vector(27, 8),
34869 => conv_std_logic_vector(28, 8),
34870 => conv_std_logic_vector(28, 8),
34871 => conv_std_logic_vector(29, 8),
34872 => conv_std_logic_vector(29, 8),
34873 => conv_std_logic_vector(30, 8),
34874 => conv_std_logic_vector(30, 8),
34875 => conv_std_logic_vector(31, 8),
34876 => conv_std_logic_vector(31, 8),
34877 => conv_std_logic_vector(32, 8),
34878 => conv_std_logic_vector(32, 8),
34879 => conv_std_logic_vector(33, 8),
34880 => conv_std_logic_vector(34, 8),
34881 => conv_std_logic_vector(34, 8),
34882 => conv_std_logic_vector(35, 8),
34883 => conv_std_logic_vector(35, 8),
34884 => conv_std_logic_vector(36, 8),
34885 => conv_std_logic_vector(36, 8),
34886 => conv_std_logic_vector(37, 8),
34887 => conv_std_logic_vector(37, 8),
34888 => conv_std_logic_vector(38, 8),
34889 => conv_std_logic_vector(38, 8),
34890 => conv_std_logic_vector(39, 8),
34891 => conv_std_logic_vector(39, 8),
34892 => conv_std_logic_vector(40, 8),
34893 => conv_std_logic_vector(40, 8),
34894 => conv_std_logic_vector(41, 8),
34895 => conv_std_logic_vector(41, 8),
34896 => conv_std_logic_vector(42, 8),
34897 => conv_std_logic_vector(43, 8),
34898 => conv_std_logic_vector(43, 8),
34899 => conv_std_logic_vector(44, 8),
34900 => conv_std_logic_vector(44, 8),
34901 => conv_std_logic_vector(45, 8),
34902 => conv_std_logic_vector(45, 8),
34903 => conv_std_logic_vector(46, 8),
34904 => conv_std_logic_vector(46, 8),
34905 => conv_std_logic_vector(47, 8),
34906 => conv_std_logic_vector(47, 8),
34907 => conv_std_logic_vector(48, 8),
34908 => conv_std_logic_vector(48, 8),
34909 => conv_std_logic_vector(49, 8),
34910 => conv_std_logic_vector(49, 8),
34911 => conv_std_logic_vector(50, 8),
34912 => conv_std_logic_vector(51, 8),
34913 => conv_std_logic_vector(51, 8),
34914 => conv_std_logic_vector(52, 8),
34915 => conv_std_logic_vector(52, 8),
34916 => conv_std_logic_vector(53, 8),
34917 => conv_std_logic_vector(53, 8),
34918 => conv_std_logic_vector(54, 8),
34919 => conv_std_logic_vector(54, 8),
34920 => conv_std_logic_vector(55, 8),
34921 => conv_std_logic_vector(55, 8),
34922 => conv_std_logic_vector(56, 8),
34923 => conv_std_logic_vector(56, 8),
34924 => conv_std_logic_vector(57, 8),
34925 => conv_std_logic_vector(57, 8),
34926 => conv_std_logic_vector(58, 8),
34927 => conv_std_logic_vector(58, 8),
34928 => conv_std_logic_vector(59, 8),
34929 => conv_std_logic_vector(60, 8),
34930 => conv_std_logic_vector(60, 8),
34931 => conv_std_logic_vector(61, 8),
34932 => conv_std_logic_vector(61, 8),
34933 => conv_std_logic_vector(62, 8),
34934 => conv_std_logic_vector(62, 8),
34935 => conv_std_logic_vector(63, 8),
34936 => conv_std_logic_vector(63, 8),
34937 => conv_std_logic_vector(64, 8),
34938 => conv_std_logic_vector(64, 8),
34939 => conv_std_logic_vector(65, 8),
34940 => conv_std_logic_vector(65, 8),
34941 => conv_std_logic_vector(66, 8),
34942 => conv_std_logic_vector(66, 8),
34943 => conv_std_logic_vector(67, 8),
34944 => conv_std_logic_vector(68, 8),
34945 => conv_std_logic_vector(68, 8),
34946 => conv_std_logic_vector(69, 8),
34947 => conv_std_logic_vector(69, 8),
34948 => conv_std_logic_vector(70, 8),
34949 => conv_std_logic_vector(70, 8),
34950 => conv_std_logic_vector(71, 8),
34951 => conv_std_logic_vector(71, 8),
34952 => conv_std_logic_vector(72, 8),
34953 => conv_std_logic_vector(72, 8),
34954 => conv_std_logic_vector(73, 8),
34955 => conv_std_logic_vector(73, 8),
34956 => conv_std_logic_vector(74, 8),
34957 => conv_std_logic_vector(74, 8),
34958 => conv_std_logic_vector(75, 8),
34959 => conv_std_logic_vector(75, 8),
34960 => conv_std_logic_vector(76, 8),
34961 => conv_std_logic_vector(77, 8),
34962 => conv_std_logic_vector(77, 8),
34963 => conv_std_logic_vector(78, 8),
34964 => conv_std_logic_vector(78, 8),
34965 => conv_std_logic_vector(79, 8),
34966 => conv_std_logic_vector(79, 8),
34967 => conv_std_logic_vector(80, 8),
34968 => conv_std_logic_vector(80, 8),
34969 => conv_std_logic_vector(81, 8),
34970 => conv_std_logic_vector(81, 8),
34971 => conv_std_logic_vector(82, 8),
34972 => conv_std_logic_vector(82, 8),
34973 => conv_std_logic_vector(83, 8),
34974 => conv_std_logic_vector(83, 8),
34975 => conv_std_logic_vector(84, 8),
34976 => conv_std_logic_vector(85, 8),
34977 => conv_std_logic_vector(85, 8),
34978 => conv_std_logic_vector(86, 8),
34979 => conv_std_logic_vector(86, 8),
34980 => conv_std_logic_vector(87, 8),
34981 => conv_std_logic_vector(87, 8),
34982 => conv_std_logic_vector(88, 8),
34983 => conv_std_logic_vector(88, 8),
34984 => conv_std_logic_vector(89, 8),
34985 => conv_std_logic_vector(89, 8),
34986 => conv_std_logic_vector(90, 8),
34987 => conv_std_logic_vector(90, 8),
34988 => conv_std_logic_vector(91, 8),
34989 => conv_std_logic_vector(91, 8),
34990 => conv_std_logic_vector(92, 8),
34991 => conv_std_logic_vector(92, 8),
34992 => conv_std_logic_vector(93, 8),
34993 => conv_std_logic_vector(94, 8),
34994 => conv_std_logic_vector(94, 8),
34995 => conv_std_logic_vector(95, 8),
34996 => conv_std_logic_vector(95, 8),
34997 => conv_std_logic_vector(96, 8),
34998 => conv_std_logic_vector(96, 8),
34999 => conv_std_logic_vector(97, 8),
35000 => conv_std_logic_vector(97, 8),
35001 => conv_std_logic_vector(98, 8),
35002 => conv_std_logic_vector(98, 8),
35003 => conv_std_logic_vector(99, 8),
35004 => conv_std_logic_vector(99, 8),
35005 => conv_std_logic_vector(100, 8),
35006 => conv_std_logic_vector(100, 8),
35007 => conv_std_logic_vector(101, 8),
35008 => conv_std_logic_vector(102, 8),
35009 => conv_std_logic_vector(102, 8),
35010 => conv_std_logic_vector(103, 8),
35011 => conv_std_logic_vector(103, 8),
35012 => conv_std_logic_vector(104, 8),
35013 => conv_std_logic_vector(104, 8),
35014 => conv_std_logic_vector(105, 8),
35015 => conv_std_logic_vector(105, 8),
35016 => conv_std_logic_vector(106, 8),
35017 => conv_std_logic_vector(106, 8),
35018 => conv_std_logic_vector(107, 8),
35019 => conv_std_logic_vector(107, 8),
35020 => conv_std_logic_vector(108, 8),
35021 => conv_std_logic_vector(108, 8),
35022 => conv_std_logic_vector(109, 8),
35023 => conv_std_logic_vector(109, 8),
35024 => conv_std_logic_vector(110, 8),
35025 => conv_std_logic_vector(111, 8),
35026 => conv_std_logic_vector(111, 8),
35027 => conv_std_logic_vector(112, 8),
35028 => conv_std_logic_vector(112, 8),
35029 => conv_std_logic_vector(113, 8),
35030 => conv_std_logic_vector(113, 8),
35031 => conv_std_logic_vector(114, 8),
35032 => conv_std_logic_vector(114, 8),
35033 => conv_std_logic_vector(115, 8),
35034 => conv_std_logic_vector(115, 8),
35035 => conv_std_logic_vector(116, 8),
35036 => conv_std_logic_vector(116, 8),
35037 => conv_std_logic_vector(117, 8),
35038 => conv_std_logic_vector(117, 8),
35039 => conv_std_logic_vector(118, 8),
35040 => conv_std_logic_vector(119, 8),
35041 => conv_std_logic_vector(119, 8),
35042 => conv_std_logic_vector(120, 8),
35043 => conv_std_logic_vector(120, 8),
35044 => conv_std_logic_vector(121, 8),
35045 => conv_std_logic_vector(121, 8),
35046 => conv_std_logic_vector(122, 8),
35047 => conv_std_logic_vector(122, 8),
35048 => conv_std_logic_vector(123, 8),
35049 => conv_std_logic_vector(123, 8),
35050 => conv_std_logic_vector(124, 8),
35051 => conv_std_logic_vector(124, 8),
35052 => conv_std_logic_vector(125, 8),
35053 => conv_std_logic_vector(125, 8),
35054 => conv_std_logic_vector(126, 8),
35055 => conv_std_logic_vector(126, 8),
35056 => conv_std_logic_vector(127, 8),
35057 => conv_std_logic_vector(128, 8),
35058 => conv_std_logic_vector(128, 8),
35059 => conv_std_logic_vector(129, 8),
35060 => conv_std_logic_vector(129, 8),
35061 => conv_std_logic_vector(130, 8),
35062 => conv_std_logic_vector(130, 8),
35063 => conv_std_logic_vector(131, 8),
35064 => conv_std_logic_vector(131, 8),
35065 => conv_std_logic_vector(132, 8),
35066 => conv_std_logic_vector(132, 8),
35067 => conv_std_logic_vector(133, 8),
35068 => conv_std_logic_vector(133, 8),
35069 => conv_std_logic_vector(134, 8),
35070 => conv_std_logic_vector(134, 8),
35071 => conv_std_logic_vector(135, 8),
35072 => conv_std_logic_vector(0, 8),
35073 => conv_std_logic_vector(0, 8),
35074 => conv_std_logic_vector(1, 8),
35075 => conv_std_logic_vector(1, 8),
35076 => conv_std_logic_vector(2, 8),
35077 => conv_std_logic_vector(2, 8),
35078 => conv_std_logic_vector(3, 8),
35079 => conv_std_logic_vector(3, 8),
35080 => conv_std_logic_vector(4, 8),
35081 => conv_std_logic_vector(4, 8),
35082 => conv_std_logic_vector(5, 8),
35083 => conv_std_logic_vector(5, 8),
35084 => conv_std_logic_vector(6, 8),
35085 => conv_std_logic_vector(6, 8),
35086 => conv_std_logic_vector(7, 8),
35087 => conv_std_logic_vector(8, 8),
35088 => conv_std_logic_vector(8, 8),
35089 => conv_std_logic_vector(9, 8),
35090 => conv_std_logic_vector(9, 8),
35091 => conv_std_logic_vector(10, 8),
35092 => conv_std_logic_vector(10, 8),
35093 => conv_std_logic_vector(11, 8),
35094 => conv_std_logic_vector(11, 8),
35095 => conv_std_logic_vector(12, 8),
35096 => conv_std_logic_vector(12, 8),
35097 => conv_std_logic_vector(13, 8),
35098 => conv_std_logic_vector(13, 8),
35099 => conv_std_logic_vector(14, 8),
35100 => conv_std_logic_vector(14, 8),
35101 => conv_std_logic_vector(15, 8),
35102 => conv_std_logic_vector(16, 8),
35103 => conv_std_logic_vector(16, 8),
35104 => conv_std_logic_vector(17, 8),
35105 => conv_std_logic_vector(17, 8),
35106 => conv_std_logic_vector(18, 8),
35107 => conv_std_logic_vector(18, 8),
35108 => conv_std_logic_vector(19, 8),
35109 => conv_std_logic_vector(19, 8),
35110 => conv_std_logic_vector(20, 8),
35111 => conv_std_logic_vector(20, 8),
35112 => conv_std_logic_vector(21, 8),
35113 => conv_std_logic_vector(21, 8),
35114 => conv_std_logic_vector(22, 8),
35115 => conv_std_logic_vector(23, 8),
35116 => conv_std_logic_vector(23, 8),
35117 => conv_std_logic_vector(24, 8),
35118 => conv_std_logic_vector(24, 8),
35119 => conv_std_logic_vector(25, 8),
35120 => conv_std_logic_vector(25, 8),
35121 => conv_std_logic_vector(26, 8),
35122 => conv_std_logic_vector(26, 8),
35123 => conv_std_logic_vector(27, 8),
35124 => conv_std_logic_vector(27, 8),
35125 => conv_std_logic_vector(28, 8),
35126 => conv_std_logic_vector(28, 8),
35127 => conv_std_logic_vector(29, 8),
35128 => conv_std_logic_vector(29, 8),
35129 => conv_std_logic_vector(30, 8),
35130 => conv_std_logic_vector(31, 8),
35131 => conv_std_logic_vector(31, 8),
35132 => conv_std_logic_vector(32, 8),
35133 => conv_std_logic_vector(32, 8),
35134 => conv_std_logic_vector(33, 8),
35135 => conv_std_logic_vector(33, 8),
35136 => conv_std_logic_vector(34, 8),
35137 => conv_std_logic_vector(34, 8),
35138 => conv_std_logic_vector(35, 8),
35139 => conv_std_logic_vector(35, 8),
35140 => conv_std_logic_vector(36, 8),
35141 => conv_std_logic_vector(36, 8),
35142 => conv_std_logic_vector(37, 8),
35143 => conv_std_logic_vector(37, 8),
35144 => conv_std_logic_vector(38, 8),
35145 => conv_std_logic_vector(39, 8),
35146 => conv_std_logic_vector(39, 8),
35147 => conv_std_logic_vector(40, 8),
35148 => conv_std_logic_vector(40, 8),
35149 => conv_std_logic_vector(41, 8),
35150 => conv_std_logic_vector(41, 8),
35151 => conv_std_logic_vector(42, 8),
35152 => conv_std_logic_vector(42, 8),
35153 => conv_std_logic_vector(43, 8),
35154 => conv_std_logic_vector(43, 8),
35155 => conv_std_logic_vector(44, 8),
35156 => conv_std_logic_vector(44, 8),
35157 => conv_std_logic_vector(45, 8),
35158 => conv_std_logic_vector(46, 8),
35159 => conv_std_logic_vector(46, 8),
35160 => conv_std_logic_vector(47, 8),
35161 => conv_std_logic_vector(47, 8),
35162 => conv_std_logic_vector(48, 8),
35163 => conv_std_logic_vector(48, 8),
35164 => conv_std_logic_vector(49, 8),
35165 => conv_std_logic_vector(49, 8),
35166 => conv_std_logic_vector(50, 8),
35167 => conv_std_logic_vector(50, 8),
35168 => conv_std_logic_vector(51, 8),
35169 => conv_std_logic_vector(51, 8),
35170 => conv_std_logic_vector(52, 8),
35171 => conv_std_logic_vector(52, 8),
35172 => conv_std_logic_vector(53, 8),
35173 => conv_std_logic_vector(54, 8),
35174 => conv_std_logic_vector(54, 8),
35175 => conv_std_logic_vector(55, 8),
35176 => conv_std_logic_vector(55, 8),
35177 => conv_std_logic_vector(56, 8),
35178 => conv_std_logic_vector(56, 8),
35179 => conv_std_logic_vector(57, 8),
35180 => conv_std_logic_vector(57, 8),
35181 => conv_std_logic_vector(58, 8),
35182 => conv_std_logic_vector(58, 8),
35183 => conv_std_logic_vector(59, 8),
35184 => conv_std_logic_vector(59, 8),
35185 => conv_std_logic_vector(60, 8),
35186 => conv_std_logic_vector(61, 8),
35187 => conv_std_logic_vector(61, 8),
35188 => conv_std_logic_vector(62, 8),
35189 => conv_std_logic_vector(62, 8),
35190 => conv_std_logic_vector(63, 8),
35191 => conv_std_logic_vector(63, 8),
35192 => conv_std_logic_vector(64, 8),
35193 => conv_std_logic_vector(64, 8),
35194 => conv_std_logic_vector(65, 8),
35195 => conv_std_logic_vector(65, 8),
35196 => conv_std_logic_vector(66, 8),
35197 => conv_std_logic_vector(66, 8),
35198 => conv_std_logic_vector(67, 8),
35199 => conv_std_logic_vector(67, 8),
35200 => conv_std_logic_vector(68, 8),
35201 => conv_std_logic_vector(69, 8),
35202 => conv_std_logic_vector(69, 8),
35203 => conv_std_logic_vector(70, 8),
35204 => conv_std_logic_vector(70, 8),
35205 => conv_std_logic_vector(71, 8),
35206 => conv_std_logic_vector(71, 8),
35207 => conv_std_logic_vector(72, 8),
35208 => conv_std_logic_vector(72, 8),
35209 => conv_std_logic_vector(73, 8),
35210 => conv_std_logic_vector(73, 8),
35211 => conv_std_logic_vector(74, 8),
35212 => conv_std_logic_vector(74, 8),
35213 => conv_std_logic_vector(75, 8),
35214 => conv_std_logic_vector(75, 8),
35215 => conv_std_logic_vector(76, 8),
35216 => conv_std_logic_vector(77, 8),
35217 => conv_std_logic_vector(77, 8),
35218 => conv_std_logic_vector(78, 8),
35219 => conv_std_logic_vector(78, 8),
35220 => conv_std_logic_vector(79, 8),
35221 => conv_std_logic_vector(79, 8),
35222 => conv_std_logic_vector(80, 8),
35223 => conv_std_logic_vector(80, 8),
35224 => conv_std_logic_vector(81, 8),
35225 => conv_std_logic_vector(81, 8),
35226 => conv_std_logic_vector(82, 8),
35227 => conv_std_logic_vector(82, 8),
35228 => conv_std_logic_vector(83, 8),
35229 => conv_std_logic_vector(84, 8),
35230 => conv_std_logic_vector(84, 8),
35231 => conv_std_logic_vector(85, 8),
35232 => conv_std_logic_vector(85, 8),
35233 => conv_std_logic_vector(86, 8),
35234 => conv_std_logic_vector(86, 8),
35235 => conv_std_logic_vector(87, 8),
35236 => conv_std_logic_vector(87, 8),
35237 => conv_std_logic_vector(88, 8),
35238 => conv_std_logic_vector(88, 8),
35239 => conv_std_logic_vector(89, 8),
35240 => conv_std_logic_vector(89, 8),
35241 => conv_std_logic_vector(90, 8),
35242 => conv_std_logic_vector(90, 8),
35243 => conv_std_logic_vector(91, 8),
35244 => conv_std_logic_vector(92, 8),
35245 => conv_std_logic_vector(92, 8),
35246 => conv_std_logic_vector(93, 8),
35247 => conv_std_logic_vector(93, 8),
35248 => conv_std_logic_vector(94, 8),
35249 => conv_std_logic_vector(94, 8),
35250 => conv_std_logic_vector(95, 8),
35251 => conv_std_logic_vector(95, 8),
35252 => conv_std_logic_vector(96, 8),
35253 => conv_std_logic_vector(96, 8),
35254 => conv_std_logic_vector(97, 8),
35255 => conv_std_logic_vector(97, 8),
35256 => conv_std_logic_vector(98, 8),
35257 => conv_std_logic_vector(99, 8),
35258 => conv_std_logic_vector(99, 8),
35259 => conv_std_logic_vector(100, 8),
35260 => conv_std_logic_vector(100, 8),
35261 => conv_std_logic_vector(101, 8),
35262 => conv_std_logic_vector(101, 8),
35263 => conv_std_logic_vector(102, 8),
35264 => conv_std_logic_vector(102, 8),
35265 => conv_std_logic_vector(103, 8),
35266 => conv_std_logic_vector(103, 8),
35267 => conv_std_logic_vector(104, 8),
35268 => conv_std_logic_vector(104, 8),
35269 => conv_std_logic_vector(105, 8),
35270 => conv_std_logic_vector(105, 8),
35271 => conv_std_logic_vector(106, 8),
35272 => conv_std_logic_vector(107, 8),
35273 => conv_std_logic_vector(107, 8),
35274 => conv_std_logic_vector(108, 8),
35275 => conv_std_logic_vector(108, 8),
35276 => conv_std_logic_vector(109, 8),
35277 => conv_std_logic_vector(109, 8),
35278 => conv_std_logic_vector(110, 8),
35279 => conv_std_logic_vector(110, 8),
35280 => conv_std_logic_vector(111, 8),
35281 => conv_std_logic_vector(111, 8),
35282 => conv_std_logic_vector(112, 8),
35283 => conv_std_logic_vector(112, 8),
35284 => conv_std_logic_vector(113, 8),
35285 => conv_std_logic_vector(113, 8),
35286 => conv_std_logic_vector(114, 8),
35287 => conv_std_logic_vector(115, 8),
35288 => conv_std_logic_vector(115, 8),
35289 => conv_std_logic_vector(116, 8),
35290 => conv_std_logic_vector(116, 8),
35291 => conv_std_logic_vector(117, 8),
35292 => conv_std_logic_vector(117, 8),
35293 => conv_std_logic_vector(118, 8),
35294 => conv_std_logic_vector(118, 8),
35295 => conv_std_logic_vector(119, 8),
35296 => conv_std_logic_vector(119, 8),
35297 => conv_std_logic_vector(120, 8),
35298 => conv_std_logic_vector(120, 8),
35299 => conv_std_logic_vector(121, 8),
35300 => conv_std_logic_vector(122, 8),
35301 => conv_std_logic_vector(122, 8),
35302 => conv_std_logic_vector(123, 8),
35303 => conv_std_logic_vector(123, 8),
35304 => conv_std_logic_vector(124, 8),
35305 => conv_std_logic_vector(124, 8),
35306 => conv_std_logic_vector(125, 8),
35307 => conv_std_logic_vector(125, 8),
35308 => conv_std_logic_vector(126, 8),
35309 => conv_std_logic_vector(126, 8),
35310 => conv_std_logic_vector(127, 8),
35311 => conv_std_logic_vector(127, 8),
35312 => conv_std_logic_vector(128, 8),
35313 => conv_std_logic_vector(128, 8),
35314 => conv_std_logic_vector(129, 8),
35315 => conv_std_logic_vector(130, 8),
35316 => conv_std_logic_vector(130, 8),
35317 => conv_std_logic_vector(131, 8),
35318 => conv_std_logic_vector(131, 8),
35319 => conv_std_logic_vector(132, 8),
35320 => conv_std_logic_vector(132, 8),
35321 => conv_std_logic_vector(133, 8),
35322 => conv_std_logic_vector(133, 8),
35323 => conv_std_logic_vector(134, 8),
35324 => conv_std_logic_vector(134, 8),
35325 => conv_std_logic_vector(135, 8),
35326 => conv_std_logic_vector(135, 8),
35327 => conv_std_logic_vector(136, 8),
35328 => conv_std_logic_vector(0, 8),
35329 => conv_std_logic_vector(0, 8),
35330 => conv_std_logic_vector(1, 8),
35331 => conv_std_logic_vector(1, 8),
35332 => conv_std_logic_vector(2, 8),
35333 => conv_std_logic_vector(2, 8),
35334 => conv_std_logic_vector(3, 8),
35335 => conv_std_logic_vector(3, 8),
35336 => conv_std_logic_vector(4, 8),
35337 => conv_std_logic_vector(4, 8),
35338 => conv_std_logic_vector(5, 8),
35339 => conv_std_logic_vector(5, 8),
35340 => conv_std_logic_vector(6, 8),
35341 => conv_std_logic_vector(7, 8),
35342 => conv_std_logic_vector(7, 8),
35343 => conv_std_logic_vector(8, 8),
35344 => conv_std_logic_vector(8, 8),
35345 => conv_std_logic_vector(9, 8),
35346 => conv_std_logic_vector(9, 8),
35347 => conv_std_logic_vector(10, 8),
35348 => conv_std_logic_vector(10, 8),
35349 => conv_std_logic_vector(11, 8),
35350 => conv_std_logic_vector(11, 8),
35351 => conv_std_logic_vector(12, 8),
35352 => conv_std_logic_vector(12, 8),
35353 => conv_std_logic_vector(13, 8),
35354 => conv_std_logic_vector(14, 8),
35355 => conv_std_logic_vector(14, 8),
35356 => conv_std_logic_vector(15, 8),
35357 => conv_std_logic_vector(15, 8),
35358 => conv_std_logic_vector(16, 8),
35359 => conv_std_logic_vector(16, 8),
35360 => conv_std_logic_vector(17, 8),
35361 => conv_std_logic_vector(17, 8),
35362 => conv_std_logic_vector(18, 8),
35363 => conv_std_logic_vector(18, 8),
35364 => conv_std_logic_vector(19, 8),
35365 => conv_std_logic_vector(19, 8),
35366 => conv_std_logic_vector(20, 8),
35367 => conv_std_logic_vector(21, 8),
35368 => conv_std_logic_vector(21, 8),
35369 => conv_std_logic_vector(22, 8),
35370 => conv_std_logic_vector(22, 8),
35371 => conv_std_logic_vector(23, 8),
35372 => conv_std_logic_vector(23, 8),
35373 => conv_std_logic_vector(24, 8),
35374 => conv_std_logic_vector(24, 8),
35375 => conv_std_logic_vector(25, 8),
35376 => conv_std_logic_vector(25, 8),
35377 => conv_std_logic_vector(26, 8),
35378 => conv_std_logic_vector(26, 8),
35379 => conv_std_logic_vector(27, 8),
35380 => conv_std_logic_vector(28, 8),
35381 => conv_std_logic_vector(28, 8),
35382 => conv_std_logic_vector(29, 8),
35383 => conv_std_logic_vector(29, 8),
35384 => conv_std_logic_vector(30, 8),
35385 => conv_std_logic_vector(30, 8),
35386 => conv_std_logic_vector(31, 8),
35387 => conv_std_logic_vector(31, 8),
35388 => conv_std_logic_vector(32, 8),
35389 => conv_std_logic_vector(32, 8),
35390 => conv_std_logic_vector(33, 8),
35391 => conv_std_logic_vector(33, 8),
35392 => conv_std_logic_vector(34, 8),
35393 => conv_std_logic_vector(35, 8),
35394 => conv_std_logic_vector(35, 8),
35395 => conv_std_logic_vector(36, 8),
35396 => conv_std_logic_vector(36, 8),
35397 => conv_std_logic_vector(37, 8),
35398 => conv_std_logic_vector(37, 8),
35399 => conv_std_logic_vector(38, 8),
35400 => conv_std_logic_vector(38, 8),
35401 => conv_std_logic_vector(39, 8),
35402 => conv_std_logic_vector(39, 8),
35403 => conv_std_logic_vector(40, 8),
35404 => conv_std_logic_vector(40, 8),
35405 => conv_std_logic_vector(41, 8),
35406 => conv_std_logic_vector(42, 8),
35407 => conv_std_logic_vector(42, 8),
35408 => conv_std_logic_vector(43, 8),
35409 => conv_std_logic_vector(43, 8),
35410 => conv_std_logic_vector(44, 8),
35411 => conv_std_logic_vector(44, 8),
35412 => conv_std_logic_vector(45, 8),
35413 => conv_std_logic_vector(45, 8),
35414 => conv_std_logic_vector(46, 8),
35415 => conv_std_logic_vector(46, 8),
35416 => conv_std_logic_vector(47, 8),
35417 => conv_std_logic_vector(47, 8),
35418 => conv_std_logic_vector(48, 8),
35419 => conv_std_logic_vector(49, 8),
35420 => conv_std_logic_vector(49, 8),
35421 => conv_std_logic_vector(50, 8),
35422 => conv_std_logic_vector(50, 8),
35423 => conv_std_logic_vector(51, 8),
35424 => conv_std_logic_vector(51, 8),
35425 => conv_std_logic_vector(52, 8),
35426 => conv_std_logic_vector(52, 8),
35427 => conv_std_logic_vector(53, 8),
35428 => conv_std_logic_vector(53, 8),
35429 => conv_std_logic_vector(54, 8),
35430 => conv_std_logic_vector(54, 8),
35431 => conv_std_logic_vector(55, 8),
35432 => conv_std_logic_vector(56, 8),
35433 => conv_std_logic_vector(56, 8),
35434 => conv_std_logic_vector(57, 8),
35435 => conv_std_logic_vector(57, 8),
35436 => conv_std_logic_vector(58, 8),
35437 => conv_std_logic_vector(58, 8),
35438 => conv_std_logic_vector(59, 8),
35439 => conv_std_logic_vector(59, 8),
35440 => conv_std_logic_vector(60, 8),
35441 => conv_std_logic_vector(60, 8),
35442 => conv_std_logic_vector(61, 8),
35443 => conv_std_logic_vector(61, 8),
35444 => conv_std_logic_vector(62, 8),
35445 => conv_std_logic_vector(63, 8),
35446 => conv_std_logic_vector(63, 8),
35447 => conv_std_logic_vector(64, 8),
35448 => conv_std_logic_vector(64, 8),
35449 => conv_std_logic_vector(65, 8),
35450 => conv_std_logic_vector(65, 8),
35451 => conv_std_logic_vector(66, 8),
35452 => conv_std_logic_vector(66, 8),
35453 => conv_std_logic_vector(67, 8),
35454 => conv_std_logic_vector(67, 8),
35455 => conv_std_logic_vector(68, 8),
35456 => conv_std_logic_vector(69, 8),
35457 => conv_std_logic_vector(69, 8),
35458 => conv_std_logic_vector(70, 8),
35459 => conv_std_logic_vector(70, 8),
35460 => conv_std_logic_vector(71, 8),
35461 => conv_std_logic_vector(71, 8),
35462 => conv_std_logic_vector(72, 8),
35463 => conv_std_logic_vector(72, 8),
35464 => conv_std_logic_vector(73, 8),
35465 => conv_std_logic_vector(73, 8),
35466 => conv_std_logic_vector(74, 8),
35467 => conv_std_logic_vector(74, 8),
35468 => conv_std_logic_vector(75, 8),
35469 => conv_std_logic_vector(76, 8),
35470 => conv_std_logic_vector(76, 8),
35471 => conv_std_logic_vector(77, 8),
35472 => conv_std_logic_vector(77, 8),
35473 => conv_std_logic_vector(78, 8),
35474 => conv_std_logic_vector(78, 8),
35475 => conv_std_logic_vector(79, 8),
35476 => conv_std_logic_vector(79, 8),
35477 => conv_std_logic_vector(80, 8),
35478 => conv_std_logic_vector(80, 8),
35479 => conv_std_logic_vector(81, 8),
35480 => conv_std_logic_vector(81, 8),
35481 => conv_std_logic_vector(82, 8),
35482 => conv_std_logic_vector(83, 8),
35483 => conv_std_logic_vector(83, 8),
35484 => conv_std_logic_vector(84, 8),
35485 => conv_std_logic_vector(84, 8),
35486 => conv_std_logic_vector(85, 8),
35487 => conv_std_logic_vector(85, 8),
35488 => conv_std_logic_vector(86, 8),
35489 => conv_std_logic_vector(86, 8),
35490 => conv_std_logic_vector(87, 8),
35491 => conv_std_logic_vector(87, 8),
35492 => conv_std_logic_vector(88, 8),
35493 => conv_std_logic_vector(88, 8),
35494 => conv_std_logic_vector(89, 8),
35495 => conv_std_logic_vector(90, 8),
35496 => conv_std_logic_vector(90, 8),
35497 => conv_std_logic_vector(91, 8),
35498 => conv_std_logic_vector(91, 8),
35499 => conv_std_logic_vector(92, 8),
35500 => conv_std_logic_vector(92, 8),
35501 => conv_std_logic_vector(93, 8),
35502 => conv_std_logic_vector(93, 8),
35503 => conv_std_logic_vector(94, 8),
35504 => conv_std_logic_vector(94, 8),
35505 => conv_std_logic_vector(95, 8),
35506 => conv_std_logic_vector(95, 8),
35507 => conv_std_logic_vector(96, 8),
35508 => conv_std_logic_vector(97, 8),
35509 => conv_std_logic_vector(97, 8),
35510 => conv_std_logic_vector(98, 8),
35511 => conv_std_logic_vector(98, 8),
35512 => conv_std_logic_vector(99, 8),
35513 => conv_std_logic_vector(99, 8),
35514 => conv_std_logic_vector(100, 8),
35515 => conv_std_logic_vector(100, 8),
35516 => conv_std_logic_vector(101, 8),
35517 => conv_std_logic_vector(101, 8),
35518 => conv_std_logic_vector(102, 8),
35519 => conv_std_logic_vector(102, 8),
35520 => conv_std_logic_vector(103, 8),
35521 => conv_std_logic_vector(104, 8),
35522 => conv_std_logic_vector(104, 8),
35523 => conv_std_logic_vector(105, 8),
35524 => conv_std_logic_vector(105, 8),
35525 => conv_std_logic_vector(106, 8),
35526 => conv_std_logic_vector(106, 8),
35527 => conv_std_logic_vector(107, 8),
35528 => conv_std_logic_vector(107, 8),
35529 => conv_std_logic_vector(108, 8),
35530 => conv_std_logic_vector(108, 8),
35531 => conv_std_logic_vector(109, 8),
35532 => conv_std_logic_vector(109, 8),
35533 => conv_std_logic_vector(110, 8),
35534 => conv_std_logic_vector(111, 8),
35535 => conv_std_logic_vector(111, 8),
35536 => conv_std_logic_vector(112, 8),
35537 => conv_std_logic_vector(112, 8),
35538 => conv_std_logic_vector(113, 8),
35539 => conv_std_logic_vector(113, 8),
35540 => conv_std_logic_vector(114, 8),
35541 => conv_std_logic_vector(114, 8),
35542 => conv_std_logic_vector(115, 8),
35543 => conv_std_logic_vector(115, 8),
35544 => conv_std_logic_vector(116, 8),
35545 => conv_std_logic_vector(116, 8),
35546 => conv_std_logic_vector(117, 8),
35547 => conv_std_logic_vector(118, 8),
35548 => conv_std_logic_vector(118, 8),
35549 => conv_std_logic_vector(119, 8),
35550 => conv_std_logic_vector(119, 8),
35551 => conv_std_logic_vector(120, 8),
35552 => conv_std_logic_vector(120, 8),
35553 => conv_std_logic_vector(121, 8),
35554 => conv_std_logic_vector(121, 8),
35555 => conv_std_logic_vector(122, 8),
35556 => conv_std_logic_vector(122, 8),
35557 => conv_std_logic_vector(123, 8),
35558 => conv_std_logic_vector(123, 8),
35559 => conv_std_logic_vector(124, 8),
35560 => conv_std_logic_vector(125, 8),
35561 => conv_std_logic_vector(125, 8),
35562 => conv_std_logic_vector(126, 8),
35563 => conv_std_logic_vector(126, 8),
35564 => conv_std_logic_vector(127, 8),
35565 => conv_std_logic_vector(127, 8),
35566 => conv_std_logic_vector(128, 8),
35567 => conv_std_logic_vector(128, 8),
35568 => conv_std_logic_vector(129, 8),
35569 => conv_std_logic_vector(129, 8),
35570 => conv_std_logic_vector(130, 8),
35571 => conv_std_logic_vector(130, 8),
35572 => conv_std_logic_vector(131, 8),
35573 => conv_std_logic_vector(132, 8),
35574 => conv_std_logic_vector(132, 8),
35575 => conv_std_logic_vector(133, 8),
35576 => conv_std_logic_vector(133, 8),
35577 => conv_std_logic_vector(134, 8),
35578 => conv_std_logic_vector(134, 8),
35579 => conv_std_logic_vector(135, 8),
35580 => conv_std_logic_vector(135, 8),
35581 => conv_std_logic_vector(136, 8),
35582 => conv_std_logic_vector(136, 8),
35583 => conv_std_logic_vector(137, 8),
35584 => conv_std_logic_vector(0, 8),
35585 => conv_std_logic_vector(0, 8),
35586 => conv_std_logic_vector(1, 8),
35587 => conv_std_logic_vector(1, 8),
35588 => conv_std_logic_vector(2, 8),
35589 => conv_std_logic_vector(2, 8),
35590 => conv_std_logic_vector(3, 8),
35591 => conv_std_logic_vector(3, 8),
35592 => conv_std_logic_vector(4, 8),
35593 => conv_std_logic_vector(4, 8),
35594 => conv_std_logic_vector(5, 8),
35595 => conv_std_logic_vector(5, 8),
35596 => conv_std_logic_vector(6, 8),
35597 => conv_std_logic_vector(7, 8),
35598 => conv_std_logic_vector(7, 8),
35599 => conv_std_logic_vector(8, 8),
35600 => conv_std_logic_vector(8, 8),
35601 => conv_std_logic_vector(9, 8),
35602 => conv_std_logic_vector(9, 8),
35603 => conv_std_logic_vector(10, 8),
35604 => conv_std_logic_vector(10, 8),
35605 => conv_std_logic_vector(11, 8),
35606 => conv_std_logic_vector(11, 8),
35607 => conv_std_logic_vector(12, 8),
35608 => conv_std_logic_vector(13, 8),
35609 => conv_std_logic_vector(13, 8),
35610 => conv_std_logic_vector(14, 8),
35611 => conv_std_logic_vector(14, 8),
35612 => conv_std_logic_vector(15, 8),
35613 => conv_std_logic_vector(15, 8),
35614 => conv_std_logic_vector(16, 8),
35615 => conv_std_logic_vector(16, 8),
35616 => conv_std_logic_vector(17, 8),
35617 => conv_std_logic_vector(17, 8),
35618 => conv_std_logic_vector(18, 8),
35619 => conv_std_logic_vector(19, 8),
35620 => conv_std_logic_vector(19, 8),
35621 => conv_std_logic_vector(20, 8),
35622 => conv_std_logic_vector(20, 8),
35623 => conv_std_logic_vector(21, 8),
35624 => conv_std_logic_vector(21, 8),
35625 => conv_std_logic_vector(22, 8),
35626 => conv_std_logic_vector(22, 8),
35627 => conv_std_logic_vector(23, 8),
35628 => conv_std_logic_vector(23, 8),
35629 => conv_std_logic_vector(24, 8),
35630 => conv_std_logic_vector(24, 8),
35631 => conv_std_logic_vector(25, 8),
35632 => conv_std_logic_vector(26, 8),
35633 => conv_std_logic_vector(26, 8),
35634 => conv_std_logic_vector(27, 8),
35635 => conv_std_logic_vector(27, 8),
35636 => conv_std_logic_vector(28, 8),
35637 => conv_std_logic_vector(28, 8),
35638 => conv_std_logic_vector(29, 8),
35639 => conv_std_logic_vector(29, 8),
35640 => conv_std_logic_vector(30, 8),
35641 => conv_std_logic_vector(30, 8),
35642 => conv_std_logic_vector(31, 8),
35643 => conv_std_logic_vector(32, 8),
35644 => conv_std_logic_vector(32, 8),
35645 => conv_std_logic_vector(33, 8),
35646 => conv_std_logic_vector(33, 8),
35647 => conv_std_logic_vector(34, 8),
35648 => conv_std_logic_vector(34, 8),
35649 => conv_std_logic_vector(35, 8),
35650 => conv_std_logic_vector(35, 8),
35651 => conv_std_logic_vector(36, 8),
35652 => conv_std_logic_vector(36, 8),
35653 => conv_std_logic_vector(37, 8),
35654 => conv_std_logic_vector(38, 8),
35655 => conv_std_logic_vector(38, 8),
35656 => conv_std_logic_vector(39, 8),
35657 => conv_std_logic_vector(39, 8),
35658 => conv_std_logic_vector(40, 8),
35659 => conv_std_logic_vector(40, 8),
35660 => conv_std_logic_vector(41, 8),
35661 => conv_std_logic_vector(41, 8),
35662 => conv_std_logic_vector(42, 8),
35663 => conv_std_logic_vector(42, 8),
35664 => conv_std_logic_vector(43, 8),
35665 => conv_std_logic_vector(43, 8),
35666 => conv_std_logic_vector(44, 8),
35667 => conv_std_logic_vector(45, 8),
35668 => conv_std_logic_vector(45, 8),
35669 => conv_std_logic_vector(46, 8),
35670 => conv_std_logic_vector(46, 8),
35671 => conv_std_logic_vector(47, 8),
35672 => conv_std_logic_vector(47, 8),
35673 => conv_std_logic_vector(48, 8),
35674 => conv_std_logic_vector(48, 8),
35675 => conv_std_logic_vector(49, 8),
35676 => conv_std_logic_vector(49, 8),
35677 => conv_std_logic_vector(50, 8),
35678 => conv_std_logic_vector(51, 8),
35679 => conv_std_logic_vector(51, 8),
35680 => conv_std_logic_vector(52, 8),
35681 => conv_std_logic_vector(52, 8),
35682 => conv_std_logic_vector(53, 8),
35683 => conv_std_logic_vector(53, 8),
35684 => conv_std_logic_vector(54, 8),
35685 => conv_std_logic_vector(54, 8),
35686 => conv_std_logic_vector(55, 8),
35687 => conv_std_logic_vector(55, 8),
35688 => conv_std_logic_vector(56, 8),
35689 => conv_std_logic_vector(57, 8),
35690 => conv_std_logic_vector(57, 8),
35691 => conv_std_logic_vector(58, 8),
35692 => conv_std_logic_vector(58, 8),
35693 => conv_std_logic_vector(59, 8),
35694 => conv_std_logic_vector(59, 8),
35695 => conv_std_logic_vector(60, 8),
35696 => conv_std_logic_vector(60, 8),
35697 => conv_std_logic_vector(61, 8),
35698 => conv_std_logic_vector(61, 8),
35699 => conv_std_logic_vector(62, 8),
35700 => conv_std_logic_vector(62, 8),
35701 => conv_std_logic_vector(63, 8),
35702 => conv_std_logic_vector(64, 8),
35703 => conv_std_logic_vector(64, 8),
35704 => conv_std_logic_vector(65, 8),
35705 => conv_std_logic_vector(65, 8),
35706 => conv_std_logic_vector(66, 8),
35707 => conv_std_logic_vector(66, 8),
35708 => conv_std_logic_vector(67, 8),
35709 => conv_std_logic_vector(67, 8),
35710 => conv_std_logic_vector(68, 8),
35711 => conv_std_logic_vector(68, 8),
35712 => conv_std_logic_vector(69, 8),
35713 => conv_std_logic_vector(70, 8),
35714 => conv_std_logic_vector(70, 8),
35715 => conv_std_logic_vector(71, 8),
35716 => conv_std_logic_vector(71, 8),
35717 => conv_std_logic_vector(72, 8),
35718 => conv_std_logic_vector(72, 8),
35719 => conv_std_logic_vector(73, 8),
35720 => conv_std_logic_vector(73, 8),
35721 => conv_std_logic_vector(74, 8),
35722 => conv_std_logic_vector(74, 8),
35723 => conv_std_logic_vector(75, 8),
35724 => conv_std_logic_vector(76, 8),
35725 => conv_std_logic_vector(76, 8),
35726 => conv_std_logic_vector(77, 8),
35727 => conv_std_logic_vector(77, 8),
35728 => conv_std_logic_vector(78, 8),
35729 => conv_std_logic_vector(78, 8),
35730 => conv_std_logic_vector(79, 8),
35731 => conv_std_logic_vector(79, 8),
35732 => conv_std_logic_vector(80, 8),
35733 => conv_std_logic_vector(80, 8),
35734 => conv_std_logic_vector(81, 8),
35735 => conv_std_logic_vector(81, 8),
35736 => conv_std_logic_vector(82, 8),
35737 => conv_std_logic_vector(83, 8),
35738 => conv_std_logic_vector(83, 8),
35739 => conv_std_logic_vector(84, 8),
35740 => conv_std_logic_vector(84, 8),
35741 => conv_std_logic_vector(85, 8),
35742 => conv_std_logic_vector(85, 8),
35743 => conv_std_logic_vector(86, 8),
35744 => conv_std_logic_vector(86, 8),
35745 => conv_std_logic_vector(87, 8),
35746 => conv_std_logic_vector(87, 8),
35747 => conv_std_logic_vector(88, 8),
35748 => conv_std_logic_vector(89, 8),
35749 => conv_std_logic_vector(89, 8),
35750 => conv_std_logic_vector(90, 8),
35751 => conv_std_logic_vector(90, 8),
35752 => conv_std_logic_vector(91, 8),
35753 => conv_std_logic_vector(91, 8),
35754 => conv_std_logic_vector(92, 8),
35755 => conv_std_logic_vector(92, 8),
35756 => conv_std_logic_vector(93, 8),
35757 => conv_std_logic_vector(93, 8),
35758 => conv_std_logic_vector(94, 8),
35759 => conv_std_logic_vector(95, 8),
35760 => conv_std_logic_vector(95, 8),
35761 => conv_std_logic_vector(96, 8),
35762 => conv_std_logic_vector(96, 8),
35763 => conv_std_logic_vector(97, 8),
35764 => conv_std_logic_vector(97, 8),
35765 => conv_std_logic_vector(98, 8),
35766 => conv_std_logic_vector(98, 8),
35767 => conv_std_logic_vector(99, 8),
35768 => conv_std_logic_vector(99, 8),
35769 => conv_std_logic_vector(100, 8),
35770 => conv_std_logic_vector(100, 8),
35771 => conv_std_logic_vector(101, 8),
35772 => conv_std_logic_vector(102, 8),
35773 => conv_std_logic_vector(102, 8),
35774 => conv_std_logic_vector(103, 8),
35775 => conv_std_logic_vector(103, 8),
35776 => conv_std_logic_vector(104, 8),
35777 => conv_std_logic_vector(104, 8),
35778 => conv_std_logic_vector(105, 8),
35779 => conv_std_logic_vector(105, 8),
35780 => conv_std_logic_vector(106, 8),
35781 => conv_std_logic_vector(106, 8),
35782 => conv_std_logic_vector(107, 8),
35783 => conv_std_logic_vector(108, 8),
35784 => conv_std_logic_vector(108, 8),
35785 => conv_std_logic_vector(109, 8),
35786 => conv_std_logic_vector(109, 8),
35787 => conv_std_logic_vector(110, 8),
35788 => conv_std_logic_vector(110, 8),
35789 => conv_std_logic_vector(111, 8),
35790 => conv_std_logic_vector(111, 8),
35791 => conv_std_logic_vector(112, 8),
35792 => conv_std_logic_vector(112, 8),
35793 => conv_std_logic_vector(113, 8),
35794 => conv_std_logic_vector(114, 8),
35795 => conv_std_logic_vector(114, 8),
35796 => conv_std_logic_vector(115, 8),
35797 => conv_std_logic_vector(115, 8),
35798 => conv_std_logic_vector(116, 8),
35799 => conv_std_logic_vector(116, 8),
35800 => conv_std_logic_vector(117, 8),
35801 => conv_std_logic_vector(117, 8),
35802 => conv_std_logic_vector(118, 8),
35803 => conv_std_logic_vector(118, 8),
35804 => conv_std_logic_vector(119, 8),
35805 => conv_std_logic_vector(119, 8),
35806 => conv_std_logic_vector(120, 8),
35807 => conv_std_logic_vector(121, 8),
35808 => conv_std_logic_vector(121, 8),
35809 => conv_std_logic_vector(122, 8),
35810 => conv_std_logic_vector(122, 8),
35811 => conv_std_logic_vector(123, 8),
35812 => conv_std_logic_vector(123, 8),
35813 => conv_std_logic_vector(124, 8),
35814 => conv_std_logic_vector(124, 8),
35815 => conv_std_logic_vector(125, 8),
35816 => conv_std_logic_vector(125, 8),
35817 => conv_std_logic_vector(126, 8),
35818 => conv_std_logic_vector(127, 8),
35819 => conv_std_logic_vector(127, 8),
35820 => conv_std_logic_vector(128, 8),
35821 => conv_std_logic_vector(128, 8),
35822 => conv_std_logic_vector(129, 8),
35823 => conv_std_logic_vector(129, 8),
35824 => conv_std_logic_vector(130, 8),
35825 => conv_std_logic_vector(130, 8),
35826 => conv_std_logic_vector(131, 8),
35827 => conv_std_logic_vector(131, 8),
35828 => conv_std_logic_vector(132, 8),
35829 => conv_std_logic_vector(133, 8),
35830 => conv_std_logic_vector(133, 8),
35831 => conv_std_logic_vector(134, 8),
35832 => conv_std_logic_vector(134, 8),
35833 => conv_std_logic_vector(135, 8),
35834 => conv_std_logic_vector(135, 8),
35835 => conv_std_logic_vector(136, 8),
35836 => conv_std_logic_vector(136, 8),
35837 => conv_std_logic_vector(137, 8),
35838 => conv_std_logic_vector(137, 8),
35839 => conv_std_logic_vector(138, 8),
35840 => conv_std_logic_vector(0, 8),
35841 => conv_std_logic_vector(0, 8),
35842 => conv_std_logic_vector(1, 8),
35843 => conv_std_logic_vector(1, 8),
35844 => conv_std_logic_vector(2, 8),
35845 => conv_std_logic_vector(2, 8),
35846 => conv_std_logic_vector(3, 8),
35847 => conv_std_logic_vector(3, 8),
35848 => conv_std_logic_vector(4, 8),
35849 => conv_std_logic_vector(4, 8),
35850 => conv_std_logic_vector(5, 8),
35851 => conv_std_logic_vector(6, 8),
35852 => conv_std_logic_vector(6, 8),
35853 => conv_std_logic_vector(7, 8),
35854 => conv_std_logic_vector(7, 8),
35855 => conv_std_logic_vector(8, 8),
35856 => conv_std_logic_vector(8, 8),
35857 => conv_std_logic_vector(9, 8),
35858 => conv_std_logic_vector(9, 8),
35859 => conv_std_logic_vector(10, 8),
35860 => conv_std_logic_vector(10, 8),
35861 => conv_std_logic_vector(11, 8),
35862 => conv_std_logic_vector(12, 8),
35863 => conv_std_logic_vector(12, 8),
35864 => conv_std_logic_vector(13, 8),
35865 => conv_std_logic_vector(13, 8),
35866 => conv_std_logic_vector(14, 8),
35867 => conv_std_logic_vector(14, 8),
35868 => conv_std_logic_vector(15, 8),
35869 => conv_std_logic_vector(15, 8),
35870 => conv_std_logic_vector(16, 8),
35871 => conv_std_logic_vector(16, 8),
35872 => conv_std_logic_vector(17, 8),
35873 => conv_std_logic_vector(18, 8),
35874 => conv_std_logic_vector(18, 8),
35875 => conv_std_logic_vector(19, 8),
35876 => conv_std_logic_vector(19, 8),
35877 => conv_std_logic_vector(20, 8),
35878 => conv_std_logic_vector(20, 8),
35879 => conv_std_logic_vector(21, 8),
35880 => conv_std_logic_vector(21, 8),
35881 => conv_std_logic_vector(22, 8),
35882 => conv_std_logic_vector(22, 8),
35883 => conv_std_logic_vector(23, 8),
35884 => conv_std_logic_vector(24, 8),
35885 => conv_std_logic_vector(24, 8),
35886 => conv_std_logic_vector(25, 8),
35887 => conv_std_logic_vector(25, 8),
35888 => conv_std_logic_vector(26, 8),
35889 => conv_std_logic_vector(26, 8),
35890 => conv_std_logic_vector(27, 8),
35891 => conv_std_logic_vector(27, 8),
35892 => conv_std_logic_vector(28, 8),
35893 => conv_std_logic_vector(28, 8),
35894 => conv_std_logic_vector(29, 8),
35895 => conv_std_logic_vector(30, 8),
35896 => conv_std_logic_vector(30, 8),
35897 => conv_std_logic_vector(31, 8),
35898 => conv_std_logic_vector(31, 8),
35899 => conv_std_logic_vector(32, 8),
35900 => conv_std_logic_vector(32, 8),
35901 => conv_std_logic_vector(33, 8),
35902 => conv_std_logic_vector(33, 8),
35903 => conv_std_logic_vector(34, 8),
35904 => conv_std_logic_vector(35, 8),
35905 => conv_std_logic_vector(35, 8),
35906 => conv_std_logic_vector(36, 8),
35907 => conv_std_logic_vector(36, 8),
35908 => conv_std_logic_vector(37, 8),
35909 => conv_std_logic_vector(37, 8),
35910 => conv_std_logic_vector(38, 8),
35911 => conv_std_logic_vector(38, 8),
35912 => conv_std_logic_vector(39, 8),
35913 => conv_std_logic_vector(39, 8),
35914 => conv_std_logic_vector(40, 8),
35915 => conv_std_logic_vector(41, 8),
35916 => conv_std_logic_vector(41, 8),
35917 => conv_std_logic_vector(42, 8),
35918 => conv_std_logic_vector(42, 8),
35919 => conv_std_logic_vector(43, 8),
35920 => conv_std_logic_vector(43, 8),
35921 => conv_std_logic_vector(44, 8),
35922 => conv_std_logic_vector(44, 8),
35923 => conv_std_logic_vector(45, 8),
35924 => conv_std_logic_vector(45, 8),
35925 => conv_std_logic_vector(46, 8),
35926 => conv_std_logic_vector(47, 8),
35927 => conv_std_logic_vector(47, 8),
35928 => conv_std_logic_vector(48, 8),
35929 => conv_std_logic_vector(48, 8),
35930 => conv_std_logic_vector(49, 8),
35931 => conv_std_logic_vector(49, 8),
35932 => conv_std_logic_vector(50, 8),
35933 => conv_std_logic_vector(50, 8),
35934 => conv_std_logic_vector(51, 8),
35935 => conv_std_logic_vector(51, 8),
35936 => conv_std_logic_vector(52, 8),
35937 => conv_std_logic_vector(53, 8),
35938 => conv_std_logic_vector(53, 8),
35939 => conv_std_logic_vector(54, 8),
35940 => conv_std_logic_vector(54, 8),
35941 => conv_std_logic_vector(55, 8),
35942 => conv_std_logic_vector(55, 8),
35943 => conv_std_logic_vector(56, 8),
35944 => conv_std_logic_vector(56, 8),
35945 => conv_std_logic_vector(57, 8),
35946 => conv_std_logic_vector(57, 8),
35947 => conv_std_logic_vector(58, 8),
35948 => conv_std_logic_vector(59, 8),
35949 => conv_std_logic_vector(59, 8),
35950 => conv_std_logic_vector(60, 8),
35951 => conv_std_logic_vector(60, 8),
35952 => conv_std_logic_vector(61, 8),
35953 => conv_std_logic_vector(61, 8),
35954 => conv_std_logic_vector(62, 8),
35955 => conv_std_logic_vector(62, 8),
35956 => conv_std_logic_vector(63, 8),
35957 => conv_std_logic_vector(63, 8),
35958 => conv_std_logic_vector(64, 8),
35959 => conv_std_logic_vector(65, 8),
35960 => conv_std_logic_vector(65, 8),
35961 => conv_std_logic_vector(66, 8),
35962 => conv_std_logic_vector(66, 8),
35963 => conv_std_logic_vector(67, 8),
35964 => conv_std_logic_vector(67, 8),
35965 => conv_std_logic_vector(68, 8),
35966 => conv_std_logic_vector(68, 8),
35967 => conv_std_logic_vector(69, 8),
35968 => conv_std_logic_vector(70, 8),
35969 => conv_std_logic_vector(70, 8),
35970 => conv_std_logic_vector(71, 8),
35971 => conv_std_logic_vector(71, 8),
35972 => conv_std_logic_vector(72, 8),
35973 => conv_std_logic_vector(72, 8),
35974 => conv_std_logic_vector(73, 8),
35975 => conv_std_logic_vector(73, 8),
35976 => conv_std_logic_vector(74, 8),
35977 => conv_std_logic_vector(74, 8),
35978 => conv_std_logic_vector(75, 8),
35979 => conv_std_logic_vector(76, 8),
35980 => conv_std_logic_vector(76, 8),
35981 => conv_std_logic_vector(77, 8),
35982 => conv_std_logic_vector(77, 8),
35983 => conv_std_logic_vector(78, 8),
35984 => conv_std_logic_vector(78, 8),
35985 => conv_std_logic_vector(79, 8),
35986 => conv_std_logic_vector(79, 8),
35987 => conv_std_logic_vector(80, 8),
35988 => conv_std_logic_vector(80, 8),
35989 => conv_std_logic_vector(81, 8),
35990 => conv_std_logic_vector(82, 8),
35991 => conv_std_logic_vector(82, 8),
35992 => conv_std_logic_vector(83, 8),
35993 => conv_std_logic_vector(83, 8),
35994 => conv_std_logic_vector(84, 8),
35995 => conv_std_logic_vector(84, 8),
35996 => conv_std_logic_vector(85, 8),
35997 => conv_std_logic_vector(85, 8),
35998 => conv_std_logic_vector(86, 8),
35999 => conv_std_logic_vector(86, 8),
36000 => conv_std_logic_vector(87, 8),
36001 => conv_std_logic_vector(88, 8),
36002 => conv_std_logic_vector(88, 8),
36003 => conv_std_logic_vector(89, 8),
36004 => conv_std_logic_vector(89, 8),
36005 => conv_std_logic_vector(90, 8),
36006 => conv_std_logic_vector(90, 8),
36007 => conv_std_logic_vector(91, 8),
36008 => conv_std_logic_vector(91, 8),
36009 => conv_std_logic_vector(92, 8),
36010 => conv_std_logic_vector(92, 8),
36011 => conv_std_logic_vector(93, 8),
36012 => conv_std_logic_vector(94, 8),
36013 => conv_std_logic_vector(94, 8),
36014 => conv_std_logic_vector(95, 8),
36015 => conv_std_logic_vector(95, 8),
36016 => conv_std_logic_vector(96, 8),
36017 => conv_std_logic_vector(96, 8),
36018 => conv_std_logic_vector(97, 8),
36019 => conv_std_logic_vector(97, 8),
36020 => conv_std_logic_vector(98, 8),
36021 => conv_std_logic_vector(98, 8),
36022 => conv_std_logic_vector(99, 8),
36023 => conv_std_logic_vector(100, 8),
36024 => conv_std_logic_vector(100, 8),
36025 => conv_std_logic_vector(101, 8),
36026 => conv_std_logic_vector(101, 8),
36027 => conv_std_logic_vector(102, 8),
36028 => conv_std_logic_vector(102, 8),
36029 => conv_std_logic_vector(103, 8),
36030 => conv_std_logic_vector(103, 8),
36031 => conv_std_logic_vector(104, 8),
36032 => conv_std_logic_vector(105, 8),
36033 => conv_std_logic_vector(105, 8),
36034 => conv_std_logic_vector(106, 8),
36035 => conv_std_logic_vector(106, 8),
36036 => conv_std_logic_vector(107, 8),
36037 => conv_std_logic_vector(107, 8),
36038 => conv_std_logic_vector(108, 8),
36039 => conv_std_logic_vector(108, 8),
36040 => conv_std_logic_vector(109, 8),
36041 => conv_std_logic_vector(109, 8),
36042 => conv_std_logic_vector(110, 8),
36043 => conv_std_logic_vector(111, 8),
36044 => conv_std_logic_vector(111, 8),
36045 => conv_std_logic_vector(112, 8),
36046 => conv_std_logic_vector(112, 8),
36047 => conv_std_logic_vector(113, 8),
36048 => conv_std_logic_vector(113, 8),
36049 => conv_std_logic_vector(114, 8),
36050 => conv_std_logic_vector(114, 8),
36051 => conv_std_logic_vector(115, 8),
36052 => conv_std_logic_vector(115, 8),
36053 => conv_std_logic_vector(116, 8),
36054 => conv_std_logic_vector(117, 8),
36055 => conv_std_logic_vector(117, 8),
36056 => conv_std_logic_vector(118, 8),
36057 => conv_std_logic_vector(118, 8),
36058 => conv_std_logic_vector(119, 8),
36059 => conv_std_logic_vector(119, 8),
36060 => conv_std_logic_vector(120, 8),
36061 => conv_std_logic_vector(120, 8),
36062 => conv_std_logic_vector(121, 8),
36063 => conv_std_logic_vector(121, 8),
36064 => conv_std_logic_vector(122, 8),
36065 => conv_std_logic_vector(123, 8),
36066 => conv_std_logic_vector(123, 8),
36067 => conv_std_logic_vector(124, 8),
36068 => conv_std_logic_vector(124, 8),
36069 => conv_std_logic_vector(125, 8),
36070 => conv_std_logic_vector(125, 8),
36071 => conv_std_logic_vector(126, 8),
36072 => conv_std_logic_vector(126, 8),
36073 => conv_std_logic_vector(127, 8),
36074 => conv_std_logic_vector(127, 8),
36075 => conv_std_logic_vector(128, 8),
36076 => conv_std_logic_vector(129, 8),
36077 => conv_std_logic_vector(129, 8),
36078 => conv_std_logic_vector(130, 8),
36079 => conv_std_logic_vector(130, 8),
36080 => conv_std_logic_vector(131, 8),
36081 => conv_std_logic_vector(131, 8),
36082 => conv_std_logic_vector(132, 8),
36083 => conv_std_logic_vector(132, 8),
36084 => conv_std_logic_vector(133, 8),
36085 => conv_std_logic_vector(133, 8),
36086 => conv_std_logic_vector(134, 8),
36087 => conv_std_logic_vector(135, 8),
36088 => conv_std_logic_vector(135, 8),
36089 => conv_std_logic_vector(136, 8),
36090 => conv_std_logic_vector(136, 8),
36091 => conv_std_logic_vector(137, 8),
36092 => conv_std_logic_vector(137, 8),
36093 => conv_std_logic_vector(138, 8),
36094 => conv_std_logic_vector(138, 8),
36095 => conv_std_logic_vector(139, 8),
36096 => conv_std_logic_vector(0, 8),
36097 => conv_std_logic_vector(0, 8),
36098 => conv_std_logic_vector(1, 8),
36099 => conv_std_logic_vector(1, 8),
36100 => conv_std_logic_vector(2, 8),
36101 => conv_std_logic_vector(2, 8),
36102 => conv_std_logic_vector(3, 8),
36103 => conv_std_logic_vector(3, 8),
36104 => conv_std_logic_vector(4, 8),
36105 => conv_std_logic_vector(4, 8),
36106 => conv_std_logic_vector(5, 8),
36107 => conv_std_logic_vector(6, 8),
36108 => conv_std_logic_vector(6, 8),
36109 => conv_std_logic_vector(7, 8),
36110 => conv_std_logic_vector(7, 8),
36111 => conv_std_logic_vector(8, 8),
36112 => conv_std_logic_vector(8, 8),
36113 => conv_std_logic_vector(9, 8),
36114 => conv_std_logic_vector(9, 8),
36115 => conv_std_logic_vector(10, 8),
36116 => conv_std_logic_vector(11, 8),
36117 => conv_std_logic_vector(11, 8),
36118 => conv_std_logic_vector(12, 8),
36119 => conv_std_logic_vector(12, 8),
36120 => conv_std_logic_vector(13, 8),
36121 => conv_std_logic_vector(13, 8),
36122 => conv_std_logic_vector(14, 8),
36123 => conv_std_logic_vector(14, 8),
36124 => conv_std_logic_vector(15, 8),
36125 => conv_std_logic_vector(15, 8),
36126 => conv_std_logic_vector(16, 8),
36127 => conv_std_logic_vector(17, 8),
36128 => conv_std_logic_vector(17, 8),
36129 => conv_std_logic_vector(18, 8),
36130 => conv_std_logic_vector(18, 8),
36131 => conv_std_logic_vector(19, 8),
36132 => conv_std_logic_vector(19, 8),
36133 => conv_std_logic_vector(20, 8),
36134 => conv_std_logic_vector(20, 8),
36135 => conv_std_logic_vector(21, 8),
36136 => conv_std_logic_vector(22, 8),
36137 => conv_std_logic_vector(22, 8),
36138 => conv_std_logic_vector(23, 8),
36139 => conv_std_logic_vector(23, 8),
36140 => conv_std_logic_vector(24, 8),
36141 => conv_std_logic_vector(24, 8),
36142 => conv_std_logic_vector(25, 8),
36143 => conv_std_logic_vector(25, 8),
36144 => conv_std_logic_vector(26, 8),
36145 => conv_std_logic_vector(26, 8),
36146 => conv_std_logic_vector(27, 8),
36147 => conv_std_logic_vector(28, 8),
36148 => conv_std_logic_vector(28, 8),
36149 => conv_std_logic_vector(29, 8),
36150 => conv_std_logic_vector(29, 8),
36151 => conv_std_logic_vector(30, 8),
36152 => conv_std_logic_vector(30, 8),
36153 => conv_std_logic_vector(31, 8),
36154 => conv_std_logic_vector(31, 8),
36155 => conv_std_logic_vector(32, 8),
36156 => conv_std_logic_vector(33, 8),
36157 => conv_std_logic_vector(33, 8),
36158 => conv_std_logic_vector(34, 8),
36159 => conv_std_logic_vector(34, 8),
36160 => conv_std_logic_vector(35, 8),
36161 => conv_std_logic_vector(35, 8),
36162 => conv_std_logic_vector(36, 8),
36163 => conv_std_logic_vector(36, 8),
36164 => conv_std_logic_vector(37, 8),
36165 => conv_std_logic_vector(38, 8),
36166 => conv_std_logic_vector(38, 8),
36167 => conv_std_logic_vector(39, 8),
36168 => conv_std_logic_vector(39, 8),
36169 => conv_std_logic_vector(40, 8),
36170 => conv_std_logic_vector(40, 8),
36171 => conv_std_logic_vector(41, 8),
36172 => conv_std_logic_vector(41, 8),
36173 => conv_std_logic_vector(42, 8),
36174 => conv_std_logic_vector(42, 8),
36175 => conv_std_logic_vector(43, 8),
36176 => conv_std_logic_vector(44, 8),
36177 => conv_std_logic_vector(44, 8),
36178 => conv_std_logic_vector(45, 8),
36179 => conv_std_logic_vector(45, 8),
36180 => conv_std_logic_vector(46, 8),
36181 => conv_std_logic_vector(46, 8),
36182 => conv_std_logic_vector(47, 8),
36183 => conv_std_logic_vector(47, 8),
36184 => conv_std_logic_vector(48, 8),
36185 => conv_std_logic_vector(49, 8),
36186 => conv_std_logic_vector(49, 8),
36187 => conv_std_logic_vector(50, 8),
36188 => conv_std_logic_vector(50, 8),
36189 => conv_std_logic_vector(51, 8),
36190 => conv_std_logic_vector(51, 8),
36191 => conv_std_logic_vector(52, 8),
36192 => conv_std_logic_vector(52, 8),
36193 => conv_std_logic_vector(53, 8),
36194 => conv_std_logic_vector(53, 8),
36195 => conv_std_logic_vector(54, 8),
36196 => conv_std_logic_vector(55, 8),
36197 => conv_std_logic_vector(55, 8),
36198 => conv_std_logic_vector(56, 8),
36199 => conv_std_logic_vector(56, 8),
36200 => conv_std_logic_vector(57, 8),
36201 => conv_std_logic_vector(57, 8),
36202 => conv_std_logic_vector(58, 8),
36203 => conv_std_logic_vector(58, 8),
36204 => conv_std_logic_vector(59, 8),
36205 => conv_std_logic_vector(60, 8),
36206 => conv_std_logic_vector(60, 8),
36207 => conv_std_logic_vector(61, 8),
36208 => conv_std_logic_vector(61, 8),
36209 => conv_std_logic_vector(62, 8),
36210 => conv_std_logic_vector(62, 8),
36211 => conv_std_logic_vector(63, 8),
36212 => conv_std_logic_vector(63, 8),
36213 => conv_std_logic_vector(64, 8),
36214 => conv_std_logic_vector(64, 8),
36215 => conv_std_logic_vector(65, 8),
36216 => conv_std_logic_vector(66, 8),
36217 => conv_std_logic_vector(66, 8),
36218 => conv_std_logic_vector(67, 8),
36219 => conv_std_logic_vector(67, 8),
36220 => conv_std_logic_vector(68, 8),
36221 => conv_std_logic_vector(68, 8),
36222 => conv_std_logic_vector(69, 8),
36223 => conv_std_logic_vector(69, 8),
36224 => conv_std_logic_vector(70, 8),
36225 => conv_std_logic_vector(71, 8),
36226 => conv_std_logic_vector(71, 8),
36227 => conv_std_logic_vector(72, 8),
36228 => conv_std_logic_vector(72, 8),
36229 => conv_std_logic_vector(73, 8),
36230 => conv_std_logic_vector(73, 8),
36231 => conv_std_logic_vector(74, 8),
36232 => conv_std_logic_vector(74, 8),
36233 => conv_std_logic_vector(75, 8),
36234 => conv_std_logic_vector(76, 8),
36235 => conv_std_logic_vector(76, 8),
36236 => conv_std_logic_vector(77, 8),
36237 => conv_std_logic_vector(77, 8),
36238 => conv_std_logic_vector(78, 8),
36239 => conv_std_logic_vector(78, 8),
36240 => conv_std_logic_vector(79, 8),
36241 => conv_std_logic_vector(79, 8),
36242 => conv_std_logic_vector(80, 8),
36243 => conv_std_logic_vector(80, 8),
36244 => conv_std_logic_vector(81, 8),
36245 => conv_std_logic_vector(82, 8),
36246 => conv_std_logic_vector(82, 8),
36247 => conv_std_logic_vector(83, 8),
36248 => conv_std_logic_vector(83, 8),
36249 => conv_std_logic_vector(84, 8),
36250 => conv_std_logic_vector(84, 8),
36251 => conv_std_logic_vector(85, 8),
36252 => conv_std_logic_vector(85, 8),
36253 => conv_std_logic_vector(86, 8),
36254 => conv_std_logic_vector(87, 8),
36255 => conv_std_logic_vector(87, 8),
36256 => conv_std_logic_vector(88, 8),
36257 => conv_std_logic_vector(88, 8),
36258 => conv_std_logic_vector(89, 8),
36259 => conv_std_logic_vector(89, 8),
36260 => conv_std_logic_vector(90, 8),
36261 => conv_std_logic_vector(90, 8),
36262 => conv_std_logic_vector(91, 8),
36263 => conv_std_logic_vector(91, 8),
36264 => conv_std_logic_vector(92, 8),
36265 => conv_std_logic_vector(93, 8),
36266 => conv_std_logic_vector(93, 8),
36267 => conv_std_logic_vector(94, 8),
36268 => conv_std_logic_vector(94, 8),
36269 => conv_std_logic_vector(95, 8),
36270 => conv_std_logic_vector(95, 8),
36271 => conv_std_logic_vector(96, 8),
36272 => conv_std_logic_vector(96, 8),
36273 => conv_std_logic_vector(97, 8),
36274 => conv_std_logic_vector(98, 8),
36275 => conv_std_logic_vector(98, 8),
36276 => conv_std_logic_vector(99, 8),
36277 => conv_std_logic_vector(99, 8),
36278 => conv_std_logic_vector(100, 8),
36279 => conv_std_logic_vector(100, 8),
36280 => conv_std_logic_vector(101, 8),
36281 => conv_std_logic_vector(101, 8),
36282 => conv_std_logic_vector(102, 8),
36283 => conv_std_logic_vector(102, 8),
36284 => conv_std_logic_vector(103, 8),
36285 => conv_std_logic_vector(104, 8),
36286 => conv_std_logic_vector(104, 8),
36287 => conv_std_logic_vector(105, 8),
36288 => conv_std_logic_vector(105, 8),
36289 => conv_std_logic_vector(106, 8),
36290 => conv_std_logic_vector(106, 8),
36291 => conv_std_logic_vector(107, 8),
36292 => conv_std_logic_vector(107, 8),
36293 => conv_std_logic_vector(108, 8),
36294 => conv_std_logic_vector(109, 8),
36295 => conv_std_logic_vector(109, 8),
36296 => conv_std_logic_vector(110, 8),
36297 => conv_std_logic_vector(110, 8),
36298 => conv_std_logic_vector(111, 8),
36299 => conv_std_logic_vector(111, 8),
36300 => conv_std_logic_vector(112, 8),
36301 => conv_std_logic_vector(112, 8),
36302 => conv_std_logic_vector(113, 8),
36303 => conv_std_logic_vector(114, 8),
36304 => conv_std_logic_vector(114, 8),
36305 => conv_std_logic_vector(115, 8),
36306 => conv_std_logic_vector(115, 8),
36307 => conv_std_logic_vector(116, 8),
36308 => conv_std_logic_vector(116, 8),
36309 => conv_std_logic_vector(117, 8),
36310 => conv_std_logic_vector(117, 8),
36311 => conv_std_logic_vector(118, 8),
36312 => conv_std_logic_vector(118, 8),
36313 => conv_std_logic_vector(119, 8),
36314 => conv_std_logic_vector(120, 8),
36315 => conv_std_logic_vector(120, 8),
36316 => conv_std_logic_vector(121, 8),
36317 => conv_std_logic_vector(121, 8),
36318 => conv_std_logic_vector(122, 8),
36319 => conv_std_logic_vector(122, 8),
36320 => conv_std_logic_vector(123, 8),
36321 => conv_std_logic_vector(123, 8),
36322 => conv_std_logic_vector(124, 8),
36323 => conv_std_logic_vector(125, 8),
36324 => conv_std_logic_vector(125, 8),
36325 => conv_std_logic_vector(126, 8),
36326 => conv_std_logic_vector(126, 8),
36327 => conv_std_logic_vector(127, 8),
36328 => conv_std_logic_vector(127, 8),
36329 => conv_std_logic_vector(128, 8),
36330 => conv_std_logic_vector(128, 8),
36331 => conv_std_logic_vector(129, 8),
36332 => conv_std_logic_vector(129, 8),
36333 => conv_std_logic_vector(130, 8),
36334 => conv_std_logic_vector(131, 8),
36335 => conv_std_logic_vector(131, 8),
36336 => conv_std_logic_vector(132, 8),
36337 => conv_std_logic_vector(132, 8),
36338 => conv_std_logic_vector(133, 8),
36339 => conv_std_logic_vector(133, 8),
36340 => conv_std_logic_vector(134, 8),
36341 => conv_std_logic_vector(134, 8),
36342 => conv_std_logic_vector(135, 8),
36343 => conv_std_logic_vector(136, 8),
36344 => conv_std_logic_vector(136, 8),
36345 => conv_std_logic_vector(137, 8),
36346 => conv_std_logic_vector(137, 8),
36347 => conv_std_logic_vector(138, 8),
36348 => conv_std_logic_vector(138, 8),
36349 => conv_std_logic_vector(139, 8),
36350 => conv_std_logic_vector(139, 8),
36351 => conv_std_logic_vector(140, 8),
36352 => conv_std_logic_vector(0, 8),
36353 => conv_std_logic_vector(0, 8),
36354 => conv_std_logic_vector(1, 8),
36355 => conv_std_logic_vector(1, 8),
36356 => conv_std_logic_vector(2, 8),
36357 => conv_std_logic_vector(2, 8),
36358 => conv_std_logic_vector(3, 8),
36359 => conv_std_logic_vector(3, 8),
36360 => conv_std_logic_vector(4, 8),
36361 => conv_std_logic_vector(4, 8),
36362 => conv_std_logic_vector(5, 8),
36363 => conv_std_logic_vector(6, 8),
36364 => conv_std_logic_vector(6, 8),
36365 => conv_std_logic_vector(7, 8),
36366 => conv_std_logic_vector(7, 8),
36367 => conv_std_logic_vector(8, 8),
36368 => conv_std_logic_vector(8, 8),
36369 => conv_std_logic_vector(9, 8),
36370 => conv_std_logic_vector(9, 8),
36371 => conv_std_logic_vector(10, 8),
36372 => conv_std_logic_vector(11, 8),
36373 => conv_std_logic_vector(11, 8),
36374 => conv_std_logic_vector(12, 8),
36375 => conv_std_logic_vector(12, 8),
36376 => conv_std_logic_vector(13, 8),
36377 => conv_std_logic_vector(13, 8),
36378 => conv_std_logic_vector(14, 8),
36379 => conv_std_logic_vector(14, 8),
36380 => conv_std_logic_vector(15, 8),
36381 => conv_std_logic_vector(16, 8),
36382 => conv_std_logic_vector(16, 8),
36383 => conv_std_logic_vector(17, 8),
36384 => conv_std_logic_vector(17, 8),
36385 => conv_std_logic_vector(18, 8),
36386 => conv_std_logic_vector(18, 8),
36387 => conv_std_logic_vector(19, 8),
36388 => conv_std_logic_vector(19, 8),
36389 => conv_std_logic_vector(20, 8),
36390 => conv_std_logic_vector(21, 8),
36391 => conv_std_logic_vector(21, 8),
36392 => conv_std_logic_vector(22, 8),
36393 => conv_std_logic_vector(22, 8),
36394 => conv_std_logic_vector(23, 8),
36395 => conv_std_logic_vector(23, 8),
36396 => conv_std_logic_vector(24, 8),
36397 => conv_std_logic_vector(24, 8),
36398 => conv_std_logic_vector(25, 8),
36399 => conv_std_logic_vector(26, 8),
36400 => conv_std_logic_vector(26, 8),
36401 => conv_std_logic_vector(27, 8),
36402 => conv_std_logic_vector(27, 8),
36403 => conv_std_logic_vector(28, 8),
36404 => conv_std_logic_vector(28, 8),
36405 => conv_std_logic_vector(29, 8),
36406 => conv_std_logic_vector(29, 8),
36407 => conv_std_logic_vector(30, 8),
36408 => conv_std_logic_vector(31, 8),
36409 => conv_std_logic_vector(31, 8),
36410 => conv_std_logic_vector(32, 8),
36411 => conv_std_logic_vector(32, 8),
36412 => conv_std_logic_vector(33, 8),
36413 => conv_std_logic_vector(33, 8),
36414 => conv_std_logic_vector(34, 8),
36415 => conv_std_logic_vector(34, 8),
36416 => conv_std_logic_vector(35, 8),
36417 => conv_std_logic_vector(36, 8),
36418 => conv_std_logic_vector(36, 8),
36419 => conv_std_logic_vector(37, 8),
36420 => conv_std_logic_vector(37, 8),
36421 => conv_std_logic_vector(38, 8),
36422 => conv_std_logic_vector(38, 8),
36423 => conv_std_logic_vector(39, 8),
36424 => conv_std_logic_vector(39, 8),
36425 => conv_std_logic_vector(40, 8),
36426 => conv_std_logic_vector(41, 8),
36427 => conv_std_logic_vector(41, 8),
36428 => conv_std_logic_vector(42, 8),
36429 => conv_std_logic_vector(42, 8),
36430 => conv_std_logic_vector(43, 8),
36431 => conv_std_logic_vector(43, 8),
36432 => conv_std_logic_vector(44, 8),
36433 => conv_std_logic_vector(44, 8),
36434 => conv_std_logic_vector(45, 8),
36435 => conv_std_logic_vector(46, 8),
36436 => conv_std_logic_vector(46, 8),
36437 => conv_std_logic_vector(47, 8),
36438 => conv_std_logic_vector(47, 8),
36439 => conv_std_logic_vector(48, 8),
36440 => conv_std_logic_vector(48, 8),
36441 => conv_std_logic_vector(49, 8),
36442 => conv_std_logic_vector(49, 8),
36443 => conv_std_logic_vector(50, 8),
36444 => conv_std_logic_vector(51, 8),
36445 => conv_std_logic_vector(51, 8),
36446 => conv_std_logic_vector(52, 8),
36447 => conv_std_logic_vector(52, 8),
36448 => conv_std_logic_vector(53, 8),
36449 => conv_std_logic_vector(53, 8),
36450 => conv_std_logic_vector(54, 8),
36451 => conv_std_logic_vector(54, 8),
36452 => conv_std_logic_vector(55, 8),
36453 => conv_std_logic_vector(56, 8),
36454 => conv_std_logic_vector(56, 8),
36455 => conv_std_logic_vector(57, 8),
36456 => conv_std_logic_vector(57, 8),
36457 => conv_std_logic_vector(58, 8),
36458 => conv_std_logic_vector(58, 8),
36459 => conv_std_logic_vector(59, 8),
36460 => conv_std_logic_vector(59, 8),
36461 => conv_std_logic_vector(60, 8),
36462 => conv_std_logic_vector(61, 8),
36463 => conv_std_logic_vector(61, 8),
36464 => conv_std_logic_vector(62, 8),
36465 => conv_std_logic_vector(62, 8),
36466 => conv_std_logic_vector(63, 8),
36467 => conv_std_logic_vector(63, 8),
36468 => conv_std_logic_vector(64, 8),
36469 => conv_std_logic_vector(64, 8),
36470 => conv_std_logic_vector(65, 8),
36471 => conv_std_logic_vector(66, 8),
36472 => conv_std_logic_vector(66, 8),
36473 => conv_std_logic_vector(67, 8),
36474 => conv_std_logic_vector(67, 8),
36475 => conv_std_logic_vector(68, 8),
36476 => conv_std_logic_vector(68, 8),
36477 => conv_std_logic_vector(69, 8),
36478 => conv_std_logic_vector(69, 8),
36479 => conv_std_logic_vector(70, 8),
36480 => conv_std_logic_vector(71, 8),
36481 => conv_std_logic_vector(71, 8),
36482 => conv_std_logic_vector(72, 8),
36483 => conv_std_logic_vector(72, 8),
36484 => conv_std_logic_vector(73, 8),
36485 => conv_std_logic_vector(73, 8),
36486 => conv_std_logic_vector(74, 8),
36487 => conv_std_logic_vector(74, 8),
36488 => conv_std_logic_vector(75, 8),
36489 => conv_std_logic_vector(75, 8),
36490 => conv_std_logic_vector(76, 8),
36491 => conv_std_logic_vector(77, 8),
36492 => conv_std_logic_vector(77, 8),
36493 => conv_std_logic_vector(78, 8),
36494 => conv_std_logic_vector(78, 8),
36495 => conv_std_logic_vector(79, 8),
36496 => conv_std_logic_vector(79, 8),
36497 => conv_std_logic_vector(80, 8),
36498 => conv_std_logic_vector(80, 8),
36499 => conv_std_logic_vector(81, 8),
36500 => conv_std_logic_vector(82, 8),
36501 => conv_std_logic_vector(82, 8),
36502 => conv_std_logic_vector(83, 8),
36503 => conv_std_logic_vector(83, 8),
36504 => conv_std_logic_vector(84, 8),
36505 => conv_std_logic_vector(84, 8),
36506 => conv_std_logic_vector(85, 8),
36507 => conv_std_logic_vector(85, 8),
36508 => conv_std_logic_vector(86, 8),
36509 => conv_std_logic_vector(87, 8),
36510 => conv_std_logic_vector(87, 8),
36511 => conv_std_logic_vector(88, 8),
36512 => conv_std_logic_vector(88, 8),
36513 => conv_std_logic_vector(89, 8),
36514 => conv_std_logic_vector(89, 8),
36515 => conv_std_logic_vector(90, 8),
36516 => conv_std_logic_vector(90, 8),
36517 => conv_std_logic_vector(91, 8),
36518 => conv_std_logic_vector(92, 8),
36519 => conv_std_logic_vector(92, 8),
36520 => conv_std_logic_vector(93, 8),
36521 => conv_std_logic_vector(93, 8),
36522 => conv_std_logic_vector(94, 8),
36523 => conv_std_logic_vector(94, 8),
36524 => conv_std_logic_vector(95, 8),
36525 => conv_std_logic_vector(95, 8),
36526 => conv_std_logic_vector(96, 8),
36527 => conv_std_logic_vector(97, 8),
36528 => conv_std_logic_vector(97, 8),
36529 => conv_std_logic_vector(98, 8),
36530 => conv_std_logic_vector(98, 8),
36531 => conv_std_logic_vector(99, 8),
36532 => conv_std_logic_vector(99, 8),
36533 => conv_std_logic_vector(100, 8),
36534 => conv_std_logic_vector(100, 8),
36535 => conv_std_logic_vector(101, 8),
36536 => conv_std_logic_vector(102, 8),
36537 => conv_std_logic_vector(102, 8),
36538 => conv_std_logic_vector(103, 8),
36539 => conv_std_logic_vector(103, 8),
36540 => conv_std_logic_vector(104, 8),
36541 => conv_std_logic_vector(104, 8),
36542 => conv_std_logic_vector(105, 8),
36543 => conv_std_logic_vector(105, 8),
36544 => conv_std_logic_vector(106, 8),
36545 => conv_std_logic_vector(107, 8),
36546 => conv_std_logic_vector(107, 8),
36547 => conv_std_logic_vector(108, 8),
36548 => conv_std_logic_vector(108, 8),
36549 => conv_std_logic_vector(109, 8),
36550 => conv_std_logic_vector(109, 8),
36551 => conv_std_logic_vector(110, 8),
36552 => conv_std_logic_vector(110, 8),
36553 => conv_std_logic_vector(111, 8),
36554 => conv_std_logic_vector(112, 8),
36555 => conv_std_logic_vector(112, 8),
36556 => conv_std_logic_vector(113, 8),
36557 => conv_std_logic_vector(113, 8),
36558 => conv_std_logic_vector(114, 8),
36559 => conv_std_logic_vector(114, 8),
36560 => conv_std_logic_vector(115, 8),
36561 => conv_std_logic_vector(115, 8),
36562 => conv_std_logic_vector(116, 8),
36563 => conv_std_logic_vector(117, 8),
36564 => conv_std_logic_vector(117, 8),
36565 => conv_std_logic_vector(118, 8),
36566 => conv_std_logic_vector(118, 8),
36567 => conv_std_logic_vector(119, 8),
36568 => conv_std_logic_vector(119, 8),
36569 => conv_std_logic_vector(120, 8),
36570 => conv_std_logic_vector(120, 8),
36571 => conv_std_logic_vector(121, 8),
36572 => conv_std_logic_vector(122, 8),
36573 => conv_std_logic_vector(122, 8),
36574 => conv_std_logic_vector(123, 8),
36575 => conv_std_logic_vector(123, 8),
36576 => conv_std_logic_vector(124, 8),
36577 => conv_std_logic_vector(124, 8),
36578 => conv_std_logic_vector(125, 8),
36579 => conv_std_logic_vector(125, 8),
36580 => conv_std_logic_vector(126, 8),
36581 => conv_std_logic_vector(127, 8),
36582 => conv_std_logic_vector(127, 8),
36583 => conv_std_logic_vector(128, 8),
36584 => conv_std_logic_vector(128, 8),
36585 => conv_std_logic_vector(129, 8),
36586 => conv_std_logic_vector(129, 8),
36587 => conv_std_logic_vector(130, 8),
36588 => conv_std_logic_vector(130, 8),
36589 => conv_std_logic_vector(131, 8),
36590 => conv_std_logic_vector(132, 8),
36591 => conv_std_logic_vector(132, 8),
36592 => conv_std_logic_vector(133, 8),
36593 => conv_std_logic_vector(133, 8),
36594 => conv_std_logic_vector(134, 8),
36595 => conv_std_logic_vector(134, 8),
36596 => conv_std_logic_vector(135, 8),
36597 => conv_std_logic_vector(135, 8),
36598 => conv_std_logic_vector(136, 8),
36599 => conv_std_logic_vector(137, 8),
36600 => conv_std_logic_vector(137, 8),
36601 => conv_std_logic_vector(138, 8),
36602 => conv_std_logic_vector(138, 8),
36603 => conv_std_logic_vector(139, 8),
36604 => conv_std_logic_vector(139, 8),
36605 => conv_std_logic_vector(140, 8),
36606 => conv_std_logic_vector(140, 8),
36607 => conv_std_logic_vector(141, 8),
36608 => conv_std_logic_vector(0, 8),
36609 => conv_std_logic_vector(0, 8),
36610 => conv_std_logic_vector(1, 8),
36611 => conv_std_logic_vector(1, 8),
36612 => conv_std_logic_vector(2, 8),
36613 => conv_std_logic_vector(2, 8),
36614 => conv_std_logic_vector(3, 8),
36615 => conv_std_logic_vector(3, 8),
36616 => conv_std_logic_vector(4, 8),
36617 => conv_std_logic_vector(5, 8),
36618 => conv_std_logic_vector(5, 8),
36619 => conv_std_logic_vector(6, 8),
36620 => conv_std_logic_vector(6, 8),
36621 => conv_std_logic_vector(7, 8),
36622 => conv_std_logic_vector(7, 8),
36623 => conv_std_logic_vector(8, 8),
36624 => conv_std_logic_vector(8, 8),
36625 => conv_std_logic_vector(9, 8),
36626 => conv_std_logic_vector(10, 8),
36627 => conv_std_logic_vector(10, 8),
36628 => conv_std_logic_vector(11, 8),
36629 => conv_std_logic_vector(11, 8),
36630 => conv_std_logic_vector(12, 8),
36631 => conv_std_logic_vector(12, 8),
36632 => conv_std_logic_vector(13, 8),
36633 => conv_std_logic_vector(13, 8),
36634 => conv_std_logic_vector(14, 8),
36635 => conv_std_logic_vector(15, 8),
36636 => conv_std_logic_vector(15, 8),
36637 => conv_std_logic_vector(16, 8),
36638 => conv_std_logic_vector(16, 8),
36639 => conv_std_logic_vector(17, 8),
36640 => conv_std_logic_vector(17, 8),
36641 => conv_std_logic_vector(18, 8),
36642 => conv_std_logic_vector(18, 8),
36643 => conv_std_logic_vector(19, 8),
36644 => conv_std_logic_vector(20, 8),
36645 => conv_std_logic_vector(20, 8),
36646 => conv_std_logic_vector(21, 8),
36647 => conv_std_logic_vector(21, 8),
36648 => conv_std_logic_vector(22, 8),
36649 => conv_std_logic_vector(22, 8),
36650 => conv_std_logic_vector(23, 8),
36651 => conv_std_logic_vector(24, 8),
36652 => conv_std_logic_vector(24, 8),
36653 => conv_std_logic_vector(25, 8),
36654 => conv_std_logic_vector(25, 8),
36655 => conv_std_logic_vector(26, 8),
36656 => conv_std_logic_vector(26, 8),
36657 => conv_std_logic_vector(27, 8),
36658 => conv_std_logic_vector(27, 8),
36659 => conv_std_logic_vector(28, 8),
36660 => conv_std_logic_vector(29, 8),
36661 => conv_std_logic_vector(29, 8),
36662 => conv_std_logic_vector(30, 8),
36663 => conv_std_logic_vector(30, 8),
36664 => conv_std_logic_vector(31, 8),
36665 => conv_std_logic_vector(31, 8),
36666 => conv_std_logic_vector(32, 8),
36667 => conv_std_logic_vector(32, 8),
36668 => conv_std_logic_vector(33, 8),
36669 => conv_std_logic_vector(34, 8),
36670 => conv_std_logic_vector(34, 8),
36671 => conv_std_logic_vector(35, 8),
36672 => conv_std_logic_vector(35, 8),
36673 => conv_std_logic_vector(36, 8),
36674 => conv_std_logic_vector(36, 8),
36675 => conv_std_logic_vector(37, 8),
36676 => conv_std_logic_vector(37, 8),
36677 => conv_std_logic_vector(38, 8),
36678 => conv_std_logic_vector(39, 8),
36679 => conv_std_logic_vector(39, 8),
36680 => conv_std_logic_vector(40, 8),
36681 => conv_std_logic_vector(40, 8),
36682 => conv_std_logic_vector(41, 8),
36683 => conv_std_logic_vector(41, 8),
36684 => conv_std_logic_vector(42, 8),
36685 => conv_std_logic_vector(43, 8),
36686 => conv_std_logic_vector(43, 8),
36687 => conv_std_logic_vector(44, 8),
36688 => conv_std_logic_vector(44, 8),
36689 => conv_std_logic_vector(45, 8),
36690 => conv_std_logic_vector(45, 8),
36691 => conv_std_logic_vector(46, 8),
36692 => conv_std_logic_vector(46, 8),
36693 => conv_std_logic_vector(47, 8),
36694 => conv_std_logic_vector(48, 8),
36695 => conv_std_logic_vector(48, 8),
36696 => conv_std_logic_vector(49, 8),
36697 => conv_std_logic_vector(49, 8),
36698 => conv_std_logic_vector(50, 8),
36699 => conv_std_logic_vector(50, 8),
36700 => conv_std_logic_vector(51, 8),
36701 => conv_std_logic_vector(51, 8),
36702 => conv_std_logic_vector(52, 8),
36703 => conv_std_logic_vector(53, 8),
36704 => conv_std_logic_vector(53, 8),
36705 => conv_std_logic_vector(54, 8),
36706 => conv_std_logic_vector(54, 8),
36707 => conv_std_logic_vector(55, 8),
36708 => conv_std_logic_vector(55, 8),
36709 => conv_std_logic_vector(56, 8),
36710 => conv_std_logic_vector(56, 8),
36711 => conv_std_logic_vector(57, 8),
36712 => conv_std_logic_vector(58, 8),
36713 => conv_std_logic_vector(58, 8),
36714 => conv_std_logic_vector(59, 8),
36715 => conv_std_logic_vector(59, 8),
36716 => conv_std_logic_vector(60, 8),
36717 => conv_std_logic_vector(60, 8),
36718 => conv_std_logic_vector(61, 8),
36719 => conv_std_logic_vector(62, 8),
36720 => conv_std_logic_vector(62, 8),
36721 => conv_std_logic_vector(63, 8),
36722 => conv_std_logic_vector(63, 8),
36723 => conv_std_logic_vector(64, 8),
36724 => conv_std_logic_vector(64, 8),
36725 => conv_std_logic_vector(65, 8),
36726 => conv_std_logic_vector(65, 8),
36727 => conv_std_logic_vector(66, 8),
36728 => conv_std_logic_vector(67, 8),
36729 => conv_std_logic_vector(67, 8),
36730 => conv_std_logic_vector(68, 8),
36731 => conv_std_logic_vector(68, 8),
36732 => conv_std_logic_vector(69, 8),
36733 => conv_std_logic_vector(69, 8),
36734 => conv_std_logic_vector(70, 8),
36735 => conv_std_logic_vector(70, 8),
36736 => conv_std_logic_vector(71, 8),
36737 => conv_std_logic_vector(72, 8),
36738 => conv_std_logic_vector(72, 8),
36739 => conv_std_logic_vector(73, 8),
36740 => conv_std_logic_vector(73, 8),
36741 => conv_std_logic_vector(74, 8),
36742 => conv_std_logic_vector(74, 8),
36743 => conv_std_logic_vector(75, 8),
36744 => conv_std_logic_vector(75, 8),
36745 => conv_std_logic_vector(76, 8),
36746 => conv_std_logic_vector(77, 8),
36747 => conv_std_logic_vector(77, 8),
36748 => conv_std_logic_vector(78, 8),
36749 => conv_std_logic_vector(78, 8),
36750 => conv_std_logic_vector(79, 8),
36751 => conv_std_logic_vector(79, 8),
36752 => conv_std_logic_vector(80, 8),
36753 => conv_std_logic_vector(80, 8),
36754 => conv_std_logic_vector(81, 8),
36755 => conv_std_logic_vector(82, 8),
36756 => conv_std_logic_vector(82, 8),
36757 => conv_std_logic_vector(83, 8),
36758 => conv_std_logic_vector(83, 8),
36759 => conv_std_logic_vector(84, 8),
36760 => conv_std_logic_vector(84, 8),
36761 => conv_std_logic_vector(85, 8),
36762 => conv_std_logic_vector(86, 8),
36763 => conv_std_logic_vector(86, 8),
36764 => conv_std_logic_vector(87, 8),
36765 => conv_std_logic_vector(87, 8),
36766 => conv_std_logic_vector(88, 8),
36767 => conv_std_logic_vector(88, 8),
36768 => conv_std_logic_vector(89, 8),
36769 => conv_std_logic_vector(89, 8),
36770 => conv_std_logic_vector(90, 8),
36771 => conv_std_logic_vector(91, 8),
36772 => conv_std_logic_vector(91, 8),
36773 => conv_std_logic_vector(92, 8),
36774 => conv_std_logic_vector(92, 8),
36775 => conv_std_logic_vector(93, 8),
36776 => conv_std_logic_vector(93, 8),
36777 => conv_std_logic_vector(94, 8),
36778 => conv_std_logic_vector(94, 8),
36779 => conv_std_logic_vector(95, 8),
36780 => conv_std_logic_vector(96, 8),
36781 => conv_std_logic_vector(96, 8),
36782 => conv_std_logic_vector(97, 8),
36783 => conv_std_logic_vector(97, 8),
36784 => conv_std_logic_vector(98, 8),
36785 => conv_std_logic_vector(98, 8),
36786 => conv_std_logic_vector(99, 8),
36787 => conv_std_logic_vector(99, 8),
36788 => conv_std_logic_vector(100, 8),
36789 => conv_std_logic_vector(101, 8),
36790 => conv_std_logic_vector(101, 8),
36791 => conv_std_logic_vector(102, 8),
36792 => conv_std_logic_vector(102, 8),
36793 => conv_std_logic_vector(103, 8),
36794 => conv_std_logic_vector(103, 8),
36795 => conv_std_logic_vector(104, 8),
36796 => conv_std_logic_vector(105, 8),
36797 => conv_std_logic_vector(105, 8),
36798 => conv_std_logic_vector(106, 8),
36799 => conv_std_logic_vector(106, 8),
36800 => conv_std_logic_vector(107, 8),
36801 => conv_std_logic_vector(107, 8),
36802 => conv_std_logic_vector(108, 8),
36803 => conv_std_logic_vector(108, 8),
36804 => conv_std_logic_vector(109, 8),
36805 => conv_std_logic_vector(110, 8),
36806 => conv_std_logic_vector(110, 8),
36807 => conv_std_logic_vector(111, 8),
36808 => conv_std_logic_vector(111, 8),
36809 => conv_std_logic_vector(112, 8),
36810 => conv_std_logic_vector(112, 8),
36811 => conv_std_logic_vector(113, 8),
36812 => conv_std_logic_vector(113, 8),
36813 => conv_std_logic_vector(114, 8),
36814 => conv_std_logic_vector(115, 8),
36815 => conv_std_logic_vector(115, 8),
36816 => conv_std_logic_vector(116, 8),
36817 => conv_std_logic_vector(116, 8),
36818 => conv_std_logic_vector(117, 8),
36819 => conv_std_logic_vector(117, 8),
36820 => conv_std_logic_vector(118, 8),
36821 => conv_std_logic_vector(118, 8),
36822 => conv_std_logic_vector(119, 8),
36823 => conv_std_logic_vector(120, 8),
36824 => conv_std_logic_vector(120, 8),
36825 => conv_std_logic_vector(121, 8),
36826 => conv_std_logic_vector(121, 8),
36827 => conv_std_logic_vector(122, 8),
36828 => conv_std_logic_vector(122, 8),
36829 => conv_std_logic_vector(123, 8),
36830 => conv_std_logic_vector(124, 8),
36831 => conv_std_logic_vector(124, 8),
36832 => conv_std_logic_vector(125, 8),
36833 => conv_std_logic_vector(125, 8),
36834 => conv_std_logic_vector(126, 8),
36835 => conv_std_logic_vector(126, 8),
36836 => conv_std_logic_vector(127, 8),
36837 => conv_std_logic_vector(127, 8),
36838 => conv_std_logic_vector(128, 8),
36839 => conv_std_logic_vector(129, 8),
36840 => conv_std_logic_vector(129, 8),
36841 => conv_std_logic_vector(130, 8),
36842 => conv_std_logic_vector(130, 8),
36843 => conv_std_logic_vector(131, 8),
36844 => conv_std_logic_vector(131, 8),
36845 => conv_std_logic_vector(132, 8),
36846 => conv_std_logic_vector(132, 8),
36847 => conv_std_logic_vector(133, 8),
36848 => conv_std_logic_vector(134, 8),
36849 => conv_std_logic_vector(134, 8),
36850 => conv_std_logic_vector(135, 8),
36851 => conv_std_logic_vector(135, 8),
36852 => conv_std_logic_vector(136, 8),
36853 => conv_std_logic_vector(136, 8),
36854 => conv_std_logic_vector(137, 8),
36855 => conv_std_logic_vector(137, 8),
36856 => conv_std_logic_vector(138, 8),
36857 => conv_std_logic_vector(139, 8),
36858 => conv_std_logic_vector(139, 8),
36859 => conv_std_logic_vector(140, 8),
36860 => conv_std_logic_vector(140, 8),
36861 => conv_std_logic_vector(141, 8),
36862 => conv_std_logic_vector(141, 8),
36863 => conv_std_logic_vector(142, 8),
36864 => conv_std_logic_vector(0, 8),
36865 => conv_std_logic_vector(0, 8),
36866 => conv_std_logic_vector(1, 8),
36867 => conv_std_logic_vector(1, 8),
36868 => conv_std_logic_vector(2, 8),
36869 => conv_std_logic_vector(2, 8),
36870 => conv_std_logic_vector(3, 8),
36871 => conv_std_logic_vector(3, 8),
36872 => conv_std_logic_vector(4, 8),
36873 => conv_std_logic_vector(5, 8),
36874 => conv_std_logic_vector(5, 8),
36875 => conv_std_logic_vector(6, 8),
36876 => conv_std_logic_vector(6, 8),
36877 => conv_std_logic_vector(7, 8),
36878 => conv_std_logic_vector(7, 8),
36879 => conv_std_logic_vector(8, 8),
36880 => conv_std_logic_vector(9, 8),
36881 => conv_std_logic_vector(9, 8),
36882 => conv_std_logic_vector(10, 8),
36883 => conv_std_logic_vector(10, 8),
36884 => conv_std_logic_vector(11, 8),
36885 => conv_std_logic_vector(11, 8),
36886 => conv_std_logic_vector(12, 8),
36887 => conv_std_logic_vector(12, 8),
36888 => conv_std_logic_vector(13, 8),
36889 => conv_std_logic_vector(14, 8),
36890 => conv_std_logic_vector(14, 8),
36891 => conv_std_logic_vector(15, 8),
36892 => conv_std_logic_vector(15, 8),
36893 => conv_std_logic_vector(16, 8),
36894 => conv_std_logic_vector(16, 8),
36895 => conv_std_logic_vector(17, 8),
36896 => conv_std_logic_vector(18, 8),
36897 => conv_std_logic_vector(18, 8),
36898 => conv_std_logic_vector(19, 8),
36899 => conv_std_logic_vector(19, 8),
36900 => conv_std_logic_vector(20, 8),
36901 => conv_std_logic_vector(20, 8),
36902 => conv_std_logic_vector(21, 8),
36903 => conv_std_logic_vector(21, 8),
36904 => conv_std_logic_vector(22, 8),
36905 => conv_std_logic_vector(23, 8),
36906 => conv_std_logic_vector(23, 8),
36907 => conv_std_logic_vector(24, 8),
36908 => conv_std_logic_vector(24, 8),
36909 => conv_std_logic_vector(25, 8),
36910 => conv_std_logic_vector(25, 8),
36911 => conv_std_logic_vector(26, 8),
36912 => conv_std_logic_vector(27, 8),
36913 => conv_std_logic_vector(27, 8),
36914 => conv_std_logic_vector(28, 8),
36915 => conv_std_logic_vector(28, 8),
36916 => conv_std_logic_vector(29, 8),
36917 => conv_std_logic_vector(29, 8),
36918 => conv_std_logic_vector(30, 8),
36919 => conv_std_logic_vector(30, 8),
36920 => conv_std_logic_vector(31, 8),
36921 => conv_std_logic_vector(32, 8),
36922 => conv_std_logic_vector(32, 8),
36923 => conv_std_logic_vector(33, 8),
36924 => conv_std_logic_vector(33, 8),
36925 => conv_std_logic_vector(34, 8),
36926 => conv_std_logic_vector(34, 8),
36927 => conv_std_logic_vector(35, 8),
36928 => conv_std_logic_vector(36, 8),
36929 => conv_std_logic_vector(36, 8),
36930 => conv_std_logic_vector(37, 8),
36931 => conv_std_logic_vector(37, 8),
36932 => conv_std_logic_vector(38, 8),
36933 => conv_std_logic_vector(38, 8),
36934 => conv_std_logic_vector(39, 8),
36935 => conv_std_logic_vector(39, 8),
36936 => conv_std_logic_vector(40, 8),
36937 => conv_std_logic_vector(41, 8),
36938 => conv_std_logic_vector(41, 8),
36939 => conv_std_logic_vector(42, 8),
36940 => conv_std_logic_vector(42, 8),
36941 => conv_std_logic_vector(43, 8),
36942 => conv_std_logic_vector(43, 8),
36943 => conv_std_logic_vector(44, 8),
36944 => conv_std_logic_vector(45, 8),
36945 => conv_std_logic_vector(45, 8),
36946 => conv_std_logic_vector(46, 8),
36947 => conv_std_logic_vector(46, 8),
36948 => conv_std_logic_vector(47, 8),
36949 => conv_std_logic_vector(47, 8),
36950 => conv_std_logic_vector(48, 8),
36951 => conv_std_logic_vector(48, 8),
36952 => conv_std_logic_vector(49, 8),
36953 => conv_std_logic_vector(50, 8),
36954 => conv_std_logic_vector(50, 8),
36955 => conv_std_logic_vector(51, 8),
36956 => conv_std_logic_vector(51, 8),
36957 => conv_std_logic_vector(52, 8),
36958 => conv_std_logic_vector(52, 8),
36959 => conv_std_logic_vector(53, 8),
36960 => conv_std_logic_vector(54, 8),
36961 => conv_std_logic_vector(54, 8),
36962 => conv_std_logic_vector(55, 8),
36963 => conv_std_logic_vector(55, 8),
36964 => conv_std_logic_vector(56, 8),
36965 => conv_std_logic_vector(56, 8),
36966 => conv_std_logic_vector(57, 8),
36967 => conv_std_logic_vector(57, 8),
36968 => conv_std_logic_vector(58, 8),
36969 => conv_std_logic_vector(59, 8),
36970 => conv_std_logic_vector(59, 8),
36971 => conv_std_logic_vector(60, 8),
36972 => conv_std_logic_vector(60, 8),
36973 => conv_std_logic_vector(61, 8),
36974 => conv_std_logic_vector(61, 8),
36975 => conv_std_logic_vector(62, 8),
36976 => conv_std_logic_vector(63, 8),
36977 => conv_std_logic_vector(63, 8),
36978 => conv_std_logic_vector(64, 8),
36979 => conv_std_logic_vector(64, 8),
36980 => conv_std_logic_vector(65, 8),
36981 => conv_std_logic_vector(65, 8),
36982 => conv_std_logic_vector(66, 8),
36983 => conv_std_logic_vector(66, 8),
36984 => conv_std_logic_vector(67, 8),
36985 => conv_std_logic_vector(68, 8),
36986 => conv_std_logic_vector(68, 8),
36987 => conv_std_logic_vector(69, 8),
36988 => conv_std_logic_vector(69, 8),
36989 => conv_std_logic_vector(70, 8),
36990 => conv_std_logic_vector(70, 8),
36991 => conv_std_logic_vector(71, 8),
36992 => conv_std_logic_vector(72, 8),
36993 => conv_std_logic_vector(72, 8),
36994 => conv_std_logic_vector(73, 8),
36995 => conv_std_logic_vector(73, 8),
36996 => conv_std_logic_vector(74, 8),
36997 => conv_std_logic_vector(74, 8),
36998 => conv_std_logic_vector(75, 8),
36999 => conv_std_logic_vector(75, 8),
37000 => conv_std_logic_vector(76, 8),
37001 => conv_std_logic_vector(77, 8),
37002 => conv_std_logic_vector(77, 8),
37003 => conv_std_logic_vector(78, 8),
37004 => conv_std_logic_vector(78, 8),
37005 => conv_std_logic_vector(79, 8),
37006 => conv_std_logic_vector(79, 8),
37007 => conv_std_logic_vector(80, 8),
37008 => conv_std_logic_vector(81, 8),
37009 => conv_std_logic_vector(81, 8),
37010 => conv_std_logic_vector(82, 8),
37011 => conv_std_logic_vector(82, 8),
37012 => conv_std_logic_vector(83, 8),
37013 => conv_std_logic_vector(83, 8),
37014 => conv_std_logic_vector(84, 8),
37015 => conv_std_logic_vector(84, 8),
37016 => conv_std_logic_vector(85, 8),
37017 => conv_std_logic_vector(86, 8),
37018 => conv_std_logic_vector(86, 8),
37019 => conv_std_logic_vector(87, 8),
37020 => conv_std_logic_vector(87, 8),
37021 => conv_std_logic_vector(88, 8),
37022 => conv_std_logic_vector(88, 8),
37023 => conv_std_logic_vector(89, 8),
37024 => conv_std_logic_vector(90, 8),
37025 => conv_std_logic_vector(90, 8),
37026 => conv_std_logic_vector(91, 8),
37027 => conv_std_logic_vector(91, 8),
37028 => conv_std_logic_vector(92, 8),
37029 => conv_std_logic_vector(92, 8),
37030 => conv_std_logic_vector(93, 8),
37031 => conv_std_logic_vector(93, 8),
37032 => conv_std_logic_vector(94, 8),
37033 => conv_std_logic_vector(95, 8),
37034 => conv_std_logic_vector(95, 8),
37035 => conv_std_logic_vector(96, 8),
37036 => conv_std_logic_vector(96, 8),
37037 => conv_std_logic_vector(97, 8),
37038 => conv_std_logic_vector(97, 8),
37039 => conv_std_logic_vector(98, 8),
37040 => conv_std_logic_vector(99, 8),
37041 => conv_std_logic_vector(99, 8),
37042 => conv_std_logic_vector(100, 8),
37043 => conv_std_logic_vector(100, 8),
37044 => conv_std_logic_vector(101, 8),
37045 => conv_std_logic_vector(101, 8),
37046 => conv_std_logic_vector(102, 8),
37047 => conv_std_logic_vector(102, 8),
37048 => conv_std_logic_vector(103, 8),
37049 => conv_std_logic_vector(104, 8),
37050 => conv_std_logic_vector(104, 8),
37051 => conv_std_logic_vector(105, 8),
37052 => conv_std_logic_vector(105, 8),
37053 => conv_std_logic_vector(106, 8),
37054 => conv_std_logic_vector(106, 8),
37055 => conv_std_logic_vector(107, 8),
37056 => conv_std_logic_vector(108, 8),
37057 => conv_std_logic_vector(108, 8),
37058 => conv_std_logic_vector(109, 8),
37059 => conv_std_logic_vector(109, 8),
37060 => conv_std_logic_vector(110, 8),
37061 => conv_std_logic_vector(110, 8),
37062 => conv_std_logic_vector(111, 8),
37063 => conv_std_logic_vector(111, 8),
37064 => conv_std_logic_vector(112, 8),
37065 => conv_std_logic_vector(113, 8),
37066 => conv_std_logic_vector(113, 8),
37067 => conv_std_logic_vector(114, 8),
37068 => conv_std_logic_vector(114, 8),
37069 => conv_std_logic_vector(115, 8),
37070 => conv_std_logic_vector(115, 8),
37071 => conv_std_logic_vector(116, 8),
37072 => conv_std_logic_vector(117, 8),
37073 => conv_std_logic_vector(117, 8),
37074 => conv_std_logic_vector(118, 8),
37075 => conv_std_logic_vector(118, 8),
37076 => conv_std_logic_vector(119, 8),
37077 => conv_std_logic_vector(119, 8),
37078 => conv_std_logic_vector(120, 8),
37079 => conv_std_logic_vector(120, 8),
37080 => conv_std_logic_vector(121, 8),
37081 => conv_std_logic_vector(122, 8),
37082 => conv_std_logic_vector(122, 8),
37083 => conv_std_logic_vector(123, 8),
37084 => conv_std_logic_vector(123, 8),
37085 => conv_std_logic_vector(124, 8),
37086 => conv_std_logic_vector(124, 8),
37087 => conv_std_logic_vector(125, 8),
37088 => conv_std_logic_vector(126, 8),
37089 => conv_std_logic_vector(126, 8),
37090 => conv_std_logic_vector(127, 8),
37091 => conv_std_logic_vector(127, 8),
37092 => conv_std_logic_vector(128, 8),
37093 => conv_std_logic_vector(128, 8),
37094 => conv_std_logic_vector(129, 8),
37095 => conv_std_logic_vector(129, 8),
37096 => conv_std_logic_vector(130, 8),
37097 => conv_std_logic_vector(131, 8),
37098 => conv_std_logic_vector(131, 8),
37099 => conv_std_logic_vector(132, 8),
37100 => conv_std_logic_vector(132, 8),
37101 => conv_std_logic_vector(133, 8),
37102 => conv_std_logic_vector(133, 8),
37103 => conv_std_logic_vector(134, 8),
37104 => conv_std_logic_vector(135, 8),
37105 => conv_std_logic_vector(135, 8),
37106 => conv_std_logic_vector(136, 8),
37107 => conv_std_logic_vector(136, 8),
37108 => conv_std_logic_vector(137, 8),
37109 => conv_std_logic_vector(137, 8),
37110 => conv_std_logic_vector(138, 8),
37111 => conv_std_logic_vector(138, 8),
37112 => conv_std_logic_vector(139, 8),
37113 => conv_std_logic_vector(140, 8),
37114 => conv_std_logic_vector(140, 8),
37115 => conv_std_logic_vector(141, 8),
37116 => conv_std_logic_vector(141, 8),
37117 => conv_std_logic_vector(142, 8),
37118 => conv_std_logic_vector(142, 8),
37119 => conv_std_logic_vector(143, 8),
37120 => conv_std_logic_vector(0, 8),
37121 => conv_std_logic_vector(0, 8),
37122 => conv_std_logic_vector(1, 8),
37123 => conv_std_logic_vector(1, 8),
37124 => conv_std_logic_vector(2, 8),
37125 => conv_std_logic_vector(2, 8),
37126 => conv_std_logic_vector(3, 8),
37127 => conv_std_logic_vector(3, 8),
37128 => conv_std_logic_vector(4, 8),
37129 => conv_std_logic_vector(5, 8),
37130 => conv_std_logic_vector(5, 8),
37131 => conv_std_logic_vector(6, 8),
37132 => conv_std_logic_vector(6, 8),
37133 => conv_std_logic_vector(7, 8),
37134 => conv_std_logic_vector(7, 8),
37135 => conv_std_logic_vector(8, 8),
37136 => conv_std_logic_vector(9, 8),
37137 => conv_std_logic_vector(9, 8),
37138 => conv_std_logic_vector(10, 8),
37139 => conv_std_logic_vector(10, 8),
37140 => conv_std_logic_vector(11, 8),
37141 => conv_std_logic_vector(11, 8),
37142 => conv_std_logic_vector(12, 8),
37143 => conv_std_logic_vector(13, 8),
37144 => conv_std_logic_vector(13, 8),
37145 => conv_std_logic_vector(14, 8),
37146 => conv_std_logic_vector(14, 8),
37147 => conv_std_logic_vector(15, 8),
37148 => conv_std_logic_vector(15, 8),
37149 => conv_std_logic_vector(16, 8),
37150 => conv_std_logic_vector(16, 8),
37151 => conv_std_logic_vector(17, 8),
37152 => conv_std_logic_vector(18, 8),
37153 => conv_std_logic_vector(18, 8),
37154 => conv_std_logic_vector(19, 8),
37155 => conv_std_logic_vector(19, 8),
37156 => conv_std_logic_vector(20, 8),
37157 => conv_std_logic_vector(20, 8),
37158 => conv_std_logic_vector(21, 8),
37159 => conv_std_logic_vector(22, 8),
37160 => conv_std_logic_vector(22, 8),
37161 => conv_std_logic_vector(23, 8),
37162 => conv_std_logic_vector(23, 8),
37163 => conv_std_logic_vector(24, 8),
37164 => conv_std_logic_vector(24, 8),
37165 => conv_std_logic_vector(25, 8),
37166 => conv_std_logic_vector(26, 8),
37167 => conv_std_logic_vector(26, 8),
37168 => conv_std_logic_vector(27, 8),
37169 => conv_std_logic_vector(27, 8),
37170 => conv_std_logic_vector(28, 8),
37171 => conv_std_logic_vector(28, 8),
37172 => conv_std_logic_vector(29, 8),
37173 => conv_std_logic_vector(30, 8),
37174 => conv_std_logic_vector(30, 8),
37175 => conv_std_logic_vector(31, 8),
37176 => conv_std_logic_vector(31, 8),
37177 => conv_std_logic_vector(32, 8),
37178 => conv_std_logic_vector(32, 8),
37179 => conv_std_logic_vector(33, 8),
37180 => conv_std_logic_vector(33, 8),
37181 => conv_std_logic_vector(34, 8),
37182 => conv_std_logic_vector(35, 8),
37183 => conv_std_logic_vector(35, 8),
37184 => conv_std_logic_vector(36, 8),
37185 => conv_std_logic_vector(36, 8),
37186 => conv_std_logic_vector(37, 8),
37187 => conv_std_logic_vector(37, 8),
37188 => conv_std_logic_vector(38, 8),
37189 => conv_std_logic_vector(39, 8),
37190 => conv_std_logic_vector(39, 8),
37191 => conv_std_logic_vector(40, 8),
37192 => conv_std_logic_vector(40, 8),
37193 => conv_std_logic_vector(41, 8),
37194 => conv_std_logic_vector(41, 8),
37195 => conv_std_logic_vector(42, 8),
37196 => conv_std_logic_vector(43, 8),
37197 => conv_std_logic_vector(43, 8),
37198 => conv_std_logic_vector(44, 8),
37199 => conv_std_logic_vector(44, 8),
37200 => conv_std_logic_vector(45, 8),
37201 => conv_std_logic_vector(45, 8),
37202 => conv_std_logic_vector(46, 8),
37203 => conv_std_logic_vector(47, 8),
37204 => conv_std_logic_vector(47, 8),
37205 => conv_std_logic_vector(48, 8),
37206 => conv_std_logic_vector(48, 8),
37207 => conv_std_logic_vector(49, 8),
37208 => conv_std_logic_vector(49, 8),
37209 => conv_std_logic_vector(50, 8),
37210 => conv_std_logic_vector(50, 8),
37211 => conv_std_logic_vector(51, 8),
37212 => conv_std_logic_vector(52, 8),
37213 => conv_std_logic_vector(52, 8),
37214 => conv_std_logic_vector(53, 8),
37215 => conv_std_logic_vector(53, 8),
37216 => conv_std_logic_vector(54, 8),
37217 => conv_std_logic_vector(54, 8),
37218 => conv_std_logic_vector(55, 8),
37219 => conv_std_logic_vector(56, 8),
37220 => conv_std_logic_vector(56, 8),
37221 => conv_std_logic_vector(57, 8),
37222 => conv_std_logic_vector(57, 8),
37223 => conv_std_logic_vector(58, 8),
37224 => conv_std_logic_vector(58, 8),
37225 => conv_std_logic_vector(59, 8),
37226 => conv_std_logic_vector(60, 8),
37227 => conv_std_logic_vector(60, 8),
37228 => conv_std_logic_vector(61, 8),
37229 => conv_std_logic_vector(61, 8),
37230 => conv_std_logic_vector(62, 8),
37231 => conv_std_logic_vector(62, 8),
37232 => conv_std_logic_vector(63, 8),
37233 => conv_std_logic_vector(64, 8),
37234 => conv_std_logic_vector(64, 8),
37235 => conv_std_logic_vector(65, 8),
37236 => conv_std_logic_vector(65, 8),
37237 => conv_std_logic_vector(66, 8),
37238 => conv_std_logic_vector(66, 8),
37239 => conv_std_logic_vector(67, 8),
37240 => conv_std_logic_vector(67, 8),
37241 => conv_std_logic_vector(68, 8),
37242 => conv_std_logic_vector(69, 8),
37243 => conv_std_logic_vector(69, 8),
37244 => conv_std_logic_vector(70, 8),
37245 => conv_std_logic_vector(70, 8),
37246 => conv_std_logic_vector(71, 8),
37247 => conv_std_logic_vector(71, 8),
37248 => conv_std_logic_vector(72, 8),
37249 => conv_std_logic_vector(73, 8),
37250 => conv_std_logic_vector(73, 8),
37251 => conv_std_logic_vector(74, 8),
37252 => conv_std_logic_vector(74, 8),
37253 => conv_std_logic_vector(75, 8),
37254 => conv_std_logic_vector(75, 8),
37255 => conv_std_logic_vector(76, 8),
37256 => conv_std_logic_vector(77, 8),
37257 => conv_std_logic_vector(77, 8),
37258 => conv_std_logic_vector(78, 8),
37259 => conv_std_logic_vector(78, 8),
37260 => conv_std_logic_vector(79, 8),
37261 => conv_std_logic_vector(79, 8),
37262 => conv_std_logic_vector(80, 8),
37263 => conv_std_logic_vector(80, 8),
37264 => conv_std_logic_vector(81, 8),
37265 => conv_std_logic_vector(82, 8),
37266 => conv_std_logic_vector(82, 8),
37267 => conv_std_logic_vector(83, 8),
37268 => conv_std_logic_vector(83, 8),
37269 => conv_std_logic_vector(84, 8),
37270 => conv_std_logic_vector(84, 8),
37271 => conv_std_logic_vector(85, 8),
37272 => conv_std_logic_vector(86, 8),
37273 => conv_std_logic_vector(86, 8),
37274 => conv_std_logic_vector(87, 8),
37275 => conv_std_logic_vector(87, 8),
37276 => conv_std_logic_vector(88, 8),
37277 => conv_std_logic_vector(88, 8),
37278 => conv_std_logic_vector(89, 8),
37279 => conv_std_logic_vector(90, 8),
37280 => conv_std_logic_vector(90, 8),
37281 => conv_std_logic_vector(91, 8),
37282 => conv_std_logic_vector(91, 8),
37283 => conv_std_logic_vector(92, 8),
37284 => conv_std_logic_vector(92, 8),
37285 => conv_std_logic_vector(93, 8),
37286 => conv_std_logic_vector(94, 8),
37287 => conv_std_logic_vector(94, 8),
37288 => conv_std_logic_vector(95, 8),
37289 => conv_std_logic_vector(95, 8),
37290 => conv_std_logic_vector(96, 8),
37291 => conv_std_logic_vector(96, 8),
37292 => conv_std_logic_vector(97, 8),
37293 => conv_std_logic_vector(97, 8),
37294 => conv_std_logic_vector(98, 8),
37295 => conv_std_logic_vector(99, 8),
37296 => conv_std_logic_vector(99, 8),
37297 => conv_std_logic_vector(100, 8),
37298 => conv_std_logic_vector(100, 8),
37299 => conv_std_logic_vector(101, 8),
37300 => conv_std_logic_vector(101, 8),
37301 => conv_std_logic_vector(102, 8),
37302 => conv_std_logic_vector(103, 8),
37303 => conv_std_logic_vector(103, 8),
37304 => conv_std_logic_vector(104, 8),
37305 => conv_std_logic_vector(104, 8),
37306 => conv_std_logic_vector(105, 8),
37307 => conv_std_logic_vector(105, 8),
37308 => conv_std_logic_vector(106, 8),
37309 => conv_std_logic_vector(107, 8),
37310 => conv_std_logic_vector(107, 8),
37311 => conv_std_logic_vector(108, 8),
37312 => conv_std_logic_vector(108, 8),
37313 => conv_std_logic_vector(109, 8),
37314 => conv_std_logic_vector(109, 8),
37315 => conv_std_logic_vector(110, 8),
37316 => conv_std_logic_vector(111, 8),
37317 => conv_std_logic_vector(111, 8),
37318 => conv_std_logic_vector(112, 8),
37319 => conv_std_logic_vector(112, 8),
37320 => conv_std_logic_vector(113, 8),
37321 => conv_std_logic_vector(113, 8),
37322 => conv_std_logic_vector(114, 8),
37323 => conv_std_logic_vector(114, 8),
37324 => conv_std_logic_vector(115, 8),
37325 => conv_std_logic_vector(116, 8),
37326 => conv_std_logic_vector(116, 8),
37327 => conv_std_logic_vector(117, 8),
37328 => conv_std_logic_vector(117, 8),
37329 => conv_std_logic_vector(118, 8),
37330 => conv_std_logic_vector(118, 8),
37331 => conv_std_logic_vector(119, 8),
37332 => conv_std_logic_vector(120, 8),
37333 => conv_std_logic_vector(120, 8),
37334 => conv_std_logic_vector(121, 8),
37335 => conv_std_logic_vector(121, 8),
37336 => conv_std_logic_vector(122, 8),
37337 => conv_std_logic_vector(122, 8),
37338 => conv_std_logic_vector(123, 8),
37339 => conv_std_logic_vector(124, 8),
37340 => conv_std_logic_vector(124, 8),
37341 => conv_std_logic_vector(125, 8),
37342 => conv_std_logic_vector(125, 8),
37343 => conv_std_logic_vector(126, 8),
37344 => conv_std_logic_vector(126, 8),
37345 => conv_std_logic_vector(127, 8),
37346 => conv_std_logic_vector(128, 8),
37347 => conv_std_logic_vector(128, 8),
37348 => conv_std_logic_vector(129, 8),
37349 => conv_std_logic_vector(129, 8),
37350 => conv_std_logic_vector(130, 8),
37351 => conv_std_logic_vector(130, 8),
37352 => conv_std_logic_vector(131, 8),
37353 => conv_std_logic_vector(131, 8),
37354 => conv_std_logic_vector(132, 8),
37355 => conv_std_logic_vector(133, 8),
37356 => conv_std_logic_vector(133, 8),
37357 => conv_std_logic_vector(134, 8),
37358 => conv_std_logic_vector(134, 8),
37359 => conv_std_logic_vector(135, 8),
37360 => conv_std_logic_vector(135, 8),
37361 => conv_std_logic_vector(136, 8),
37362 => conv_std_logic_vector(137, 8),
37363 => conv_std_logic_vector(137, 8),
37364 => conv_std_logic_vector(138, 8),
37365 => conv_std_logic_vector(138, 8),
37366 => conv_std_logic_vector(139, 8),
37367 => conv_std_logic_vector(139, 8),
37368 => conv_std_logic_vector(140, 8),
37369 => conv_std_logic_vector(141, 8),
37370 => conv_std_logic_vector(141, 8),
37371 => conv_std_logic_vector(142, 8),
37372 => conv_std_logic_vector(142, 8),
37373 => conv_std_logic_vector(143, 8),
37374 => conv_std_logic_vector(143, 8),
37375 => conv_std_logic_vector(144, 8),
37376 => conv_std_logic_vector(0, 8),
37377 => conv_std_logic_vector(0, 8),
37378 => conv_std_logic_vector(1, 8),
37379 => conv_std_logic_vector(1, 8),
37380 => conv_std_logic_vector(2, 8),
37381 => conv_std_logic_vector(2, 8),
37382 => conv_std_logic_vector(3, 8),
37383 => conv_std_logic_vector(3, 8),
37384 => conv_std_logic_vector(4, 8),
37385 => conv_std_logic_vector(5, 8),
37386 => conv_std_logic_vector(5, 8),
37387 => conv_std_logic_vector(6, 8),
37388 => conv_std_logic_vector(6, 8),
37389 => conv_std_logic_vector(7, 8),
37390 => conv_std_logic_vector(7, 8),
37391 => conv_std_logic_vector(8, 8),
37392 => conv_std_logic_vector(9, 8),
37393 => conv_std_logic_vector(9, 8),
37394 => conv_std_logic_vector(10, 8),
37395 => conv_std_logic_vector(10, 8),
37396 => conv_std_logic_vector(11, 8),
37397 => conv_std_logic_vector(11, 8),
37398 => conv_std_logic_vector(12, 8),
37399 => conv_std_logic_vector(13, 8),
37400 => conv_std_logic_vector(13, 8),
37401 => conv_std_logic_vector(14, 8),
37402 => conv_std_logic_vector(14, 8),
37403 => conv_std_logic_vector(15, 8),
37404 => conv_std_logic_vector(15, 8),
37405 => conv_std_logic_vector(16, 8),
37406 => conv_std_logic_vector(17, 8),
37407 => conv_std_logic_vector(17, 8),
37408 => conv_std_logic_vector(18, 8),
37409 => conv_std_logic_vector(18, 8),
37410 => conv_std_logic_vector(19, 8),
37411 => conv_std_logic_vector(19, 8),
37412 => conv_std_logic_vector(20, 8),
37413 => conv_std_logic_vector(21, 8),
37414 => conv_std_logic_vector(21, 8),
37415 => conv_std_logic_vector(22, 8),
37416 => conv_std_logic_vector(22, 8),
37417 => conv_std_logic_vector(23, 8),
37418 => conv_std_logic_vector(23, 8),
37419 => conv_std_logic_vector(24, 8),
37420 => conv_std_logic_vector(25, 8),
37421 => conv_std_logic_vector(25, 8),
37422 => conv_std_logic_vector(26, 8),
37423 => conv_std_logic_vector(26, 8),
37424 => conv_std_logic_vector(27, 8),
37425 => conv_std_logic_vector(27, 8),
37426 => conv_std_logic_vector(28, 8),
37427 => conv_std_logic_vector(29, 8),
37428 => conv_std_logic_vector(29, 8),
37429 => conv_std_logic_vector(30, 8),
37430 => conv_std_logic_vector(30, 8),
37431 => conv_std_logic_vector(31, 8),
37432 => conv_std_logic_vector(31, 8),
37433 => conv_std_logic_vector(32, 8),
37434 => conv_std_logic_vector(33, 8),
37435 => conv_std_logic_vector(33, 8),
37436 => conv_std_logic_vector(34, 8),
37437 => conv_std_logic_vector(34, 8),
37438 => conv_std_logic_vector(35, 8),
37439 => conv_std_logic_vector(35, 8),
37440 => conv_std_logic_vector(36, 8),
37441 => conv_std_logic_vector(37, 8),
37442 => conv_std_logic_vector(37, 8),
37443 => conv_std_logic_vector(38, 8),
37444 => conv_std_logic_vector(38, 8),
37445 => conv_std_logic_vector(39, 8),
37446 => conv_std_logic_vector(39, 8),
37447 => conv_std_logic_vector(40, 8),
37448 => conv_std_logic_vector(41, 8),
37449 => conv_std_logic_vector(41, 8),
37450 => conv_std_logic_vector(42, 8),
37451 => conv_std_logic_vector(42, 8),
37452 => conv_std_logic_vector(43, 8),
37453 => conv_std_logic_vector(43, 8),
37454 => conv_std_logic_vector(44, 8),
37455 => conv_std_logic_vector(45, 8),
37456 => conv_std_logic_vector(45, 8),
37457 => conv_std_logic_vector(46, 8),
37458 => conv_std_logic_vector(46, 8),
37459 => conv_std_logic_vector(47, 8),
37460 => conv_std_logic_vector(47, 8),
37461 => conv_std_logic_vector(48, 8),
37462 => conv_std_logic_vector(49, 8),
37463 => conv_std_logic_vector(49, 8),
37464 => conv_std_logic_vector(50, 8),
37465 => conv_std_logic_vector(50, 8),
37466 => conv_std_logic_vector(51, 8),
37467 => conv_std_logic_vector(51, 8),
37468 => conv_std_logic_vector(52, 8),
37469 => conv_std_logic_vector(53, 8),
37470 => conv_std_logic_vector(53, 8),
37471 => conv_std_logic_vector(54, 8),
37472 => conv_std_logic_vector(54, 8),
37473 => conv_std_logic_vector(55, 8),
37474 => conv_std_logic_vector(55, 8),
37475 => conv_std_logic_vector(56, 8),
37476 => conv_std_logic_vector(57, 8),
37477 => conv_std_logic_vector(57, 8),
37478 => conv_std_logic_vector(58, 8),
37479 => conv_std_logic_vector(58, 8),
37480 => conv_std_logic_vector(59, 8),
37481 => conv_std_logic_vector(59, 8),
37482 => conv_std_logic_vector(60, 8),
37483 => conv_std_logic_vector(61, 8),
37484 => conv_std_logic_vector(61, 8),
37485 => conv_std_logic_vector(62, 8),
37486 => conv_std_logic_vector(62, 8),
37487 => conv_std_logic_vector(63, 8),
37488 => conv_std_logic_vector(63, 8),
37489 => conv_std_logic_vector(64, 8),
37490 => conv_std_logic_vector(65, 8),
37491 => conv_std_logic_vector(65, 8),
37492 => conv_std_logic_vector(66, 8),
37493 => conv_std_logic_vector(66, 8),
37494 => conv_std_logic_vector(67, 8),
37495 => conv_std_logic_vector(67, 8),
37496 => conv_std_logic_vector(68, 8),
37497 => conv_std_logic_vector(69, 8),
37498 => conv_std_logic_vector(69, 8),
37499 => conv_std_logic_vector(70, 8),
37500 => conv_std_logic_vector(70, 8),
37501 => conv_std_logic_vector(71, 8),
37502 => conv_std_logic_vector(71, 8),
37503 => conv_std_logic_vector(72, 8),
37504 => conv_std_logic_vector(73, 8),
37505 => conv_std_logic_vector(73, 8),
37506 => conv_std_logic_vector(74, 8),
37507 => conv_std_logic_vector(74, 8),
37508 => conv_std_logic_vector(75, 8),
37509 => conv_std_logic_vector(75, 8),
37510 => conv_std_logic_vector(76, 8),
37511 => conv_std_logic_vector(76, 8),
37512 => conv_std_logic_vector(77, 8),
37513 => conv_std_logic_vector(78, 8),
37514 => conv_std_logic_vector(78, 8),
37515 => conv_std_logic_vector(79, 8),
37516 => conv_std_logic_vector(79, 8),
37517 => conv_std_logic_vector(80, 8),
37518 => conv_std_logic_vector(80, 8),
37519 => conv_std_logic_vector(81, 8),
37520 => conv_std_logic_vector(82, 8),
37521 => conv_std_logic_vector(82, 8),
37522 => conv_std_logic_vector(83, 8),
37523 => conv_std_logic_vector(83, 8),
37524 => conv_std_logic_vector(84, 8),
37525 => conv_std_logic_vector(84, 8),
37526 => conv_std_logic_vector(85, 8),
37527 => conv_std_logic_vector(86, 8),
37528 => conv_std_logic_vector(86, 8),
37529 => conv_std_logic_vector(87, 8),
37530 => conv_std_logic_vector(87, 8),
37531 => conv_std_logic_vector(88, 8),
37532 => conv_std_logic_vector(88, 8),
37533 => conv_std_logic_vector(89, 8),
37534 => conv_std_logic_vector(90, 8),
37535 => conv_std_logic_vector(90, 8),
37536 => conv_std_logic_vector(91, 8),
37537 => conv_std_logic_vector(91, 8),
37538 => conv_std_logic_vector(92, 8),
37539 => conv_std_logic_vector(92, 8),
37540 => conv_std_logic_vector(93, 8),
37541 => conv_std_logic_vector(94, 8),
37542 => conv_std_logic_vector(94, 8),
37543 => conv_std_logic_vector(95, 8),
37544 => conv_std_logic_vector(95, 8),
37545 => conv_std_logic_vector(96, 8),
37546 => conv_std_logic_vector(96, 8),
37547 => conv_std_logic_vector(97, 8),
37548 => conv_std_logic_vector(98, 8),
37549 => conv_std_logic_vector(98, 8),
37550 => conv_std_logic_vector(99, 8),
37551 => conv_std_logic_vector(99, 8),
37552 => conv_std_logic_vector(100, 8),
37553 => conv_std_logic_vector(100, 8),
37554 => conv_std_logic_vector(101, 8),
37555 => conv_std_logic_vector(102, 8),
37556 => conv_std_logic_vector(102, 8),
37557 => conv_std_logic_vector(103, 8),
37558 => conv_std_logic_vector(103, 8),
37559 => conv_std_logic_vector(104, 8),
37560 => conv_std_logic_vector(104, 8),
37561 => conv_std_logic_vector(105, 8),
37562 => conv_std_logic_vector(106, 8),
37563 => conv_std_logic_vector(106, 8),
37564 => conv_std_logic_vector(107, 8),
37565 => conv_std_logic_vector(107, 8),
37566 => conv_std_logic_vector(108, 8),
37567 => conv_std_logic_vector(108, 8),
37568 => conv_std_logic_vector(109, 8),
37569 => conv_std_logic_vector(110, 8),
37570 => conv_std_logic_vector(110, 8),
37571 => conv_std_logic_vector(111, 8),
37572 => conv_std_logic_vector(111, 8),
37573 => conv_std_logic_vector(112, 8),
37574 => conv_std_logic_vector(112, 8),
37575 => conv_std_logic_vector(113, 8),
37576 => conv_std_logic_vector(114, 8),
37577 => conv_std_logic_vector(114, 8),
37578 => conv_std_logic_vector(115, 8),
37579 => conv_std_logic_vector(115, 8),
37580 => conv_std_logic_vector(116, 8),
37581 => conv_std_logic_vector(116, 8),
37582 => conv_std_logic_vector(117, 8),
37583 => conv_std_logic_vector(118, 8),
37584 => conv_std_logic_vector(118, 8),
37585 => conv_std_logic_vector(119, 8),
37586 => conv_std_logic_vector(119, 8),
37587 => conv_std_logic_vector(120, 8),
37588 => conv_std_logic_vector(120, 8),
37589 => conv_std_logic_vector(121, 8),
37590 => conv_std_logic_vector(122, 8),
37591 => conv_std_logic_vector(122, 8),
37592 => conv_std_logic_vector(123, 8),
37593 => conv_std_logic_vector(123, 8),
37594 => conv_std_logic_vector(124, 8),
37595 => conv_std_logic_vector(124, 8),
37596 => conv_std_logic_vector(125, 8),
37597 => conv_std_logic_vector(126, 8),
37598 => conv_std_logic_vector(126, 8),
37599 => conv_std_logic_vector(127, 8),
37600 => conv_std_logic_vector(127, 8),
37601 => conv_std_logic_vector(128, 8),
37602 => conv_std_logic_vector(128, 8),
37603 => conv_std_logic_vector(129, 8),
37604 => conv_std_logic_vector(130, 8),
37605 => conv_std_logic_vector(130, 8),
37606 => conv_std_logic_vector(131, 8),
37607 => conv_std_logic_vector(131, 8),
37608 => conv_std_logic_vector(132, 8),
37609 => conv_std_logic_vector(132, 8),
37610 => conv_std_logic_vector(133, 8),
37611 => conv_std_logic_vector(134, 8),
37612 => conv_std_logic_vector(134, 8),
37613 => conv_std_logic_vector(135, 8),
37614 => conv_std_logic_vector(135, 8),
37615 => conv_std_logic_vector(136, 8),
37616 => conv_std_logic_vector(136, 8),
37617 => conv_std_logic_vector(137, 8),
37618 => conv_std_logic_vector(138, 8),
37619 => conv_std_logic_vector(138, 8),
37620 => conv_std_logic_vector(139, 8),
37621 => conv_std_logic_vector(139, 8),
37622 => conv_std_logic_vector(140, 8),
37623 => conv_std_logic_vector(140, 8),
37624 => conv_std_logic_vector(141, 8),
37625 => conv_std_logic_vector(142, 8),
37626 => conv_std_logic_vector(142, 8),
37627 => conv_std_logic_vector(143, 8),
37628 => conv_std_logic_vector(143, 8),
37629 => conv_std_logic_vector(144, 8),
37630 => conv_std_logic_vector(144, 8),
37631 => conv_std_logic_vector(145, 8),
37632 => conv_std_logic_vector(0, 8),
37633 => conv_std_logic_vector(0, 8),
37634 => conv_std_logic_vector(1, 8),
37635 => conv_std_logic_vector(1, 8),
37636 => conv_std_logic_vector(2, 8),
37637 => conv_std_logic_vector(2, 8),
37638 => conv_std_logic_vector(3, 8),
37639 => conv_std_logic_vector(4, 8),
37640 => conv_std_logic_vector(4, 8),
37641 => conv_std_logic_vector(5, 8),
37642 => conv_std_logic_vector(5, 8),
37643 => conv_std_logic_vector(6, 8),
37644 => conv_std_logic_vector(6, 8),
37645 => conv_std_logic_vector(7, 8),
37646 => conv_std_logic_vector(8, 8),
37647 => conv_std_logic_vector(8, 8),
37648 => conv_std_logic_vector(9, 8),
37649 => conv_std_logic_vector(9, 8),
37650 => conv_std_logic_vector(10, 8),
37651 => conv_std_logic_vector(10, 8),
37652 => conv_std_logic_vector(11, 8),
37653 => conv_std_logic_vector(12, 8),
37654 => conv_std_logic_vector(12, 8),
37655 => conv_std_logic_vector(13, 8),
37656 => conv_std_logic_vector(13, 8),
37657 => conv_std_logic_vector(14, 8),
37658 => conv_std_logic_vector(14, 8),
37659 => conv_std_logic_vector(15, 8),
37660 => conv_std_logic_vector(16, 8),
37661 => conv_std_logic_vector(16, 8),
37662 => conv_std_logic_vector(17, 8),
37663 => conv_std_logic_vector(17, 8),
37664 => conv_std_logic_vector(18, 8),
37665 => conv_std_logic_vector(18, 8),
37666 => conv_std_logic_vector(19, 8),
37667 => conv_std_logic_vector(20, 8),
37668 => conv_std_logic_vector(20, 8),
37669 => conv_std_logic_vector(21, 8),
37670 => conv_std_logic_vector(21, 8),
37671 => conv_std_logic_vector(22, 8),
37672 => conv_std_logic_vector(22, 8),
37673 => conv_std_logic_vector(23, 8),
37674 => conv_std_logic_vector(24, 8),
37675 => conv_std_logic_vector(24, 8),
37676 => conv_std_logic_vector(25, 8),
37677 => conv_std_logic_vector(25, 8),
37678 => conv_std_logic_vector(26, 8),
37679 => conv_std_logic_vector(26, 8),
37680 => conv_std_logic_vector(27, 8),
37681 => conv_std_logic_vector(28, 8),
37682 => conv_std_logic_vector(28, 8),
37683 => conv_std_logic_vector(29, 8),
37684 => conv_std_logic_vector(29, 8),
37685 => conv_std_logic_vector(30, 8),
37686 => conv_std_logic_vector(31, 8),
37687 => conv_std_logic_vector(31, 8),
37688 => conv_std_logic_vector(32, 8),
37689 => conv_std_logic_vector(32, 8),
37690 => conv_std_logic_vector(33, 8),
37691 => conv_std_logic_vector(33, 8),
37692 => conv_std_logic_vector(34, 8),
37693 => conv_std_logic_vector(35, 8),
37694 => conv_std_logic_vector(35, 8),
37695 => conv_std_logic_vector(36, 8),
37696 => conv_std_logic_vector(36, 8),
37697 => conv_std_logic_vector(37, 8),
37698 => conv_std_logic_vector(37, 8),
37699 => conv_std_logic_vector(38, 8),
37700 => conv_std_logic_vector(39, 8),
37701 => conv_std_logic_vector(39, 8),
37702 => conv_std_logic_vector(40, 8),
37703 => conv_std_logic_vector(40, 8),
37704 => conv_std_logic_vector(41, 8),
37705 => conv_std_logic_vector(41, 8),
37706 => conv_std_logic_vector(42, 8),
37707 => conv_std_logic_vector(43, 8),
37708 => conv_std_logic_vector(43, 8),
37709 => conv_std_logic_vector(44, 8),
37710 => conv_std_logic_vector(44, 8),
37711 => conv_std_logic_vector(45, 8),
37712 => conv_std_logic_vector(45, 8),
37713 => conv_std_logic_vector(46, 8),
37714 => conv_std_logic_vector(47, 8),
37715 => conv_std_logic_vector(47, 8),
37716 => conv_std_logic_vector(48, 8),
37717 => conv_std_logic_vector(48, 8),
37718 => conv_std_logic_vector(49, 8),
37719 => conv_std_logic_vector(49, 8),
37720 => conv_std_logic_vector(50, 8),
37721 => conv_std_logic_vector(51, 8),
37722 => conv_std_logic_vector(51, 8),
37723 => conv_std_logic_vector(52, 8),
37724 => conv_std_logic_vector(52, 8),
37725 => conv_std_logic_vector(53, 8),
37726 => conv_std_logic_vector(53, 8),
37727 => conv_std_logic_vector(54, 8),
37728 => conv_std_logic_vector(55, 8),
37729 => conv_std_logic_vector(55, 8),
37730 => conv_std_logic_vector(56, 8),
37731 => conv_std_logic_vector(56, 8),
37732 => conv_std_logic_vector(57, 8),
37733 => conv_std_logic_vector(57, 8),
37734 => conv_std_logic_vector(58, 8),
37735 => conv_std_logic_vector(59, 8),
37736 => conv_std_logic_vector(59, 8),
37737 => conv_std_logic_vector(60, 8),
37738 => conv_std_logic_vector(60, 8),
37739 => conv_std_logic_vector(61, 8),
37740 => conv_std_logic_vector(62, 8),
37741 => conv_std_logic_vector(62, 8),
37742 => conv_std_logic_vector(63, 8),
37743 => conv_std_logic_vector(63, 8),
37744 => conv_std_logic_vector(64, 8),
37745 => conv_std_logic_vector(64, 8),
37746 => conv_std_logic_vector(65, 8),
37747 => conv_std_logic_vector(66, 8),
37748 => conv_std_logic_vector(66, 8),
37749 => conv_std_logic_vector(67, 8),
37750 => conv_std_logic_vector(67, 8),
37751 => conv_std_logic_vector(68, 8),
37752 => conv_std_logic_vector(68, 8),
37753 => conv_std_logic_vector(69, 8),
37754 => conv_std_logic_vector(70, 8),
37755 => conv_std_logic_vector(70, 8),
37756 => conv_std_logic_vector(71, 8),
37757 => conv_std_logic_vector(71, 8),
37758 => conv_std_logic_vector(72, 8),
37759 => conv_std_logic_vector(72, 8),
37760 => conv_std_logic_vector(73, 8),
37761 => conv_std_logic_vector(74, 8),
37762 => conv_std_logic_vector(74, 8),
37763 => conv_std_logic_vector(75, 8),
37764 => conv_std_logic_vector(75, 8),
37765 => conv_std_logic_vector(76, 8),
37766 => conv_std_logic_vector(76, 8),
37767 => conv_std_logic_vector(77, 8),
37768 => conv_std_logic_vector(78, 8),
37769 => conv_std_logic_vector(78, 8),
37770 => conv_std_logic_vector(79, 8),
37771 => conv_std_logic_vector(79, 8),
37772 => conv_std_logic_vector(80, 8),
37773 => conv_std_logic_vector(80, 8),
37774 => conv_std_logic_vector(81, 8),
37775 => conv_std_logic_vector(82, 8),
37776 => conv_std_logic_vector(82, 8),
37777 => conv_std_logic_vector(83, 8),
37778 => conv_std_logic_vector(83, 8),
37779 => conv_std_logic_vector(84, 8),
37780 => conv_std_logic_vector(84, 8),
37781 => conv_std_logic_vector(85, 8),
37782 => conv_std_logic_vector(86, 8),
37783 => conv_std_logic_vector(86, 8),
37784 => conv_std_logic_vector(87, 8),
37785 => conv_std_logic_vector(87, 8),
37786 => conv_std_logic_vector(88, 8),
37787 => conv_std_logic_vector(89, 8),
37788 => conv_std_logic_vector(89, 8),
37789 => conv_std_logic_vector(90, 8),
37790 => conv_std_logic_vector(90, 8),
37791 => conv_std_logic_vector(91, 8),
37792 => conv_std_logic_vector(91, 8),
37793 => conv_std_logic_vector(92, 8),
37794 => conv_std_logic_vector(93, 8),
37795 => conv_std_logic_vector(93, 8),
37796 => conv_std_logic_vector(94, 8),
37797 => conv_std_logic_vector(94, 8),
37798 => conv_std_logic_vector(95, 8),
37799 => conv_std_logic_vector(95, 8),
37800 => conv_std_logic_vector(96, 8),
37801 => conv_std_logic_vector(97, 8),
37802 => conv_std_logic_vector(97, 8),
37803 => conv_std_logic_vector(98, 8),
37804 => conv_std_logic_vector(98, 8),
37805 => conv_std_logic_vector(99, 8),
37806 => conv_std_logic_vector(99, 8),
37807 => conv_std_logic_vector(100, 8),
37808 => conv_std_logic_vector(101, 8),
37809 => conv_std_logic_vector(101, 8),
37810 => conv_std_logic_vector(102, 8),
37811 => conv_std_logic_vector(102, 8),
37812 => conv_std_logic_vector(103, 8),
37813 => conv_std_logic_vector(103, 8),
37814 => conv_std_logic_vector(104, 8),
37815 => conv_std_logic_vector(105, 8),
37816 => conv_std_logic_vector(105, 8),
37817 => conv_std_logic_vector(106, 8),
37818 => conv_std_logic_vector(106, 8),
37819 => conv_std_logic_vector(107, 8),
37820 => conv_std_logic_vector(107, 8),
37821 => conv_std_logic_vector(108, 8),
37822 => conv_std_logic_vector(109, 8),
37823 => conv_std_logic_vector(109, 8),
37824 => conv_std_logic_vector(110, 8),
37825 => conv_std_logic_vector(110, 8),
37826 => conv_std_logic_vector(111, 8),
37827 => conv_std_logic_vector(111, 8),
37828 => conv_std_logic_vector(112, 8),
37829 => conv_std_logic_vector(113, 8),
37830 => conv_std_logic_vector(113, 8),
37831 => conv_std_logic_vector(114, 8),
37832 => conv_std_logic_vector(114, 8),
37833 => conv_std_logic_vector(115, 8),
37834 => conv_std_logic_vector(115, 8),
37835 => conv_std_logic_vector(116, 8),
37836 => conv_std_logic_vector(117, 8),
37837 => conv_std_logic_vector(117, 8),
37838 => conv_std_logic_vector(118, 8),
37839 => conv_std_logic_vector(118, 8),
37840 => conv_std_logic_vector(119, 8),
37841 => conv_std_logic_vector(120, 8),
37842 => conv_std_logic_vector(120, 8),
37843 => conv_std_logic_vector(121, 8),
37844 => conv_std_logic_vector(121, 8),
37845 => conv_std_logic_vector(122, 8),
37846 => conv_std_logic_vector(122, 8),
37847 => conv_std_logic_vector(123, 8),
37848 => conv_std_logic_vector(124, 8),
37849 => conv_std_logic_vector(124, 8),
37850 => conv_std_logic_vector(125, 8),
37851 => conv_std_logic_vector(125, 8),
37852 => conv_std_logic_vector(126, 8),
37853 => conv_std_logic_vector(126, 8),
37854 => conv_std_logic_vector(127, 8),
37855 => conv_std_logic_vector(128, 8),
37856 => conv_std_logic_vector(128, 8),
37857 => conv_std_logic_vector(129, 8),
37858 => conv_std_logic_vector(129, 8),
37859 => conv_std_logic_vector(130, 8),
37860 => conv_std_logic_vector(130, 8),
37861 => conv_std_logic_vector(131, 8),
37862 => conv_std_logic_vector(132, 8),
37863 => conv_std_logic_vector(132, 8),
37864 => conv_std_logic_vector(133, 8),
37865 => conv_std_logic_vector(133, 8),
37866 => conv_std_logic_vector(134, 8),
37867 => conv_std_logic_vector(134, 8),
37868 => conv_std_logic_vector(135, 8),
37869 => conv_std_logic_vector(136, 8),
37870 => conv_std_logic_vector(136, 8),
37871 => conv_std_logic_vector(137, 8),
37872 => conv_std_logic_vector(137, 8),
37873 => conv_std_logic_vector(138, 8),
37874 => conv_std_logic_vector(138, 8),
37875 => conv_std_logic_vector(139, 8),
37876 => conv_std_logic_vector(140, 8),
37877 => conv_std_logic_vector(140, 8),
37878 => conv_std_logic_vector(141, 8),
37879 => conv_std_logic_vector(141, 8),
37880 => conv_std_logic_vector(142, 8),
37881 => conv_std_logic_vector(142, 8),
37882 => conv_std_logic_vector(143, 8),
37883 => conv_std_logic_vector(144, 8),
37884 => conv_std_logic_vector(144, 8),
37885 => conv_std_logic_vector(145, 8),
37886 => conv_std_logic_vector(145, 8),
37887 => conv_std_logic_vector(146, 8),
37888 => conv_std_logic_vector(0, 8),
37889 => conv_std_logic_vector(0, 8),
37890 => conv_std_logic_vector(1, 8),
37891 => conv_std_logic_vector(1, 8),
37892 => conv_std_logic_vector(2, 8),
37893 => conv_std_logic_vector(2, 8),
37894 => conv_std_logic_vector(3, 8),
37895 => conv_std_logic_vector(4, 8),
37896 => conv_std_logic_vector(4, 8),
37897 => conv_std_logic_vector(5, 8),
37898 => conv_std_logic_vector(5, 8),
37899 => conv_std_logic_vector(6, 8),
37900 => conv_std_logic_vector(6, 8),
37901 => conv_std_logic_vector(7, 8),
37902 => conv_std_logic_vector(8, 8),
37903 => conv_std_logic_vector(8, 8),
37904 => conv_std_logic_vector(9, 8),
37905 => conv_std_logic_vector(9, 8),
37906 => conv_std_logic_vector(10, 8),
37907 => conv_std_logic_vector(10, 8),
37908 => conv_std_logic_vector(11, 8),
37909 => conv_std_logic_vector(12, 8),
37910 => conv_std_logic_vector(12, 8),
37911 => conv_std_logic_vector(13, 8),
37912 => conv_std_logic_vector(13, 8),
37913 => conv_std_logic_vector(14, 8),
37914 => conv_std_logic_vector(15, 8),
37915 => conv_std_logic_vector(15, 8),
37916 => conv_std_logic_vector(16, 8),
37917 => conv_std_logic_vector(16, 8),
37918 => conv_std_logic_vector(17, 8),
37919 => conv_std_logic_vector(17, 8),
37920 => conv_std_logic_vector(18, 8),
37921 => conv_std_logic_vector(19, 8),
37922 => conv_std_logic_vector(19, 8),
37923 => conv_std_logic_vector(20, 8),
37924 => conv_std_logic_vector(20, 8),
37925 => conv_std_logic_vector(21, 8),
37926 => conv_std_logic_vector(21, 8),
37927 => conv_std_logic_vector(22, 8),
37928 => conv_std_logic_vector(23, 8),
37929 => conv_std_logic_vector(23, 8),
37930 => conv_std_logic_vector(24, 8),
37931 => conv_std_logic_vector(24, 8),
37932 => conv_std_logic_vector(25, 8),
37933 => conv_std_logic_vector(26, 8),
37934 => conv_std_logic_vector(26, 8),
37935 => conv_std_logic_vector(27, 8),
37936 => conv_std_logic_vector(27, 8),
37937 => conv_std_logic_vector(28, 8),
37938 => conv_std_logic_vector(28, 8),
37939 => conv_std_logic_vector(29, 8),
37940 => conv_std_logic_vector(30, 8),
37941 => conv_std_logic_vector(30, 8),
37942 => conv_std_logic_vector(31, 8),
37943 => conv_std_logic_vector(31, 8),
37944 => conv_std_logic_vector(32, 8),
37945 => conv_std_logic_vector(32, 8),
37946 => conv_std_logic_vector(33, 8),
37947 => conv_std_logic_vector(34, 8),
37948 => conv_std_logic_vector(34, 8),
37949 => conv_std_logic_vector(35, 8),
37950 => conv_std_logic_vector(35, 8),
37951 => conv_std_logic_vector(36, 8),
37952 => conv_std_logic_vector(37, 8),
37953 => conv_std_logic_vector(37, 8),
37954 => conv_std_logic_vector(38, 8),
37955 => conv_std_logic_vector(38, 8),
37956 => conv_std_logic_vector(39, 8),
37957 => conv_std_logic_vector(39, 8),
37958 => conv_std_logic_vector(40, 8),
37959 => conv_std_logic_vector(41, 8),
37960 => conv_std_logic_vector(41, 8),
37961 => conv_std_logic_vector(42, 8),
37962 => conv_std_logic_vector(42, 8),
37963 => conv_std_logic_vector(43, 8),
37964 => conv_std_logic_vector(43, 8),
37965 => conv_std_logic_vector(44, 8),
37966 => conv_std_logic_vector(45, 8),
37967 => conv_std_logic_vector(45, 8),
37968 => conv_std_logic_vector(46, 8),
37969 => conv_std_logic_vector(46, 8),
37970 => conv_std_logic_vector(47, 8),
37971 => conv_std_logic_vector(47, 8),
37972 => conv_std_logic_vector(48, 8),
37973 => conv_std_logic_vector(49, 8),
37974 => conv_std_logic_vector(49, 8),
37975 => conv_std_logic_vector(50, 8),
37976 => conv_std_logic_vector(50, 8),
37977 => conv_std_logic_vector(51, 8),
37978 => conv_std_logic_vector(52, 8),
37979 => conv_std_logic_vector(52, 8),
37980 => conv_std_logic_vector(53, 8),
37981 => conv_std_logic_vector(53, 8),
37982 => conv_std_logic_vector(54, 8),
37983 => conv_std_logic_vector(54, 8),
37984 => conv_std_logic_vector(55, 8),
37985 => conv_std_logic_vector(56, 8),
37986 => conv_std_logic_vector(56, 8),
37987 => conv_std_logic_vector(57, 8),
37988 => conv_std_logic_vector(57, 8),
37989 => conv_std_logic_vector(58, 8),
37990 => conv_std_logic_vector(58, 8),
37991 => conv_std_logic_vector(59, 8),
37992 => conv_std_logic_vector(60, 8),
37993 => conv_std_logic_vector(60, 8),
37994 => conv_std_logic_vector(61, 8),
37995 => conv_std_logic_vector(61, 8),
37996 => conv_std_logic_vector(62, 8),
37997 => conv_std_logic_vector(63, 8),
37998 => conv_std_logic_vector(63, 8),
37999 => conv_std_logic_vector(64, 8),
38000 => conv_std_logic_vector(64, 8),
38001 => conv_std_logic_vector(65, 8),
38002 => conv_std_logic_vector(65, 8),
38003 => conv_std_logic_vector(66, 8),
38004 => conv_std_logic_vector(67, 8),
38005 => conv_std_logic_vector(67, 8),
38006 => conv_std_logic_vector(68, 8),
38007 => conv_std_logic_vector(68, 8),
38008 => conv_std_logic_vector(69, 8),
38009 => conv_std_logic_vector(69, 8),
38010 => conv_std_logic_vector(70, 8),
38011 => conv_std_logic_vector(71, 8),
38012 => conv_std_logic_vector(71, 8),
38013 => conv_std_logic_vector(72, 8),
38014 => conv_std_logic_vector(72, 8),
38015 => conv_std_logic_vector(73, 8),
38016 => conv_std_logic_vector(74, 8),
38017 => conv_std_logic_vector(74, 8),
38018 => conv_std_logic_vector(75, 8),
38019 => conv_std_logic_vector(75, 8),
38020 => conv_std_logic_vector(76, 8),
38021 => conv_std_logic_vector(76, 8),
38022 => conv_std_logic_vector(77, 8),
38023 => conv_std_logic_vector(78, 8),
38024 => conv_std_logic_vector(78, 8),
38025 => conv_std_logic_vector(79, 8),
38026 => conv_std_logic_vector(79, 8),
38027 => conv_std_logic_vector(80, 8),
38028 => conv_std_logic_vector(80, 8),
38029 => conv_std_logic_vector(81, 8),
38030 => conv_std_logic_vector(82, 8),
38031 => conv_std_logic_vector(82, 8),
38032 => conv_std_logic_vector(83, 8),
38033 => conv_std_logic_vector(83, 8),
38034 => conv_std_logic_vector(84, 8),
38035 => conv_std_logic_vector(84, 8),
38036 => conv_std_logic_vector(85, 8),
38037 => conv_std_logic_vector(86, 8),
38038 => conv_std_logic_vector(86, 8),
38039 => conv_std_logic_vector(87, 8),
38040 => conv_std_logic_vector(87, 8),
38041 => conv_std_logic_vector(88, 8),
38042 => conv_std_logic_vector(89, 8),
38043 => conv_std_logic_vector(89, 8),
38044 => conv_std_logic_vector(90, 8),
38045 => conv_std_logic_vector(90, 8),
38046 => conv_std_logic_vector(91, 8),
38047 => conv_std_logic_vector(91, 8),
38048 => conv_std_logic_vector(92, 8),
38049 => conv_std_logic_vector(93, 8),
38050 => conv_std_logic_vector(93, 8),
38051 => conv_std_logic_vector(94, 8),
38052 => conv_std_logic_vector(94, 8),
38053 => conv_std_logic_vector(95, 8),
38054 => conv_std_logic_vector(95, 8),
38055 => conv_std_logic_vector(96, 8),
38056 => conv_std_logic_vector(97, 8),
38057 => conv_std_logic_vector(97, 8),
38058 => conv_std_logic_vector(98, 8),
38059 => conv_std_logic_vector(98, 8),
38060 => conv_std_logic_vector(99, 8),
38061 => conv_std_logic_vector(100, 8),
38062 => conv_std_logic_vector(100, 8),
38063 => conv_std_logic_vector(101, 8),
38064 => conv_std_logic_vector(101, 8),
38065 => conv_std_logic_vector(102, 8),
38066 => conv_std_logic_vector(102, 8),
38067 => conv_std_logic_vector(103, 8),
38068 => conv_std_logic_vector(104, 8),
38069 => conv_std_logic_vector(104, 8),
38070 => conv_std_logic_vector(105, 8),
38071 => conv_std_logic_vector(105, 8),
38072 => conv_std_logic_vector(106, 8),
38073 => conv_std_logic_vector(106, 8),
38074 => conv_std_logic_vector(107, 8),
38075 => conv_std_logic_vector(108, 8),
38076 => conv_std_logic_vector(108, 8),
38077 => conv_std_logic_vector(109, 8),
38078 => conv_std_logic_vector(109, 8),
38079 => conv_std_logic_vector(110, 8),
38080 => conv_std_logic_vector(111, 8),
38081 => conv_std_logic_vector(111, 8),
38082 => conv_std_logic_vector(112, 8),
38083 => conv_std_logic_vector(112, 8),
38084 => conv_std_logic_vector(113, 8),
38085 => conv_std_logic_vector(113, 8),
38086 => conv_std_logic_vector(114, 8),
38087 => conv_std_logic_vector(115, 8),
38088 => conv_std_logic_vector(115, 8),
38089 => conv_std_logic_vector(116, 8),
38090 => conv_std_logic_vector(116, 8),
38091 => conv_std_logic_vector(117, 8),
38092 => conv_std_logic_vector(117, 8),
38093 => conv_std_logic_vector(118, 8),
38094 => conv_std_logic_vector(119, 8),
38095 => conv_std_logic_vector(119, 8),
38096 => conv_std_logic_vector(120, 8),
38097 => conv_std_logic_vector(120, 8),
38098 => conv_std_logic_vector(121, 8),
38099 => conv_std_logic_vector(121, 8),
38100 => conv_std_logic_vector(122, 8),
38101 => conv_std_logic_vector(123, 8),
38102 => conv_std_logic_vector(123, 8),
38103 => conv_std_logic_vector(124, 8),
38104 => conv_std_logic_vector(124, 8),
38105 => conv_std_logic_vector(125, 8),
38106 => conv_std_logic_vector(126, 8),
38107 => conv_std_logic_vector(126, 8),
38108 => conv_std_logic_vector(127, 8),
38109 => conv_std_logic_vector(127, 8),
38110 => conv_std_logic_vector(128, 8),
38111 => conv_std_logic_vector(128, 8),
38112 => conv_std_logic_vector(129, 8),
38113 => conv_std_logic_vector(130, 8),
38114 => conv_std_logic_vector(130, 8),
38115 => conv_std_logic_vector(131, 8),
38116 => conv_std_logic_vector(131, 8),
38117 => conv_std_logic_vector(132, 8),
38118 => conv_std_logic_vector(132, 8),
38119 => conv_std_logic_vector(133, 8),
38120 => conv_std_logic_vector(134, 8),
38121 => conv_std_logic_vector(134, 8),
38122 => conv_std_logic_vector(135, 8),
38123 => conv_std_logic_vector(135, 8),
38124 => conv_std_logic_vector(136, 8),
38125 => conv_std_logic_vector(137, 8),
38126 => conv_std_logic_vector(137, 8),
38127 => conv_std_logic_vector(138, 8),
38128 => conv_std_logic_vector(138, 8),
38129 => conv_std_logic_vector(139, 8),
38130 => conv_std_logic_vector(139, 8),
38131 => conv_std_logic_vector(140, 8),
38132 => conv_std_logic_vector(141, 8),
38133 => conv_std_logic_vector(141, 8),
38134 => conv_std_logic_vector(142, 8),
38135 => conv_std_logic_vector(142, 8),
38136 => conv_std_logic_vector(143, 8),
38137 => conv_std_logic_vector(143, 8),
38138 => conv_std_logic_vector(144, 8),
38139 => conv_std_logic_vector(145, 8),
38140 => conv_std_logic_vector(145, 8),
38141 => conv_std_logic_vector(146, 8),
38142 => conv_std_logic_vector(146, 8),
38143 => conv_std_logic_vector(147, 8),
38144 => conv_std_logic_vector(0, 8),
38145 => conv_std_logic_vector(0, 8),
38146 => conv_std_logic_vector(1, 8),
38147 => conv_std_logic_vector(1, 8),
38148 => conv_std_logic_vector(2, 8),
38149 => conv_std_logic_vector(2, 8),
38150 => conv_std_logic_vector(3, 8),
38151 => conv_std_logic_vector(4, 8),
38152 => conv_std_logic_vector(4, 8),
38153 => conv_std_logic_vector(5, 8),
38154 => conv_std_logic_vector(5, 8),
38155 => conv_std_logic_vector(6, 8),
38156 => conv_std_logic_vector(6, 8),
38157 => conv_std_logic_vector(7, 8),
38158 => conv_std_logic_vector(8, 8),
38159 => conv_std_logic_vector(8, 8),
38160 => conv_std_logic_vector(9, 8),
38161 => conv_std_logic_vector(9, 8),
38162 => conv_std_logic_vector(10, 8),
38163 => conv_std_logic_vector(11, 8),
38164 => conv_std_logic_vector(11, 8),
38165 => conv_std_logic_vector(12, 8),
38166 => conv_std_logic_vector(12, 8),
38167 => conv_std_logic_vector(13, 8),
38168 => conv_std_logic_vector(13, 8),
38169 => conv_std_logic_vector(14, 8),
38170 => conv_std_logic_vector(15, 8),
38171 => conv_std_logic_vector(15, 8),
38172 => conv_std_logic_vector(16, 8),
38173 => conv_std_logic_vector(16, 8),
38174 => conv_std_logic_vector(17, 8),
38175 => conv_std_logic_vector(18, 8),
38176 => conv_std_logic_vector(18, 8),
38177 => conv_std_logic_vector(19, 8),
38178 => conv_std_logic_vector(19, 8),
38179 => conv_std_logic_vector(20, 8),
38180 => conv_std_logic_vector(20, 8),
38181 => conv_std_logic_vector(21, 8),
38182 => conv_std_logic_vector(22, 8),
38183 => conv_std_logic_vector(22, 8),
38184 => conv_std_logic_vector(23, 8),
38185 => conv_std_logic_vector(23, 8),
38186 => conv_std_logic_vector(24, 8),
38187 => conv_std_logic_vector(25, 8),
38188 => conv_std_logic_vector(25, 8),
38189 => conv_std_logic_vector(26, 8),
38190 => conv_std_logic_vector(26, 8),
38191 => conv_std_logic_vector(27, 8),
38192 => conv_std_logic_vector(27, 8),
38193 => conv_std_logic_vector(28, 8),
38194 => conv_std_logic_vector(29, 8),
38195 => conv_std_logic_vector(29, 8),
38196 => conv_std_logic_vector(30, 8),
38197 => conv_std_logic_vector(30, 8),
38198 => conv_std_logic_vector(31, 8),
38199 => conv_std_logic_vector(32, 8),
38200 => conv_std_logic_vector(32, 8),
38201 => conv_std_logic_vector(33, 8),
38202 => conv_std_logic_vector(33, 8),
38203 => conv_std_logic_vector(34, 8),
38204 => conv_std_logic_vector(34, 8),
38205 => conv_std_logic_vector(35, 8),
38206 => conv_std_logic_vector(36, 8),
38207 => conv_std_logic_vector(36, 8),
38208 => conv_std_logic_vector(37, 8),
38209 => conv_std_logic_vector(37, 8),
38210 => conv_std_logic_vector(38, 8),
38211 => conv_std_logic_vector(38, 8),
38212 => conv_std_logic_vector(39, 8),
38213 => conv_std_logic_vector(40, 8),
38214 => conv_std_logic_vector(40, 8),
38215 => conv_std_logic_vector(41, 8),
38216 => conv_std_logic_vector(41, 8),
38217 => conv_std_logic_vector(42, 8),
38218 => conv_std_logic_vector(43, 8),
38219 => conv_std_logic_vector(43, 8),
38220 => conv_std_logic_vector(44, 8),
38221 => conv_std_logic_vector(44, 8),
38222 => conv_std_logic_vector(45, 8),
38223 => conv_std_logic_vector(45, 8),
38224 => conv_std_logic_vector(46, 8),
38225 => conv_std_logic_vector(47, 8),
38226 => conv_std_logic_vector(47, 8),
38227 => conv_std_logic_vector(48, 8),
38228 => conv_std_logic_vector(48, 8),
38229 => conv_std_logic_vector(49, 8),
38230 => conv_std_logic_vector(50, 8),
38231 => conv_std_logic_vector(50, 8),
38232 => conv_std_logic_vector(51, 8),
38233 => conv_std_logic_vector(51, 8),
38234 => conv_std_logic_vector(52, 8),
38235 => conv_std_logic_vector(52, 8),
38236 => conv_std_logic_vector(53, 8),
38237 => conv_std_logic_vector(54, 8),
38238 => conv_std_logic_vector(54, 8),
38239 => conv_std_logic_vector(55, 8),
38240 => conv_std_logic_vector(55, 8),
38241 => conv_std_logic_vector(56, 8),
38242 => conv_std_logic_vector(57, 8),
38243 => conv_std_logic_vector(57, 8),
38244 => conv_std_logic_vector(58, 8),
38245 => conv_std_logic_vector(58, 8),
38246 => conv_std_logic_vector(59, 8),
38247 => conv_std_logic_vector(59, 8),
38248 => conv_std_logic_vector(60, 8),
38249 => conv_std_logic_vector(61, 8),
38250 => conv_std_logic_vector(61, 8),
38251 => conv_std_logic_vector(62, 8),
38252 => conv_std_logic_vector(62, 8),
38253 => conv_std_logic_vector(63, 8),
38254 => conv_std_logic_vector(64, 8),
38255 => conv_std_logic_vector(64, 8),
38256 => conv_std_logic_vector(65, 8),
38257 => conv_std_logic_vector(65, 8),
38258 => conv_std_logic_vector(66, 8),
38259 => conv_std_logic_vector(66, 8),
38260 => conv_std_logic_vector(67, 8),
38261 => conv_std_logic_vector(68, 8),
38262 => conv_std_logic_vector(68, 8),
38263 => conv_std_logic_vector(69, 8),
38264 => conv_std_logic_vector(69, 8),
38265 => conv_std_logic_vector(70, 8),
38266 => conv_std_logic_vector(71, 8),
38267 => conv_std_logic_vector(71, 8),
38268 => conv_std_logic_vector(72, 8),
38269 => conv_std_logic_vector(72, 8),
38270 => conv_std_logic_vector(73, 8),
38271 => conv_std_logic_vector(73, 8),
38272 => conv_std_logic_vector(74, 8),
38273 => conv_std_logic_vector(75, 8),
38274 => conv_std_logic_vector(75, 8),
38275 => conv_std_logic_vector(76, 8),
38276 => conv_std_logic_vector(76, 8),
38277 => conv_std_logic_vector(77, 8),
38278 => conv_std_logic_vector(77, 8),
38279 => conv_std_logic_vector(78, 8),
38280 => conv_std_logic_vector(79, 8),
38281 => conv_std_logic_vector(79, 8),
38282 => conv_std_logic_vector(80, 8),
38283 => conv_std_logic_vector(80, 8),
38284 => conv_std_logic_vector(81, 8),
38285 => conv_std_logic_vector(82, 8),
38286 => conv_std_logic_vector(82, 8),
38287 => conv_std_logic_vector(83, 8),
38288 => conv_std_logic_vector(83, 8),
38289 => conv_std_logic_vector(84, 8),
38290 => conv_std_logic_vector(84, 8),
38291 => conv_std_logic_vector(85, 8),
38292 => conv_std_logic_vector(86, 8),
38293 => conv_std_logic_vector(86, 8),
38294 => conv_std_logic_vector(87, 8),
38295 => conv_std_logic_vector(87, 8),
38296 => conv_std_logic_vector(88, 8),
38297 => conv_std_logic_vector(89, 8),
38298 => conv_std_logic_vector(89, 8),
38299 => conv_std_logic_vector(90, 8),
38300 => conv_std_logic_vector(90, 8),
38301 => conv_std_logic_vector(91, 8),
38302 => conv_std_logic_vector(91, 8),
38303 => conv_std_logic_vector(92, 8),
38304 => conv_std_logic_vector(93, 8),
38305 => conv_std_logic_vector(93, 8),
38306 => conv_std_logic_vector(94, 8),
38307 => conv_std_logic_vector(94, 8),
38308 => conv_std_logic_vector(95, 8),
38309 => conv_std_logic_vector(96, 8),
38310 => conv_std_logic_vector(96, 8),
38311 => conv_std_logic_vector(97, 8),
38312 => conv_std_logic_vector(97, 8),
38313 => conv_std_logic_vector(98, 8),
38314 => conv_std_logic_vector(98, 8),
38315 => conv_std_logic_vector(99, 8),
38316 => conv_std_logic_vector(100, 8),
38317 => conv_std_logic_vector(100, 8),
38318 => conv_std_logic_vector(101, 8),
38319 => conv_std_logic_vector(101, 8),
38320 => conv_std_logic_vector(102, 8),
38321 => conv_std_logic_vector(103, 8),
38322 => conv_std_logic_vector(103, 8),
38323 => conv_std_logic_vector(104, 8),
38324 => conv_std_logic_vector(104, 8),
38325 => conv_std_logic_vector(105, 8),
38326 => conv_std_logic_vector(105, 8),
38327 => conv_std_logic_vector(106, 8),
38328 => conv_std_logic_vector(107, 8),
38329 => conv_std_logic_vector(107, 8),
38330 => conv_std_logic_vector(108, 8),
38331 => conv_std_logic_vector(108, 8),
38332 => conv_std_logic_vector(109, 8),
38333 => conv_std_logic_vector(110, 8),
38334 => conv_std_logic_vector(110, 8),
38335 => conv_std_logic_vector(111, 8),
38336 => conv_std_logic_vector(111, 8),
38337 => conv_std_logic_vector(112, 8),
38338 => conv_std_logic_vector(112, 8),
38339 => conv_std_logic_vector(113, 8),
38340 => conv_std_logic_vector(114, 8),
38341 => conv_std_logic_vector(114, 8),
38342 => conv_std_logic_vector(115, 8),
38343 => conv_std_logic_vector(115, 8),
38344 => conv_std_logic_vector(116, 8),
38345 => conv_std_logic_vector(116, 8),
38346 => conv_std_logic_vector(117, 8),
38347 => conv_std_logic_vector(118, 8),
38348 => conv_std_logic_vector(118, 8),
38349 => conv_std_logic_vector(119, 8),
38350 => conv_std_logic_vector(119, 8),
38351 => conv_std_logic_vector(120, 8),
38352 => conv_std_logic_vector(121, 8),
38353 => conv_std_logic_vector(121, 8),
38354 => conv_std_logic_vector(122, 8),
38355 => conv_std_logic_vector(122, 8),
38356 => conv_std_logic_vector(123, 8),
38357 => conv_std_logic_vector(123, 8),
38358 => conv_std_logic_vector(124, 8),
38359 => conv_std_logic_vector(125, 8),
38360 => conv_std_logic_vector(125, 8),
38361 => conv_std_logic_vector(126, 8),
38362 => conv_std_logic_vector(126, 8),
38363 => conv_std_logic_vector(127, 8),
38364 => conv_std_logic_vector(128, 8),
38365 => conv_std_logic_vector(128, 8),
38366 => conv_std_logic_vector(129, 8),
38367 => conv_std_logic_vector(129, 8),
38368 => conv_std_logic_vector(130, 8),
38369 => conv_std_logic_vector(130, 8),
38370 => conv_std_logic_vector(131, 8),
38371 => conv_std_logic_vector(132, 8),
38372 => conv_std_logic_vector(132, 8),
38373 => conv_std_logic_vector(133, 8),
38374 => conv_std_logic_vector(133, 8),
38375 => conv_std_logic_vector(134, 8),
38376 => conv_std_logic_vector(135, 8),
38377 => conv_std_logic_vector(135, 8),
38378 => conv_std_logic_vector(136, 8),
38379 => conv_std_logic_vector(136, 8),
38380 => conv_std_logic_vector(137, 8),
38381 => conv_std_logic_vector(137, 8),
38382 => conv_std_logic_vector(138, 8),
38383 => conv_std_logic_vector(139, 8),
38384 => conv_std_logic_vector(139, 8),
38385 => conv_std_logic_vector(140, 8),
38386 => conv_std_logic_vector(140, 8),
38387 => conv_std_logic_vector(141, 8),
38388 => conv_std_logic_vector(142, 8),
38389 => conv_std_logic_vector(142, 8),
38390 => conv_std_logic_vector(143, 8),
38391 => conv_std_logic_vector(143, 8),
38392 => conv_std_logic_vector(144, 8),
38393 => conv_std_logic_vector(144, 8),
38394 => conv_std_logic_vector(145, 8),
38395 => conv_std_logic_vector(146, 8),
38396 => conv_std_logic_vector(146, 8),
38397 => conv_std_logic_vector(147, 8),
38398 => conv_std_logic_vector(147, 8),
38399 => conv_std_logic_vector(148, 8),
38400 => conv_std_logic_vector(0, 8),
38401 => conv_std_logic_vector(0, 8),
38402 => conv_std_logic_vector(1, 8),
38403 => conv_std_logic_vector(1, 8),
38404 => conv_std_logic_vector(2, 8),
38405 => conv_std_logic_vector(2, 8),
38406 => conv_std_logic_vector(3, 8),
38407 => conv_std_logic_vector(4, 8),
38408 => conv_std_logic_vector(4, 8),
38409 => conv_std_logic_vector(5, 8),
38410 => conv_std_logic_vector(5, 8),
38411 => conv_std_logic_vector(6, 8),
38412 => conv_std_logic_vector(7, 8),
38413 => conv_std_logic_vector(7, 8),
38414 => conv_std_logic_vector(8, 8),
38415 => conv_std_logic_vector(8, 8),
38416 => conv_std_logic_vector(9, 8),
38417 => conv_std_logic_vector(9, 8),
38418 => conv_std_logic_vector(10, 8),
38419 => conv_std_logic_vector(11, 8),
38420 => conv_std_logic_vector(11, 8),
38421 => conv_std_logic_vector(12, 8),
38422 => conv_std_logic_vector(12, 8),
38423 => conv_std_logic_vector(13, 8),
38424 => conv_std_logic_vector(14, 8),
38425 => conv_std_logic_vector(14, 8),
38426 => conv_std_logic_vector(15, 8),
38427 => conv_std_logic_vector(15, 8),
38428 => conv_std_logic_vector(16, 8),
38429 => conv_std_logic_vector(16, 8),
38430 => conv_std_logic_vector(17, 8),
38431 => conv_std_logic_vector(18, 8),
38432 => conv_std_logic_vector(18, 8),
38433 => conv_std_logic_vector(19, 8),
38434 => conv_std_logic_vector(19, 8),
38435 => conv_std_logic_vector(20, 8),
38436 => conv_std_logic_vector(21, 8),
38437 => conv_std_logic_vector(21, 8),
38438 => conv_std_logic_vector(22, 8),
38439 => conv_std_logic_vector(22, 8),
38440 => conv_std_logic_vector(23, 8),
38441 => conv_std_logic_vector(24, 8),
38442 => conv_std_logic_vector(24, 8),
38443 => conv_std_logic_vector(25, 8),
38444 => conv_std_logic_vector(25, 8),
38445 => conv_std_logic_vector(26, 8),
38446 => conv_std_logic_vector(26, 8),
38447 => conv_std_logic_vector(27, 8),
38448 => conv_std_logic_vector(28, 8),
38449 => conv_std_logic_vector(28, 8),
38450 => conv_std_logic_vector(29, 8),
38451 => conv_std_logic_vector(29, 8),
38452 => conv_std_logic_vector(30, 8),
38453 => conv_std_logic_vector(31, 8),
38454 => conv_std_logic_vector(31, 8),
38455 => conv_std_logic_vector(32, 8),
38456 => conv_std_logic_vector(32, 8),
38457 => conv_std_logic_vector(33, 8),
38458 => conv_std_logic_vector(33, 8),
38459 => conv_std_logic_vector(34, 8),
38460 => conv_std_logic_vector(35, 8),
38461 => conv_std_logic_vector(35, 8),
38462 => conv_std_logic_vector(36, 8),
38463 => conv_std_logic_vector(36, 8),
38464 => conv_std_logic_vector(37, 8),
38465 => conv_std_logic_vector(38, 8),
38466 => conv_std_logic_vector(38, 8),
38467 => conv_std_logic_vector(39, 8),
38468 => conv_std_logic_vector(39, 8),
38469 => conv_std_logic_vector(40, 8),
38470 => conv_std_logic_vector(41, 8),
38471 => conv_std_logic_vector(41, 8),
38472 => conv_std_logic_vector(42, 8),
38473 => conv_std_logic_vector(42, 8),
38474 => conv_std_logic_vector(43, 8),
38475 => conv_std_logic_vector(43, 8),
38476 => conv_std_logic_vector(44, 8),
38477 => conv_std_logic_vector(45, 8),
38478 => conv_std_logic_vector(45, 8),
38479 => conv_std_logic_vector(46, 8),
38480 => conv_std_logic_vector(46, 8),
38481 => conv_std_logic_vector(47, 8),
38482 => conv_std_logic_vector(48, 8),
38483 => conv_std_logic_vector(48, 8),
38484 => conv_std_logic_vector(49, 8),
38485 => conv_std_logic_vector(49, 8),
38486 => conv_std_logic_vector(50, 8),
38487 => conv_std_logic_vector(50, 8),
38488 => conv_std_logic_vector(51, 8),
38489 => conv_std_logic_vector(52, 8),
38490 => conv_std_logic_vector(52, 8),
38491 => conv_std_logic_vector(53, 8),
38492 => conv_std_logic_vector(53, 8),
38493 => conv_std_logic_vector(54, 8),
38494 => conv_std_logic_vector(55, 8),
38495 => conv_std_logic_vector(55, 8),
38496 => conv_std_logic_vector(56, 8),
38497 => conv_std_logic_vector(56, 8),
38498 => conv_std_logic_vector(57, 8),
38499 => conv_std_logic_vector(58, 8),
38500 => conv_std_logic_vector(58, 8),
38501 => conv_std_logic_vector(59, 8),
38502 => conv_std_logic_vector(59, 8),
38503 => conv_std_logic_vector(60, 8),
38504 => conv_std_logic_vector(60, 8),
38505 => conv_std_logic_vector(61, 8),
38506 => conv_std_logic_vector(62, 8),
38507 => conv_std_logic_vector(62, 8),
38508 => conv_std_logic_vector(63, 8),
38509 => conv_std_logic_vector(63, 8),
38510 => conv_std_logic_vector(64, 8),
38511 => conv_std_logic_vector(65, 8),
38512 => conv_std_logic_vector(65, 8),
38513 => conv_std_logic_vector(66, 8),
38514 => conv_std_logic_vector(66, 8),
38515 => conv_std_logic_vector(67, 8),
38516 => conv_std_logic_vector(67, 8),
38517 => conv_std_logic_vector(68, 8),
38518 => conv_std_logic_vector(69, 8),
38519 => conv_std_logic_vector(69, 8),
38520 => conv_std_logic_vector(70, 8),
38521 => conv_std_logic_vector(70, 8),
38522 => conv_std_logic_vector(71, 8),
38523 => conv_std_logic_vector(72, 8),
38524 => conv_std_logic_vector(72, 8),
38525 => conv_std_logic_vector(73, 8),
38526 => conv_std_logic_vector(73, 8),
38527 => conv_std_logic_vector(74, 8),
38528 => conv_std_logic_vector(75, 8),
38529 => conv_std_logic_vector(75, 8),
38530 => conv_std_logic_vector(76, 8),
38531 => conv_std_logic_vector(76, 8),
38532 => conv_std_logic_vector(77, 8),
38533 => conv_std_logic_vector(77, 8),
38534 => conv_std_logic_vector(78, 8),
38535 => conv_std_logic_vector(79, 8),
38536 => conv_std_logic_vector(79, 8),
38537 => conv_std_logic_vector(80, 8),
38538 => conv_std_logic_vector(80, 8),
38539 => conv_std_logic_vector(81, 8),
38540 => conv_std_logic_vector(82, 8),
38541 => conv_std_logic_vector(82, 8),
38542 => conv_std_logic_vector(83, 8),
38543 => conv_std_logic_vector(83, 8),
38544 => conv_std_logic_vector(84, 8),
38545 => conv_std_logic_vector(84, 8),
38546 => conv_std_logic_vector(85, 8),
38547 => conv_std_logic_vector(86, 8),
38548 => conv_std_logic_vector(86, 8),
38549 => conv_std_logic_vector(87, 8),
38550 => conv_std_logic_vector(87, 8),
38551 => conv_std_logic_vector(88, 8),
38552 => conv_std_logic_vector(89, 8),
38553 => conv_std_logic_vector(89, 8),
38554 => conv_std_logic_vector(90, 8),
38555 => conv_std_logic_vector(90, 8),
38556 => conv_std_logic_vector(91, 8),
38557 => conv_std_logic_vector(91, 8),
38558 => conv_std_logic_vector(92, 8),
38559 => conv_std_logic_vector(93, 8),
38560 => conv_std_logic_vector(93, 8),
38561 => conv_std_logic_vector(94, 8),
38562 => conv_std_logic_vector(94, 8),
38563 => conv_std_logic_vector(95, 8),
38564 => conv_std_logic_vector(96, 8),
38565 => conv_std_logic_vector(96, 8),
38566 => conv_std_logic_vector(97, 8),
38567 => conv_std_logic_vector(97, 8),
38568 => conv_std_logic_vector(98, 8),
38569 => conv_std_logic_vector(99, 8),
38570 => conv_std_logic_vector(99, 8),
38571 => conv_std_logic_vector(100, 8),
38572 => conv_std_logic_vector(100, 8),
38573 => conv_std_logic_vector(101, 8),
38574 => conv_std_logic_vector(101, 8),
38575 => conv_std_logic_vector(102, 8),
38576 => conv_std_logic_vector(103, 8),
38577 => conv_std_logic_vector(103, 8),
38578 => conv_std_logic_vector(104, 8),
38579 => conv_std_logic_vector(104, 8),
38580 => conv_std_logic_vector(105, 8),
38581 => conv_std_logic_vector(106, 8),
38582 => conv_std_logic_vector(106, 8),
38583 => conv_std_logic_vector(107, 8),
38584 => conv_std_logic_vector(107, 8),
38585 => conv_std_logic_vector(108, 8),
38586 => conv_std_logic_vector(108, 8),
38587 => conv_std_logic_vector(109, 8),
38588 => conv_std_logic_vector(110, 8),
38589 => conv_std_logic_vector(110, 8),
38590 => conv_std_logic_vector(111, 8),
38591 => conv_std_logic_vector(111, 8),
38592 => conv_std_logic_vector(112, 8),
38593 => conv_std_logic_vector(113, 8),
38594 => conv_std_logic_vector(113, 8),
38595 => conv_std_logic_vector(114, 8),
38596 => conv_std_logic_vector(114, 8),
38597 => conv_std_logic_vector(115, 8),
38598 => conv_std_logic_vector(116, 8),
38599 => conv_std_logic_vector(116, 8),
38600 => conv_std_logic_vector(117, 8),
38601 => conv_std_logic_vector(117, 8),
38602 => conv_std_logic_vector(118, 8),
38603 => conv_std_logic_vector(118, 8),
38604 => conv_std_logic_vector(119, 8),
38605 => conv_std_logic_vector(120, 8),
38606 => conv_std_logic_vector(120, 8),
38607 => conv_std_logic_vector(121, 8),
38608 => conv_std_logic_vector(121, 8),
38609 => conv_std_logic_vector(122, 8),
38610 => conv_std_logic_vector(123, 8),
38611 => conv_std_logic_vector(123, 8),
38612 => conv_std_logic_vector(124, 8),
38613 => conv_std_logic_vector(124, 8),
38614 => conv_std_logic_vector(125, 8),
38615 => conv_std_logic_vector(125, 8),
38616 => conv_std_logic_vector(126, 8),
38617 => conv_std_logic_vector(127, 8),
38618 => conv_std_logic_vector(127, 8),
38619 => conv_std_logic_vector(128, 8),
38620 => conv_std_logic_vector(128, 8),
38621 => conv_std_logic_vector(129, 8),
38622 => conv_std_logic_vector(130, 8),
38623 => conv_std_logic_vector(130, 8),
38624 => conv_std_logic_vector(131, 8),
38625 => conv_std_logic_vector(131, 8),
38626 => conv_std_logic_vector(132, 8),
38627 => conv_std_logic_vector(133, 8),
38628 => conv_std_logic_vector(133, 8),
38629 => conv_std_logic_vector(134, 8),
38630 => conv_std_logic_vector(134, 8),
38631 => conv_std_logic_vector(135, 8),
38632 => conv_std_logic_vector(135, 8),
38633 => conv_std_logic_vector(136, 8),
38634 => conv_std_logic_vector(137, 8),
38635 => conv_std_logic_vector(137, 8),
38636 => conv_std_logic_vector(138, 8),
38637 => conv_std_logic_vector(138, 8),
38638 => conv_std_logic_vector(139, 8),
38639 => conv_std_logic_vector(140, 8),
38640 => conv_std_logic_vector(140, 8),
38641 => conv_std_logic_vector(141, 8),
38642 => conv_std_logic_vector(141, 8),
38643 => conv_std_logic_vector(142, 8),
38644 => conv_std_logic_vector(142, 8),
38645 => conv_std_logic_vector(143, 8),
38646 => conv_std_logic_vector(144, 8),
38647 => conv_std_logic_vector(144, 8),
38648 => conv_std_logic_vector(145, 8),
38649 => conv_std_logic_vector(145, 8),
38650 => conv_std_logic_vector(146, 8),
38651 => conv_std_logic_vector(147, 8),
38652 => conv_std_logic_vector(147, 8),
38653 => conv_std_logic_vector(148, 8),
38654 => conv_std_logic_vector(148, 8),
38655 => conv_std_logic_vector(149, 8),
38656 => conv_std_logic_vector(0, 8),
38657 => conv_std_logic_vector(0, 8),
38658 => conv_std_logic_vector(1, 8),
38659 => conv_std_logic_vector(1, 8),
38660 => conv_std_logic_vector(2, 8),
38661 => conv_std_logic_vector(2, 8),
38662 => conv_std_logic_vector(3, 8),
38663 => conv_std_logic_vector(4, 8),
38664 => conv_std_logic_vector(4, 8),
38665 => conv_std_logic_vector(5, 8),
38666 => conv_std_logic_vector(5, 8),
38667 => conv_std_logic_vector(6, 8),
38668 => conv_std_logic_vector(7, 8),
38669 => conv_std_logic_vector(7, 8),
38670 => conv_std_logic_vector(8, 8),
38671 => conv_std_logic_vector(8, 8),
38672 => conv_std_logic_vector(9, 8),
38673 => conv_std_logic_vector(10, 8),
38674 => conv_std_logic_vector(10, 8),
38675 => conv_std_logic_vector(11, 8),
38676 => conv_std_logic_vector(11, 8),
38677 => conv_std_logic_vector(12, 8),
38678 => conv_std_logic_vector(12, 8),
38679 => conv_std_logic_vector(13, 8),
38680 => conv_std_logic_vector(14, 8),
38681 => conv_std_logic_vector(14, 8),
38682 => conv_std_logic_vector(15, 8),
38683 => conv_std_logic_vector(15, 8),
38684 => conv_std_logic_vector(16, 8),
38685 => conv_std_logic_vector(17, 8),
38686 => conv_std_logic_vector(17, 8),
38687 => conv_std_logic_vector(18, 8),
38688 => conv_std_logic_vector(18, 8),
38689 => conv_std_logic_vector(19, 8),
38690 => conv_std_logic_vector(20, 8),
38691 => conv_std_logic_vector(20, 8),
38692 => conv_std_logic_vector(21, 8),
38693 => conv_std_logic_vector(21, 8),
38694 => conv_std_logic_vector(22, 8),
38695 => conv_std_logic_vector(23, 8),
38696 => conv_std_logic_vector(23, 8),
38697 => conv_std_logic_vector(24, 8),
38698 => conv_std_logic_vector(24, 8),
38699 => conv_std_logic_vector(25, 8),
38700 => conv_std_logic_vector(25, 8),
38701 => conv_std_logic_vector(26, 8),
38702 => conv_std_logic_vector(27, 8),
38703 => conv_std_logic_vector(27, 8),
38704 => conv_std_logic_vector(28, 8),
38705 => conv_std_logic_vector(28, 8),
38706 => conv_std_logic_vector(29, 8),
38707 => conv_std_logic_vector(30, 8),
38708 => conv_std_logic_vector(30, 8),
38709 => conv_std_logic_vector(31, 8),
38710 => conv_std_logic_vector(31, 8),
38711 => conv_std_logic_vector(32, 8),
38712 => conv_std_logic_vector(33, 8),
38713 => conv_std_logic_vector(33, 8),
38714 => conv_std_logic_vector(34, 8),
38715 => conv_std_logic_vector(34, 8),
38716 => conv_std_logic_vector(35, 8),
38717 => conv_std_logic_vector(35, 8),
38718 => conv_std_logic_vector(36, 8),
38719 => conv_std_logic_vector(37, 8),
38720 => conv_std_logic_vector(37, 8),
38721 => conv_std_logic_vector(38, 8),
38722 => conv_std_logic_vector(38, 8),
38723 => conv_std_logic_vector(39, 8),
38724 => conv_std_logic_vector(40, 8),
38725 => conv_std_logic_vector(40, 8),
38726 => conv_std_logic_vector(41, 8),
38727 => conv_std_logic_vector(41, 8),
38728 => conv_std_logic_vector(42, 8),
38729 => conv_std_logic_vector(43, 8),
38730 => conv_std_logic_vector(43, 8),
38731 => conv_std_logic_vector(44, 8),
38732 => conv_std_logic_vector(44, 8),
38733 => conv_std_logic_vector(45, 8),
38734 => conv_std_logic_vector(46, 8),
38735 => conv_std_logic_vector(46, 8),
38736 => conv_std_logic_vector(47, 8),
38737 => conv_std_logic_vector(47, 8),
38738 => conv_std_logic_vector(48, 8),
38739 => conv_std_logic_vector(48, 8),
38740 => conv_std_logic_vector(49, 8),
38741 => conv_std_logic_vector(50, 8),
38742 => conv_std_logic_vector(50, 8),
38743 => conv_std_logic_vector(51, 8),
38744 => conv_std_logic_vector(51, 8),
38745 => conv_std_logic_vector(52, 8),
38746 => conv_std_logic_vector(53, 8),
38747 => conv_std_logic_vector(53, 8),
38748 => conv_std_logic_vector(54, 8),
38749 => conv_std_logic_vector(54, 8),
38750 => conv_std_logic_vector(55, 8),
38751 => conv_std_logic_vector(56, 8),
38752 => conv_std_logic_vector(56, 8),
38753 => conv_std_logic_vector(57, 8),
38754 => conv_std_logic_vector(57, 8),
38755 => conv_std_logic_vector(58, 8),
38756 => conv_std_logic_vector(58, 8),
38757 => conv_std_logic_vector(59, 8),
38758 => conv_std_logic_vector(60, 8),
38759 => conv_std_logic_vector(60, 8),
38760 => conv_std_logic_vector(61, 8),
38761 => conv_std_logic_vector(61, 8),
38762 => conv_std_logic_vector(62, 8),
38763 => conv_std_logic_vector(63, 8),
38764 => conv_std_logic_vector(63, 8),
38765 => conv_std_logic_vector(64, 8),
38766 => conv_std_logic_vector(64, 8),
38767 => conv_std_logic_vector(65, 8),
38768 => conv_std_logic_vector(66, 8),
38769 => conv_std_logic_vector(66, 8),
38770 => conv_std_logic_vector(67, 8),
38771 => conv_std_logic_vector(67, 8),
38772 => conv_std_logic_vector(68, 8),
38773 => conv_std_logic_vector(69, 8),
38774 => conv_std_logic_vector(69, 8),
38775 => conv_std_logic_vector(70, 8),
38776 => conv_std_logic_vector(70, 8),
38777 => conv_std_logic_vector(71, 8),
38778 => conv_std_logic_vector(71, 8),
38779 => conv_std_logic_vector(72, 8),
38780 => conv_std_logic_vector(73, 8),
38781 => conv_std_logic_vector(73, 8),
38782 => conv_std_logic_vector(74, 8),
38783 => conv_std_logic_vector(74, 8),
38784 => conv_std_logic_vector(75, 8),
38785 => conv_std_logic_vector(76, 8),
38786 => conv_std_logic_vector(76, 8),
38787 => conv_std_logic_vector(77, 8),
38788 => conv_std_logic_vector(77, 8),
38789 => conv_std_logic_vector(78, 8),
38790 => conv_std_logic_vector(79, 8),
38791 => conv_std_logic_vector(79, 8),
38792 => conv_std_logic_vector(80, 8),
38793 => conv_std_logic_vector(80, 8),
38794 => conv_std_logic_vector(81, 8),
38795 => conv_std_logic_vector(81, 8),
38796 => conv_std_logic_vector(82, 8),
38797 => conv_std_logic_vector(83, 8),
38798 => conv_std_logic_vector(83, 8),
38799 => conv_std_logic_vector(84, 8),
38800 => conv_std_logic_vector(84, 8),
38801 => conv_std_logic_vector(85, 8),
38802 => conv_std_logic_vector(86, 8),
38803 => conv_std_logic_vector(86, 8),
38804 => conv_std_logic_vector(87, 8),
38805 => conv_std_logic_vector(87, 8),
38806 => conv_std_logic_vector(88, 8),
38807 => conv_std_logic_vector(89, 8),
38808 => conv_std_logic_vector(89, 8),
38809 => conv_std_logic_vector(90, 8),
38810 => conv_std_logic_vector(90, 8),
38811 => conv_std_logic_vector(91, 8),
38812 => conv_std_logic_vector(92, 8),
38813 => conv_std_logic_vector(92, 8),
38814 => conv_std_logic_vector(93, 8),
38815 => conv_std_logic_vector(93, 8),
38816 => conv_std_logic_vector(94, 8),
38817 => conv_std_logic_vector(94, 8),
38818 => conv_std_logic_vector(95, 8),
38819 => conv_std_logic_vector(96, 8),
38820 => conv_std_logic_vector(96, 8),
38821 => conv_std_logic_vector(97, 8),
38822 => conv_std_logic_vector(97, 8),
38823 => conv_std_logic_vector(98, 8),
38824 => conv_std_logic_vector(99, 8),
38825 => conv_std_logic_vector(99, 8),
38826 => conv_std_logic_vector(100, 8),
38827 => conv_std_logic_vector(100, 8),
38828 => conv_std_logic_vector(101, 8),
38829 => conv_std_logic_vector(102, 8),
38830 => conv_std_logic_vector(102, 8),
38831 => conv_std_logic_vector(103, 8),
38832 => conv_std_logic_vector(103, 8),
38833 => conv_std_logic_vector(104, 8),
38834 => conv_std_logic_vector(104, 8),
38835 => conv_std_logic_vector(105, 8),
38836 => conv_std_logic_vector(106, 8),
38837 => conv_std_logic_vector(106, 8),
38838 => conv_std_logic_vector(107, 8),
38839 => conv_std_logic_vector(107, 8),
38840 => conv_std_logic_vector(108, 8),
38841 => conv_std_logic_vector(109, 8),
38842 => conv_std_logic_vector(109, 8),
38843 => conv_std_logic_vector(110, 8),
38844 => conv_std_logic_vector(110, 8),
38845 => conv_std_logic_vector(111, 8),
38846 => conv_std_logic_vector(112, 8),
38847 => conv_std_logic_vector(112, 8),
38848 => conv_std_logic_vector(113, 8),
38849 => conv_std_logic_vector(113, 8),
38850 => conv_std_logic_vector(114, 8),
38851 => conv_std_logic_vector(115, 8),
38852 => conv_std_logic_vector(115, 8),
38853 => conv_std_logic_vector(116, 8),
38854 => conv_std_logic_vector(116, 8),
38855 => conv_std_logic_vector(117, 8),
38856 => conv_std_logic_vector(117, 8),
38857 => conv_std_logic_vector(118, 8),
38858 => conv_std_logic_vector(119, 8),
38859 => conv_std_logic_vector(119, 8),
38860 => conv_std_logic_vector(120, 8),
38861 => conv_std_logic_vector(120, 8),
38862 => conv_std_logic_vector(121, 8),
38863 => conv_std_logic_vector(122, 8),
38864 => conv_std_logic_vector(122, 8),
38865 => conv_std_logic_vector(123, 8),
38866 => conv_std_logic_vector(123, 8),
38867 => conv_std_logic_vector(124, 8),
38868 => conv_std_logic_vector(125, 8),
38869 => conv_std_logic_vector(125, 8),
38870 => conv_std_logic_vector(126, 8),
38871 => conv_std_logic_vector(126, 8),
38872 => conv_std_logic_vector(127, 8),
38873 => conv_std_logic_vector(127, 8),
38874 => conv_std_logic_vector(128, 8),
38875 => conv_std_logic_vector(129, 8),
38876 => conv_std_logic_vector(129, 8),
38877 => conv_std_logic_vector(130, 8),
38878 => conv_std_logic_vector(130, 8),
38879 => conv_std_logic_vector(131, 8),
38880 => conv_std_logic_vector(132, 8),
38881 => conv_std_logic_vector(132, 8),
38882 => conv_std_logic_vector(133, 8),
38883 => conv_std_logic_vector(133, 8),
38884 => conv_std_logic_vector(134, 8),
38885 => conv_std_logic_vector(135, 8),
38886 => conv_std_logic_vector(135, 8),
38887 => conv_std_logic_vector(136, 8),
38888 => conv_std_logic_vector(136, 8),
38889 => conv_std_logic_vector(137, 8),
38890 => conv_std_logic_vector(138, 8),
38891 => conv_std_logic_vector(138, 8),
38892 => conv_std_logic_vector(139, 8),
38893 => conv_std_logic_vector(139, 8),
38894 => conv_std_logic_vector(140, 8),
38895 => conv_std_logic_vector(140, 8),
38896 => conv_std_logic_vector(141, 8),
38897 => conv_std_logic_vector(142, 8),
38898 => conv_std_logic_vector(142, 8),
38899 => conv_std_logic_vector(143, 8),
38900 => conv_std_logic_vector(143, 8),
38901 => conv_std_logic_vector(144, 8),
38902 => conv_std_logic_vector(145, 8),
38903 => conv_std_logic_vector(145, 8),
38904 => conv_std_logic_vector(146, 8),
38905 => conv_std_logic_vector(146, 8),
38906 => conv_std_logic_vector(147, 8),
38907 => conv_std_logic_vector(148, 8),
38908 => conv_std_logic_vector(148, 8),
38909 => conv_std_logic_vector(149, 8),
38910 => conv_std_logic_vector(149, 8),
38911 => conv_std_logic_vector(150, 8),
38912 => conv_std_logic_vector(0, 8),
38913 => conv_std_logic_vector(0, 8),
38914 => conv_std_logic_vector(1, 8),
38915 => conv_std_logic_vector(1, 8),
38916 => conv_std_logic_vector(2, 8),
38917 => conv_std_logic_vector(2, 8),
38918 => conv_std_logic_vector(3, 8),
38919 => conv_std_logic_vector(4, 8),
38920 => conv_std_logic_vector(4, 8),
38921 => conv_std_logic_vector(5, 8),
38922 => conv_std_logic_vector(5, 8),
38923 => conv_std_logic_vector(6, 8),
38924 => conv_std_logic_vector(7, 8),
38925 => conv_std_logic_vector(7, 8),
38926 => conv_std_logic_vector(8, 8),
38927 => conv_std_logic_vector(8, 8),
38928 => conv_std_logic_vector(9, 8),
38929 => conv_std_logic_vector(10, 8),
38930 => conv_std_logic_vector(10, 8),
38931 => conv_std_logic_vector(11, 8),
38932 => conv_std_logic_vector(11, 8),
38933 => conv_std_logic_vector(12, 8),
38934 => conv_std_logic_vector(13, 8),
38935 => conv_std_logic_vector(13, 8),
38936 => conv_std_logic_vector(14, 8),
38937 => conv_std_logic_vector(14, 8),
38938 => conv_std_logic_vector(15, 8),
38939 => conv_std_logic_vector(16, 8),
38940 => conv_std_logic_vector(16, 8),
38941 => conv_std_logic_vector(17, 8),
38942 => conv_std_logic_vector(17, 8),
38943 => conv_std_logic_vector(18, 8),
38944 => conv_std_logic_vector(19, 8),
38945 => conv_std_logic_vector(19, 8),
38946 => conv_std_logic_vector(20, 8),
38947 => conv_std_logic_vector(20, 8),
38948 => conv_std_logic_vector(21, 8),
38949 => conv_std_logic_vector(21, 8),
38950 => conv_std_logic_vector(22, 8),
38951 => conv_std_logic_vector(23, 8),
38952 => conv_std_logic_vector(23, 8),
38953 => conv_std_logic_vector(24, 8),
38954 => conv_std_logic_vector(24, 8),
38955 => conv_std_logic_vector(25, 8),
38956 => conv_std_logic_vector(26, 8),
38957 => conv_std_logic_vector(26, 8),
38958 => conv_std_logic_vector(27, 8),
38959 => conv_std_logic_vector(27, 8),
38960 => conv_std_logic_vector(28, 8),
38961 => conv_std_logic_vector(29, 8),
38962 => conv_std_logic_vector(29, 8),
38963 => conv_std_logic_vector(30, 8),
38964 => conv_std_logic_vector(30, 8),
38965 => conv_std_logic_vector(31, 8),
38966 => conv_std_logic_vector(32, 8),
38967 => conv_std_logic_vector(32, 8),
38968 => conv_std_logic_vector(33, 8),
38969 => conv_std_logic_vector(33, 8),
38970 => conv_std_logic_vector(34, 8),
38971 => conv_std_logic_vector(35, 8),
38972 => conv_std_logic_vector(35, 8),
38973 => conv_std_logic_vector(36, 8),
38974 => conv_std_logic_vector(36, 8),
38975 => conv_std_logic_vector(37, 8),
38976 => conv_std_logic_vector(38, 8),
38977 => conv_std_logic_vector(38, 8),
38978 => conv_std_logic_vector(39, 8),
38979 => conv_std_logic_vector(39, 8),
38980 => conv_std_logic_vector(40, 8),
38981 => conv_std_logic_vector(40, 8),
38982 => conv_std_logic_vector(41, 8),
38983 => conv_std_logic_vector(42, 8),
38984 => conv_std_logic_vector(42, 8),
38985 => conv_std_logic_vector(43, 8),
38986 => conv_std_logic_vector(43, 8),
38987 => conv_std_logic_vector(44, 8),
38988 => conv_std_logic_vector(45, 8),
38989 => conv_std_logic_vector(45, 8),
38990 => conv_std_logic_vector(46, 8),
38991 => conv_std_logic_vector(46, 8),
38992 => conv_std_logic_vector(47, 8),
38993 => conv_std_logic_vector(48, 8),
38994 => conv_std_logic_vector(48, 8),
38995 => conv_std_logic_vector(49, 8),
38996 => conv_std_logic_vector(49, 8),
38997 => conv_std_logic_vector(50, 8),
38998 => conv_std_logic_vector(51, 8),
38999 => conv_std_logic_vector(51, 8),
39000 => conv_std_logic_vector(52, 8),
39001 => conv_std_logic_vector(52, 8),
39002 => conv_std_logic_vector(53, 8),
39003 => conv_std_logic_vector(54, 8),
39004 => conv_std_logic_vector(54, 8),
39005 => conv_std_logic_vector(55, 8),
39006 => conv_std_logic_vector(55, 8),
39007 => conv_std_logic_vector(56, 8),
39008 => conv_std_logic_vector(57, 8),
39009 => conv_std_logic_vector(57, 8),
39010 => conv_std_logic_vector(58, 8),
39011 => conv_std_logic_vector(58, 8),
39012 => conv_std_logic_vector(59, 8),
39013 => conv_std_logic_vector(59, 8),
39014 => conv_std_logic_vector(60, 8),
39015 => conv_std_logic_vector(61, 8),
39016 => conv_std_logic_vector(61, 8),
39017 => conv_std_logic_vector(62, 8),
39018 => conv_std_logic_vector(62, 8),
39019 => conv_std_logic_vector(63, 8),
39020 => conv_std_logic_vector(64, 8),
39021 => conv_std_logic_vector(64, 8),
39022 => conv_std_logic_vector(65, 8),
39023 => conv_std_logic_vector(65, 8),
39024 => conv_std_logic_vector(66, 8),
39025 => conv_std_logic_vector(67, 8),
39026 => conv_std_logic_vector(67, 8),
39027 => conv_std_logic_vector(68, 8),
39028 => conv_std_logic_vector(68, 8),
39029 => conv_std_logic_vector(69, 8),
39030 => conv_std_logic_vector(70, 8),
39031 => conv_std_logic_vector(70, 8),
39032 => conv_std_logic_vector(71, 8),
39033 => conv_std_logic_vector(71, 8),
39034 => conv_std_logic_vector(72, 8),
39035 => conv_std_logic_vector(73, 8),
39036 => conv_std_logic_vector(73, 8),
39037 => conv_std_logic_vector(74, 8),
39038 => conv_std_logic_vector(74, 8),
39039 => conv_std_logic_vector(75, 8),
39040 => conv_std_logic_vector(76, 8),
39041 => conv_std_logic_vector(76, 8),
39042 => conv_std_logic_vector(77, 8),
39043 => conv_std_logic_vector(77, 8),
39044 => conv_std_logic_vector(78, 8),
39045 => conv_std_logic_vector(78, 8),
39046 => conv_std_logic_vector(79, 8),
39047 => conv_std_logic_vector(80, 8),
39048 => conv_std_logic_vector(80, 8),
39049 => conv_std_logic_vector(81, 8),
39050 => conv_std_logic_vector(81, 8),
39051 => conv_std_logic_vector(82, 8),
39052 => conv_std_logic_vector(83, 8),
39053 => conv_std_logic_vector(83, 8),
39054 => conv_std_logic_vector(84, 8),
39055 => conv_std_logic_vector(84, 8),
39056 => conv_std_logic_vector(85, 8),
39057 => conv_std_logic_vector(86, 8),
39058 => conv_std_logic_vector(86, 8),
39059 => conv_std_logic_vector(87, 8),
39060 => conv_std_logic_vector(87, 8),
39061 => conv_std_logic_vector(88, 8),
39062 => conv_std_logic_vector(89, 8),
39063 => conv_std_logic_vector(89, 8),
39064 => conv_std_logic_vector(90, 8),
39065 => conv_std_logic_vector(90, 8),
39066 => conv_std_logic_vector(91, 8),
39067 => conv_std_logic_vector(92, 8),
39068 => conv_std_logic_vector(92, 8),
39069 => conv_std_logic_vector(93, 8),
39070 => conv_std_logic_vector(93, 8),
39071 => conv_std_logic_vector(94, 8),
39072 => conv_std_logic_vector(95, 8),
39073 => conv_std_logic_vector(95, 8),
39074 => conv_std_logic_vector(96, 8),
39075 => conv_std_logic_vector(96, 8),
39076 => conv_std_logic_vector(97, 8),
39077 => conv_std_logic_vector(97, 8),
39078 => conv_std_logic_vector(98, 8),
39079 => conv_std_logic_vector(99, 8),
39080 => conv_std_logic_vector(99, 8),
39081 => conv_std_logic_vector(100, 8),
39082 => conv_std_logic_vector(100, 8),
39083 => conv_std_logic_vector(101, 8),
39084 => conv_std_logic_vector(102, 8),
39085 => conv_std_logic_vector(102, 8),
39086 => conv_std_logic_vector(103, 8),
39087 => conv_std_logic_vector(103, 8),
39088 => conv_std_logic_vector(104, 8),
39089 => conv_std_logic_vector(105, 8),
39090 => conv_std_logic_vector(105, 8),
39091 => conv_std_logic_vector(106, 8),
39092 => conv_std_logic_vector(106, 8),
39093 => conv_std_logic_vector(107, 8),
39094 => conv_std_logic_vector(108, 8),
39095 => conv_std_logic_vector(108, 8),
39096 => conv_std_logic_vector(109, 8),
39097 => conv_std_logic_vector(109, 8),
39098 => conv_std_logic_vector(110, 8),
39099 => conv_std_logic_vector(111, 8),
39100 => conv_std_logic_vector(111, 8),
39101 => conv_std_logic_vector(112, 8),
39102 => conv_std_logic_vector(112, 8),
39103 => conv_std_logic_vector(113, 8),
39104 => conv_std_logic_vector(114, 8),
39105 => conv_std_logic_vector(114, 8),
39106 => conv_std_logic_vector(115, 8),
39107 => conv_std_logic_vector(115, 8),
39108 => conv_std_logic_vector(116, 8),
39109 => conv_std_logic_vector(116, 8),
39110 => conv_std_logic_vector(117, 8),
39111 => conv_std_logic_vector(118, 8),
39112 => conv_std_logic_vector(118, 8),
39113 => conv_std_logic_vector(119, 8),
39114 => conv_std_logic_vector(119, 8),
39115 => conv_std_logic_vector(120, 8),
39116 => conv_std_logic_vector(121, 8),
39117 => conv_std_logic_vector(121, 8),
39118 => conv_std_logic_vector(122, 8),
39119 => conv_std_logic_vector(122, 8),
39120 => conv_std_logic_vector(123, 8),
39121 => conv_std_logic_vector(124, 8),
39122 => conv_std_logic_vector(124, 8),
39123 => conv_std_logic_vector(125, 8),
39124 => conv_std_logic_vector(125, 8),
39125 => conv_std_logic_vector(126, 8),
39126 => conv_std_logic_vector(127, 8),
39127 => conv_std_logic_vector(127, 8),
39128 => conv_std_logic_vector(128, 8),
39129 => conv_std_logic_vector(128, 8),
39130 => conv_std_logic_vector(129, 8),
39131 => conv_std_logic_vector(130, 8),
39132 => conv_std_logic_vector(130, 8),
39133 => conv_std_logic_vector(131, 8),
39134 => conv_std_logic_vector(131, 8),
39135 => conv_std_logic_vector(132, 8),
39136 => conv_std_logic_vector(133, 8),
39137 => conv_std_logic_vector(133, 8),
39138 => conv_std_logic_vector(134, 8),
39139 => conv_std_logic_vector(134, 8),
39140 => conv_std_logic_vector(135, 8),
39141 => conv_std_logic_vector(135, 8),
39142 => conv_std_logic_vector(136, 8),
39143 => conv_std_logic_vector(137, 8),
39144 => conv_std_logic_vector(137, 8),
39145 => conv_std_logic_vector(138, 8),
39146 => conv_std_logic_vector(138, 8),
39147 => conv_std_logic_vector(139, 8),
39148 => conv_std_logic_vector(140, 8),
39149 => conv_std_logic_vector(140, 8),
39150 => conv_std_logic_vector(141, 8),
39151 => conv_std_logic_vector(141, 8),
39152 => conv_std_logic_vector(142, 8),
39153 => conv_std_logic_vector(143, 8),
39154 => conv_std_logic_vector(143, 8),
39155 => conv_std_logic_vector(144, 8),
39156 => conv_std_logic_vector(144, 8),
39157 => conv_std_logic_vector(145, 8),
39158 => conv_std_logic_vector(146, 8),
39159 => conv_std_logic_vector(146, 8),
39160 => conv_std_logic_vector(147, 8),
39161 => conv_std_logic_vector(147, 8),
39162 => conv_std_logic_vector(148, 8),
39163 => conv_std_logic_vector(149, 8),
39164 => conv_std_logic_vector(149, 8),
39165 => conv_std_logic_vector(150, 8),
39166 => conv_std_logic_vector(150, 8),
39167 => conv_std_logic_vector(151, 8),
39168 => conv_std_logic_vector(0, 8),
39169 => conv_std_logic_vector(0, 8),
39170 => conv_std_logic_vector(1, 8),
39171 => conv_std_logic_vector(1, 8),
39172 => conv_std_logic_vector(2, 8),
39173 => conv_std_logic_vector(2, 8),
39174 => conv_std_logic_vector(3, 8),
39175 => conv_std_logic_vector(4, 8),
39176 => conv_std_logic_vector(4, 8),
39177 => conv_std_logic_vector(5, 8),
39178 => conv_std_logic_vector(5, 8),
39179 => conv_std_logic_vector(6, 8),
39180 => conv_std_logic_vector(7, 8),
39181 => conv_std_logic_vector(7, 8),
39182 => conv_std_logic_vector(8, 8),
39183 => conv_std_logic_vector(8, 8),
39184 => conv_std_logic_vector(9, 8),
39185 => conv_std_logic_vector(10, 8),
39186 => conv_std_logic_vector(10, 8),
39187 => conv_std_logic_vector(11, 8),
39188 => conv_std_logic_vector(11, 8),
39189 => conv_std_logic_vector(12, 8),
39190 => conv_std_logic_vector(13, 8),
39191 => conv_std_logic_vector(13, 8),
39192 => conv_std_logic_vector(14, 8),
39193 => conv_std_logic_vector(14, 8),
39194 => conv_std_logic_vector(15, 8),
39195 => conv_std_logic_vector(16, 8),
39196 => conv_std_logic_vector(16, 8),
39197 => conv_std_logic_vector(17, 8),
39198 => conv_std_logic_vector(17, 8),
39199 => conv_std_logic_vector(18, 8),
39200 => conv_std_logic_vector(19, 8),
39201 => conv_std_logic_vector(19, 8),
39202 => conv_std_logic_vector(20, 8),
39203 => conv_std_logic_vector(20, 8),
39204 => conv_std_logic_vector(21, 8),
39205 => conv_std_logic_vector(22, 8),
39206 => conv_std_logic_vector(22, 8),
39207 => conv_std_logic_vector(23, 8),
39208 => conv_std_logic_vector(23, 8),
39209 => conv_std_logic_vector(24, 8),
39210 => conv_std_logic_vector(25, 8),
39211 => conv_std_logic_vector(25, 8),
39212 => conv_std_logic_vector(26, 8),
39213 => conv_std_logic_vector(26, 8),
39214 => conv_std_logic_vector(27, 8),
39215 => conv_std_logic_vector(28, 8),
39216 => conv_std_logic_vector(28, 8),
39217 => conv_std_logic_vector(29, 8),
39218 => conv_std_logic_vector(29, 8),
39219 => conv_std_logic_vector(30, 8),
39220 => conv_std_logic_vector(31, 8),
39221 => conv_std_logic_vector(31, 8),
39222 => conv_std_logic_vector(32, 8),
39223 => conv_std_logic_vector(32, 8),
39224 => conv_std_logic_vector(33, 8),
39225 => conv_std_logic_vector(34, 8),
39226 => conv_std_logic_vector(34, 8),
39227 => conv_std_logic_vector(35, 8),
39228 => conv_std_logic_vector(35, 8),
39229 => conv_std_logic_vector(36, 8),
39230 => conv_std_logic_vector(37, 8),
39231 => conv_std_logic_vector(37, 8),
39232 => conv_std_logic_vector(38, 8),
39233 => conv_std_logic_vector(38, 8),
39234 => conv_std_logic_vector(39, 8),
39235 => conv_std_logic_vector(40, 8),
39236 => conv_std_logic_vector(40, 8),
39237 => conv_std_logic_vector(41, 8),
39238 => conv_std_logic_vector(41, 8),
39239 => conv_std_logic_vector(42, 8),
39240 => conv_std_logic_vector(43, 8),
39241 => conv_std_logic_vector(43, 8),
39242 => conv_std_logic_vector(44, 8),
39243 => conv_std_logic_vector(44, 8),
39244 => conv_std_logic_vector(45, 8),
39245 => conv_std_logic_vector(46, 8),
39246 => conv_std_logic_vector(46, 8),
39247 => conv_std_logic_vector(47, 8),
39248 => conv_std_logic_vector(47, 8),
39249 => conv_std_logic_vector(48, 8),
39250 => conv_std_logic_vector(49, 8),
39251 => conv_std_logic_vector(49, 8),
39252 => conv_std_logic_vector(50, 8),
39253 => conv_std_logic_vector(50, 8),
39254 => conv_std_logic_vector(51, 8),
39255 => conv_std_logic_vector(51, 8),
39256 => conv_std_logic_vector(52, 8),
39257 => conv_std_logic_vector(53, 8),
39258 => conv_std_logic_vector(53, 8),
39259 => conv_std_logic_vector(54, 8),
39260 => conv_std_logic_vector(54, 8),
39261 => conv_std_logic_vector(55, 8),
39262 => conv_std_logic_vector(56, 8),
39263 => conv_std_logic_vector(56, 8),
39264 => conv_std_logic_vector(57, 8),
39265 => conv_std_logic_vector(57, 8),
39266 => conv_std_logic_vector(58, 8),
39267 => conv_std_logic_vector(59, 8),
39268 => conv_std_logic_vector(59, 8),
39269 => conv_std_logic_vector(60, 8),
39270 => conv_std_logic_vector(60, 8),
39271 => conv_std_logic_vector(61, 8),
39272 => conv_std_logic_vector(62, 8),
39273 => conv_std_logic_vector(62, 8),
39274 => conv_std_logic_vector(63, 8),
39275 => conv_std_logic_vector(63, 8),
39276 => conv_std_logic_vector(64, 8),
39277 => conv_std_logic_vector(65, 8),
39278 => conv_std_logic_vector(65, 8),
39279 => conv_std_logic_vector(66, 8),
39280 => conv_std_logic_vector(66, 8),
39281 => conv_std_logic_vector(67, 8),
39282 => conv_std_logic_vector(68, 8),
39283 => conv_std_logic_vector(68, 8),
39284 => conv_std_logic_vector(69, 8),
39285 => conv_std_logic_vector(69, 8),
39286 => conv_std_logic_vector(70, 8),
39287 => conv_std_logic_vector(71, 8),
39288 => conv_std_logic_vector(71, 8),
39289 => conv_std_logic_vector(72, 8),
39290 => conv_std_logic_vector(72, 8),
39291 => conv_std_logic_vector(73, 8),
39292 => conv_std_logic_vector(74, 8),
39293 => conv_std_logic_vector(74, 8),
39294 => conv_std_logic_vector(75, 8),
39295 => conv_std_logic_vector(75, 8),
39296 => conv_std_logic_vector(76, 8),
39297 => conv_std_logic_vector(77, 8),
39298 => conv_std_logic_vector(77, 8),
39299 => conv_std_logic_vector(78, 8),
39300 => conv_std_logic_vector(78, 8),
39301 => conv_std_logic_vector(79, 8),
39302 => conv_std_logic_vector(80, 8),
39303 => conv_std_logic_vector(80, 8),
39304 => conv_std_logic_vector(81, 8),
39305 => conv_std_logic_vector(81, 8),
39306 => conv_std_logic_vector(82, 8),
39307 => conv_std_logic_vector(83, 8),
39308 => conv_std_logic_vector(83, 8),
39309 => conv_std_logic_vector(84, 8),
39310 => conv_std_logic_vector(84, 8),
39311 => conv_std_logic_vector(85, 8),
39312 => conv_std_logic_vector(86, 8),
39313 => conv_std_logic_vector(86, 8),
39314 => conv_std_logic_vector(87, 8),
39315 => conv_std_logic_vector(87, 8),
39316 => conv_std_logic_vector(88, 8),
39317 => conv_std_logic_vector(89, 8),
39318 => conv_std_logic_vector(89, 8),
39319 => conv_std_logic_vector(90, 8),
39320 => conv_std_logic_vector(90, 8),
39321 => conv_std_logic_vector(91, 8),
39322 => conv_std_logic_vector(92, 8),
39323 => conv_std_logic_vector(92, 8),
39324 => conv_std_logic_vector(93, 8),
39325 => conv_std_logic_vector(93, 8),
39326 => conv_std_logic_vector(94, 8),
39327 => conv_std_logic_vector(95, 8),
39328 => conv_std_logic_vector(95, 8),
39329 => conv_std_logic_vector(96, 8),
39330 => conv_std_logic_vector(96, 8),
39331 => conv_std_logic_vector(97, 8),
39332 => conv_std_logic_vector(98, 8),
39333 => conv_std_logic_vector(98, 8),
39334 => conv_std_logic_vector(99, 8),
39335 => conv_std_logic_vector(99, 8),
39336 => conv_std_logic_vector(100, 8),
39337 => conv_std_logic_vector(101, 8),
39338 => conv_std_logic_vector(101, 8),
39339 => conv_std_logic_vector(102, 8),
39340 => conv_std_logic_vector(102, 8),
39341 => conv_std_logic_vector(103, 8),
39342 => conv_std_logic_vector(103, 8),
39343 => conv_std_logic_vector(104, 8),
39344 => conv_std_logic_vector(105, 8),
39345 => conv_std_logic_vector(105, 8),
39346 => conv_std_logic_vector(106, 8),
39347 => conv_std_logic_vector(106, 8),
39348 => conv_std_logic_vector(107, 8),
39349 => conv_std_logic_vector(108, 8),
39350 => conv_std_logic_vector(108, 8),
39351 => conv_std_logic_vector(109, 8),
39352 => conv_std_logic_vector(109, 8),
39353 => conv_std_logic_vector(110, 8),
39354 => conv_std_logic_vector(111, 8),
39355 => conv_std_logic_vector(111, 8),
39356 => conv_std_logic_vector(112, 8),
39357 => conv_std_logic_vector(112, 8),
39358 => conv_std_logic_vector(113, 8),
39359 => conv_std_logic_vector(114, 8),
39360 => conv_std_logic_vector(114, 8),
39361 => conv_std_logic_vector(115, 8),
39362 => conv_std_logic_vector(115, 8),
39363 => conv_std_logic_vector(116, 8),
39364 => conv_std_logic_vector(117, 8),
39365 => conv_std_logic_vector(117, 8),
39366 => conv_std_logic_vector(118, 8),
39367 => conv_std_logic_vector(118, 8),
39368 => conv_std_logic_vector(119, 8),
39369 => conv_std_logic_vector(120, 8),
39370 => conv_std_logic_vector(120, 8),
39371 => conv_std_logic_vector(121, 8),
39372 => conv_std_logic_vector(121, 8),
39373 => conv_std_logic_vector(122, 8),
39374 => conv_std_logic_vector(123, 8),
39375 => conv_std_logic_vector(123, 8),
39376 => conv_std_logic_vector(124, 8),
39377 => conv_std_logic_vector(124, 8),
39378 => conv_std_logic_vector(125, 8),
39379 => conv_std_logic_vector(126, 8),
39380 => conv_std_logic_vector(126, 8),
39381 => conv_std_logic_vector(127, 8),
39382 => conv_std_logic_vector(127, 8),
39383 => conv_std_logic_vector(128, 8),
39384 => conv_std_logic_vector(129, 8),
39385 => conv_std_logic_vector(129, 8),
39386 => conv_std_logic_vector(130, 8),
39387 => conv_std_logic_vector(130, 8),
39388 => conv_std_logic_vector(131, 8),
39389 => conv_std_logic_vector(132, 8),
39390 => conv_std_logic_vector(132, 8),
39391 => conv_std_logic_vector(133, 8),
39392 => conv_std_logic_vector(133, 8),
39393 => conv_std_logic_vector(134, 8),
39394 => conv_std_logic_vector(135, 8),
39395 => conv_std_logic_vector(135, 8),
39396 => conv_std_logic_vector(136, 8),
39397 => conv_std_logic_vector(136, 8),
39398 => conv_std_logic_vector(137, 8),
39399 => conv_std_logic_vector(138, 8),
39400 => conv_std_logic_vector(138, 8),
39401 => conv_std_logic_vector(139, 8),
39402 => conv_std_logic_vector(139, 8),
39403 => conv_std_logic_vector(140, 8),
39404 => conv_std_logic_vector(141, 8),
39405 => conv_std_logic_vector(141, 8),
39406 => conv_std_logic_vector(142, 8),
39407 => conv_std_logic_vector(142, 8),
39408 => conv_std_logic_vector(143, 8),
39409 => conv_std_logic_vector(144, 8),
39410 => conv_std_logic_vector(144, 8),
39411 => conv_std_logic_vector(145, 8),
39412 => conv_std_logic_vector(145, 8),
39413 => conv_std_logic_vector(146, 8),
39414 => conv_std_logic_vector(147, 8),
39415 => conv_std_logic_vector(147, 8),
39416 => conv_std_logic_vector(148, 8),
39417 => conv_std_logic_vector(148, 8),
39418 => conv_std_logic_vector(149, 8),
39419 => conv_std_logic_vector(150, 8),
39420 => conv_std_logic_vector(150, 8),
39421 => conv_std_logic_vector(151, 8),
39422 => conv_std_logic_vector(151, 8),
39423 => conv_std_logic_vector(152, 8),
39424 => conv_std_logic_vector(0, 8),
39425 => conv_std_logic_vector(0, 8),
39426 => conv_std_logic_vector(1, 8),
39427 => conv_std_logic_vector(1, 8),
39428 => conv_std_logic_vector(2, 8),
39429 => conv_std_logic_vector(3, 8),
39430 => conv_std_logic_vector(3, 8),
39431 => conv_std_logic_vector(4, 8),
39432 => conv_std_logic_vector(4, 8),
39433 => conv_std_logic_vector(5, 8),
39434 => conv_std_logic_vector(6, 8),
39435 => conv_std_logic_vector(6, 8),
39436 => conv_std_logic_vector(7, 8),
39437 => conv_std_logic_vector(7, 8),
39438 => conv_std_logic_vector(8, 8),
39439 => conv_std_logic_vector(9, 8),
39440 => conv_std_logic_vector(9, 8),
39441 => conv_std_logic_vector(10, 8),
39442 => conv_std_logic_vector(10, 8),
39443 => conv_std_logic_vector(11, 8),
39444 => conv_std_logic_vector(12, 8),
39445 => conv_std_logic_vector(12, 8),
39446 => conv_std_logic_vector(13, 8),
39447 => conv_std_logic_vector(13, 8),
39448 => conv_std_logic_vector(14, 8),
39449 => conv_std_logic_vector(15, 8),
39450 => conv_std_logic_vector(15, 8),
39451 => conv_std_logic_vector(16, 8),
39452 => conv_std_logic_vector(16, 8),
39453 => conv_std_logic_vector(17, 8),
39454 => conv_std_logic_vector(18, 8),
39455 => conv_std_logic_vector(18, 8),
39456 => conv_std_logic_vector(19, 8),
39457 => conv_std_logic_vector(19, 8),
39458 => conv_std_logic_vector(20, 8),
39459 => conv_std_logic_vector(21, 8),
39460 => conv_std_logic_vector(21, 8),
39461 => conv_std_logic_vector(22, 8),
39462 => conv_std_logic_vector(22, 8),
39463 => conv_std_logic_vector(23, 8),
39464 => conv_std_logic_vector(24, 8),
39465 => conv_std_logic_vector(24, 8),
39466 => conv_std_logic_vector(25, 8),
39467 => conv_std_logic_vector(25, 8),
39468 => conv_std_logic_vector(26, 8),
39469 => conv_std_logic_vector(27, 8),
39470 => conv_std_logic_vector(27, 8),
39471 => conv_std_logic_vector(28, 8),
39472 => conv_std_logic_vector(28, 8),
39473 => conv_std_logic_vector(29, 8),
39474 => conv_std_logic_vector(30, 8),
39475 => conv_std_logic_vector(30, 8),
39476 => conv_std_logic_vector(31, 8),
39477 => conv_std_logic_vector(31, 8),
39478 => conv_std_logic_vector(32, 8),
39479 => conv_std_logic_vector(33, 8),
39480 => conv_std_logic_vector(33, 8),
39481 => conv_std_logic_vector(34, 8),
39482 => conv_std_logic_vector(34, 8),
39483 => conv_std_logic_vector(35, 8),
39484 => conv_std_logic_vector(36, 8),
39485 => conv_std_logic_vector(36, 8),
39486 => conv_std_logic_vector(37, 8),
39487 => conv_std_logic_vector(37, 8),
39488 => conv_std_logic_vector(38, 8),
39489 => conv_std_logic_vector(39, 8),
39490 => conv_std_logic_vector(39, 8),
39491 => conv_std_logic_vector(40, 8),
39492 => conv_std_logic_vector(40, 8),
39493 => conv_std_logic_vector(41, 8),
39494 => conv_std_logic_vector(42, 8),
39495 => conv_std_logic_vector(42, 8),
39496 => conv_std_logic_vector(43, 8),
39497 => conv_std_logic_vector(43, 8),
39498 => conv_std_logic_vector(44, 8),
39499 => conv_std_logic_vector(45, 8),
39500 => conv_std_logic_vector(45, 8),
39501 => conv_std_logic_vector(46, 8),
39502 => conv_std_logic_vector(46, 8),
39503 => conv_std_logic_vector(47, 8),
39504 => conv_std_logic_vector(48, 8),
39505 => conv_std_logic_vector(48, 8),
39506 => conv_std_logic_vector(49, 8),
39507 => conv_std_logic_vector(49, 8),
39508 => conv_std_logic_vector(50, 8),
39509 => conv_std_logic_vector(51, 8),
39510 => conv_std_logic_vector(51, 8),
39511 => conv_std_logic_vector(52, 8),
39512 => conv_std_logic_vector(52, 8),
39513 => conv_std_logic_vector(53, 8),
39514 => conv_std_logic_vector(54, 8),
39515 => conv_std_logic_vector(54, 8),
39516 => conv_std_logic_vector(55, 8),
39517 => conv_std_logic_vector(55, 8),
39518 => conv_std_logic_vector(56, 8),
39519 => conv_std_logic_vector(57, 8),
39520 => conv_std_logic_vector(57, 8),
39521 => conv_std_logic_vector(58, 8),
39522 => conv_std_logic_vector(58, 8),
39523 => conv_std_logic_vector(59, 8),
39524 => conv_std_logic_vector(60, 8),
39525 => conv_std_logic_vector(60, 8),
39526 => conv_std_logic_vector(61, 8),
39527 => conv_std_logic_vector(61, 8),
39528 => conv_std_logic_vector(62, 8),
39529 => conv_std_logic_vector(63, 8),
39530 => conv_std_logic_vector(63, 8),
39531 => conv_std_logic_vector(64, 8),
39532 => conv_std_logic_vector(64, 8),
39533 => conv_std_logic_vector(65, 8),
39534 => conv_std_logic_vector(66, 8),
39535 => conv_std_logic_vector(66, 8),
39536 => conv_std_logic_vector(67, 8),
39537 => conv_std_logic_vector(67, 8),
39538 => conv_std_logic_vector(68, 8),
39539 => conv_std_logic_vector(69, 8),
39540 => conv_std_logic_vector(69, 8),
39541 => conv_std_logic_vector(70, 8),
39542 => conv_std_logic_vector(70, 8),
39543 => conv_std_logic_vector(71, 8),
39544 => conv_std_logic_vector(72, 8),
39545 => conv_std_logic_vector(72, 8),
39546 => conv_std_logic_vector(73, 8),
39547 => conv_std_logic_vector(73, 8),
39548 => conv_std_logic_vector(74, 8),
39549 => conv_std_logic_vector(75, 8),
39550 => conv_std_logic_vector(75, 8),
39551 => conv_std_logic_vector(76, 8),
39552 => conv_std_logic_vector(77, 8),
39553 => conv_std_logic_vector(77, 8),
39554 => conv_std_logic_vector(78, 8),
39555 => conv_std_logic_vector(78, 8),
39556 => conv_std_logic_vector(79, 8),
39557 => conv_std_logic_vector(80, 8),
39558 => conv_std_logic_vector(80, 8),
39559 => conv_std_logic_vector(81, 8),
39560 => conv_std_logic_vector(81, 8),
39561 => conv_std_logic_vector(82, 8),
39562 => conv_std_logic_vector(83, 8),
39563 => conv_std_logic_vector(83, 8),
39564 => conv_std_logic_vector(84, 8),
39565 => conv_std_logic_vector(84, 8),
39566 => conv_std_logic_vector(85, 8),
39567 => conv_std_logic_vector(86, 8),
39568 => conv_std_logic_vector(86, 8),
39569 => conv_std_logic_vector(87, 8),
39570 => conv_std_logic_vector(87, 8),
39571 => conv_std_logic_vector(88, 8),
39572 => conv_std_logic_vector(89, 8),
39573 => conv_std_logic_vector(89, 8),
39574 => conv_std_logic_vector(90, 8),
39575 => conv_std_logic_vector(90, 8),
39576 => conv_std_logic_vector(91, 8),
39577 => conv_std_logic_vector(92, 8),
39578 => conv_std_logic_vector(92, 8),
39579 => conv_std_logic_vector(93, 8),
39580 => conv_std_logic_vector(93, 8),
39581 => conv_std_logic_vector(94, 8),
39582 => conv_std_logic_vector(95, 8),
39583 => conv_std_logic_vector(95, 8),
39584 => conv_std_logic_vector(96, 8),
39585 => conv_std_logic_vector(96, 8),
39586 => conv_std_logic_vector(97, 8),
39587 => conv_std_logic_vector(98, 8),
39588 => conv_std_logic_vector(98, 8),
39589 => conv_std_logic_vector(99, 8),
39590 => conv_std_logic_vector(99, 8),
39591 => conv_std_logic_vector(100, 8),
39592 => conv_std_logic_vector(101, 8),
39593 => conv_std_logic_vector(101, 8),
39594 => conv_std_logic_vector(102, 8),
39595 => conv_std_logic_vector(102, 8),
39596 => conv_std_logic_vector(103, 8),
39597 => conv_std_logic_vector(104, 8),
39598 => conv_std_logic_vector(104, 8),
39599 => conv_std_logic_vector(105, 8),
39600 => conv_std_logic_vector(105, 8),
39601 => conv_std_logic_vector(106, 8),
39602 => conv_std_logic_vector(107, 8),
39603 => conv_std_logic_vector(107, 8),
39604 => conv_std_logic_vector(108, 8),
39605 => conv_std_logic_vector(108, 8),
39606 => conv_std_logic_vector(109, 8),
39607 => conv_std_logic_vector(110, 8),
39608 => conv_std_logic_vector(110, 8),
39609 => conv_std_logic_vector(111, 8),
39610 => conv_std_logic_vector(111, 8),
39611 => conv_std_logic_vector(112, 8),
39612 => conv_std_logic_vector(113, 8),
39613 => conv_std_logic_vector(113, 8),
39614 => conv_std_logic_vector(114, 8),
39615 => conv_std_logic_vector(114, 8),
39616 => conv_std_logic_vector(115, 8),
39617 => conv_std_logic_vector(116, 8),
39618 => conv_std_logic_vector(116, 8),
39619 => conv_std_logic_vector(117, 8),
39620 => conv_std_logic_vector(117, 8),
39621 => conv_std_logic_vector(118, 8),
39622 => conv_std_logic_vector(119, 8),
39623 => conv_std_logic_vector(119, 8),
39624 => conv_std_logic_vector(120, 8),
39625 => conv_std_logic_vector(120, 8),
39626 => conv_std_logic_vector(121, 8),
39627 => conv_std_logic_vector(122, 8),
39628 => conv_std_logic_vector(122, 8),
39629 => conv_std_logic_vector(123, 8),
39630 => conv_std_logic_vector(123, 8),
39631 => conv_std_logic_vector(124, 8),
39632 => conv_std_logic_vector(125, 8),
39633 => conv_std_logic_vector(125, 8),
39634 => conv_std_logic_vector(126, 8),
39635 => conv_std_logic_vector(126, 8),
39636 => conv_std_logic_vector(127, 8),
39637 => conv_std_logic_vector(128, 8),
39638 => conv_std_logic_vector(128, 8),
39639 => conv_std_logic_vector(129, 8),
39640 => conv_std_logic_vector(129, 8),
39641 => conv_std_logic_vector(130, 8),
39642 => conv_std_logic_vector(131, 8),
39643 => conv_std_logic_vector(131, 8),
39644 => conv_std_logic_vector(132, 8),
39645 => conv_std_logic_vector(132, 8),
39646 => conv_std_logic_vector(133, 8),
39647 => conv_std_logic_vector(134, 8),
39648 => conv_std_logic_vector(134, 8),
39649 => conv_std_logic_vector(135, 8),
39650 => conv_std_logic_vector(135, 8),
39651 => conv_std_logic_vector(136, 8),
39652 => conv_std_logic_vector(137, 8),
39653 => conv_std_logic_vector(137, 8),
39654 => conv_std_logic_vector(138, 8),
39655 => conv_std_logic_vector(138, 8),
39656 => conv_std_logic_vector(139, 8),
39657 => conv_std_logic_vector(140, 8),
39658 => conv_std_logic_vector(140, 8),
39659 => conv_std_logic_vector(141, 8),
39660 => conv_std_logic_vector(141, 8),
39661 => conv_std_logic_vector(142, 8),
39662 => conv_std_logic_vector(143, 8),
39663 => conv_std_logic_vector(143, 8),
39664 => conv_std_logic_vector(144, 8),
39665 => conv_std_logic_vector(144, 8),
39666 => conv_std_logic_vector(145, 8),
39667 => conv_std_logic_vector(146, 8),
39668 => conv_std_logic_vector(146, 8),
39669 => conv_std_logic_vector(147, 8),
39670 => conv_std_logic_vector(147, 8),
39671 => conv_std_logic_vector(148, 8),
39672 => conv_std_logic_vector(149, 8),
39673 => conv_std_logic_vector(149, 8),
39674 => conv_std_logic_vector(150, 8),
39675 => conv_std_logic_vector(150, 8),
39676 => conv_std_logic_vector(151, 8),
39677 => conv_std_logic_vector(152, 8),
39678 => conv_std_logic_vector(152, 8),
39679 => conv_std_logic_vector(153, 8),
39680 => conv_std_logic_vector(0, 8),
39681 => conv_std_logic_vector(0, 8),
39682 => conv_std_logic_vector(1, 8),
39683 => conv_std_logic_vector(1, 8),
39684 => conv_std_logic_vector(2, 8),
39685 => conv_std_logic_vector(3, 8),
39686 => conv_std_logic_vector(3, 8),
39687 => conv_std_logic_vector(4, 8),
39688 => conv_std_logic_vector(4, 8),
39689 => conv_std_logic_vector(5, 8),
39690 => conv_std_logic_vector(6, 8),
39691 => conv_std_logic_vector(6, 8),
39692 => conv_std_logic_vector(7, 8),
39693 => conv_std_logic_vector(7, 8),
39694 => conv_std_logic_vector(8, 8),
39695 => conv_std_logic_vector(9, 8),
39696 => conv_std_logic_vector(9, 8),
39697 => conv_std_logic_vector(10, 8),
39698 => conv_std_logic_vector(10, 8),
39699 => conv_std_logic_vector(11, 8),
39700 => conv_std_logic_vector(12, 8),
39701 => conv_std_logic_vector(12, 8),
39702 => conv_std_logic_vector(13, 8),
39703 => conv_std_logic_vector(13, 8),
39704 => conv_std_logic_vector(14, 8),
39705 => conv_std_logic_vector(15, 8),
39706 => conv_std_logic_vector(15, 8),
39707 => conv_std_logic_vector(16, 8),
39708 => conv_std_logic_vector(16, 8),
39709 => conv_std_logic_vector(17, 8),
39710 => conv_std_logic_vector(18, 8),
39711 => conv_std_logic_vector(18, 8),
39712 => conv_std_logic_vector(19, 8),
39713 => conv_std_logic_vector(19, 8),
39714 => conv_std_logic_vector(20, 8),
39715 => conv_std_logic_vector(21, 8),
39716 => conv_std_logic_vector(21, 8),
39717 => conv_std_logic_vector(22, 8),
39718 => conv_std_logic_vector(23, 8),
39719 => conv_std_logic_vector(23, 8),
39720 => conv_std_logic_vector(24, 8),
39721 => conv_std_logic_vector(24, 8),
39722 => conv_std_logic_vector(25, 8),
39723 => conv_std_logic_vector(26, 8),
39724 => conv_std_logic_vector(26, 8),
39725 => conv_std_logic_vector(27, 8),
39726 => conv_std_logic_vector(27, 8),
39727 => conv_std_logic_vector(28, 8),
39728 => conv_std_logic_vector(29, 8),
39729 => conv_std_logic_vector(29, 8),
39730 => conv_std_logic_vector(30, 8),
39731 => conv_std_logic_vector(30, 8),
39732 => conv_std_logic_vector(31, 8),
39733 => conv_std_logic_vector(32, 8),
39734 => conv_std_logic_vector(32, 8),
39735 => conv_std_logic_vector(33, 8),
39736 => conv_std_logic_vector(33, 8),
39737 => conv_std_logic_vector(34, 8),
39738 => conv_std_logic_vector(35, 8),
39739 => conv_std_logic_vector(35, 8),
39740 => conv_std_logic_vector(36, 8),
39741 => conv_std_logic_vector(36, 8),
39742 => conv_std_logic_vector(37, 8),
39743 => conv_std_logic_vector(38, 8),
39744 => conv_std_logic_vector(38, 8),
39745 => conv_std_logic_vector(39, 8),
39746 => conv_std_logic_vector(39, 8),
39747 => conv_std_logic_vector(40, 8),
39748 => conv_std_logic_vector(41, 8),
39749 => conv_std_logic_vector(41, 8),
39750 => conv_std_logic_vector(42, 8),
39751 => conv_std_logic_vector(42, 8),
39752 => conv_std_logic_vector(43, 8),
39753 => conv_std_logic_vector(44, 8),
39754 => conv_std_logic_vector(44, 8),
39755 => conv_std_logic_vector(45, 8),
39756 => conv_std_logic_vector(46, 8),
39757 => conv_std_logic_vector(46, 8),
39758 => conv_std_logic_vector(47, 8),
39759 => conv_std_logic_vector(47, 8),
39760 => conv_std_logic_vector(48, 8),
39761 => conv_std_logic_vector(49, 8),
39762 => conv_std_logic_vector(49, 8),
39763 => conv_std_logic_vector(50, 8),
39764 => conv_std_logic_vector(50, 8),
39765 => conv_std_logic_vector(51, 8),
39766 => conv_std_logic_vector(52, 8),
39767 => conv_std_logic_vector(52, 8),
39768 => conv_std_logic_vector(53, 8),
39769 => conv_std_logic_vector(53, 8),
39770 => conv_std_logic_vector(54, 8),
39771 => conv_std_logic_vector(55, 8),
39772 => conv_std_logic_vector(55, 8),
39773 => conv_std_logic_vector(56, 8),
39774 => conv_std_logic_vector(56, 8),
39775 => conv_std_logic_vector(57, 8),
39776 => conv_std_logic_vector(58, 8),
39777 => conv_std_logic_vector(58, 8),
39778 => conv_std_logic_vector(59, 8),
39779 => conv_std_logic_vector(59, 8),
39780 => conv_std_logic_vector(60, 8),
39781 => conv_std_logic_vector(61, 8),
39782 => conv_std_logic_vector(61, 8),
39783 => conv_std_logic_vector(62, 8),
39784 => conv_std_logic_vector(62, 8),
39785 => conv_std_logic_vector(63, 8),
39786 => conv_std_logic_vector(64, 8),
39787 => conv_std_logic_vector(64, 8),
39788 => conv_std_logic_vector(65, 8),
39789 => conv_std_logic_vector(65, 8),
39790 => conv_std_logic_vector(66, 8),
39791 => conv_std_logic_vector(67, 8),
39792 => conv_std_logic_vector(67, 8),
39793 => conv_std_logic_vector(68, 8),
39794 => conv_std_logic_vector(69, 8),
39795 => conv_std_logic_vector(69, 8),
39796 => conv_std_logic_vector(70, 8),
39797 => conv_std_logic_vector(70, 8),
39798 => conv_std_logic_vector(71, 8),
39799 => conv_std_logic_vector(72, 8),
39800 => conv_std_logic_vector(72, 8),
39801 => conv_std_logic_vector(73, 8),
39802 => conv_std_logic_vector(73, 8),
39803 => conv_std_logic_vector(74, 8),
39804 => conv_std_logic_vector(75, 8),
39805 => conv_std_logic_vector(75, 8),
39806 => conv_std_logic_vector(76, 8),
39807 => conv_std_logic_vector(76, 8),
39808 => conv_std_logic_vector(77, 8),
39809 => conv_std_logic_vector(78, 8),
39810 => conv_std_logic_vector(78, 8),
39811 => conv_std_logic_vector(79, 8),
39812 => conv_std_logic_vector(79, 8),
39813 => conv_std_logic_vector(80, 8),
39814 => conv_std_logic_vector(81, 8),
39815 => conv_std_logic_vector(81, 8),
39816 => conv_std_logic_vector(82, 8),
39817 => conv_std_logic_vector(82, 8),
39818 => conv_std_logic_vector(83, 8),
39819 => conv_std_logic_vector(84, 8),
39820 => conv_std_logic_vector(84, 8),
39821 => conv_std_logic_vector(85, 8),
39822 => conv_std_logic_vector(85, 8),
39823 => conv_std_logic_vector(86, 8),
39824 => conv_std_logic_vector(87, 8),
39825 => conv_std_logic_vector(87, 8),
39826 => conv_std_logic_vector(88, 8),
39827 => conv_std_logic_vector(89, 8),
39828 => conv_std_logic_vector(89, 8),
39829 => conv_std_logic_vector(90, 8),
39830 => conv_std_logic_vector(90, 8),
39831 => conv_std_logic_vector(91, 8),
39832 => conv_std_logic_vector(92, 8),
39833 => conv_std_logic_vector(92, 8),
39834 => conv_std_logic_vector(93, 8),
39835 => conv_std_logic_vector(93, 8),
39836 => conv_std_logic_vector(94, 8),
39837 => conv_std_logic_vector(95, 8),
39838 => conv_std_logic_vector(95, 8),
39839 => conv_std_logic_vector(96, 8),
39840 => conv_std_logic_vector(96, 8),
39841 => conv_std_logic_vector(97, 8),
39842 => conv_std_logic_vector(98, 8),
39843 => conv_std_logic_vector(98, 8),
39844 => conv_std_logic_vector(99, 8),
39845 => conv_std_logic_vector(99, 8),
39846 => conv_std_logic_vector(100, 8),
39847 => conv_std_logic_vector(101, 8),
39848 => conv_std_logic_vector(101, 8),
39849 => conv_std_logic_vector(102, 8),
39850 => conv_std_logic_vector(102, 8),
39851 => conv_std_logic_vector(103, 8),
39852 => conv_std_logic_vector(104, 8),
39853 => conv_std_logic_vector(104, 8),
39854 => conv_std_logic_vector(105, 8),
39855 => conv_std_logic_vector(105, 8),
39856 => conv_std_logic_vector(106, 8),
39857 => conv_std_logic_vector(107, 8),
39858 => conv_std_logic_vector(107, 8),
39859 => conv_std_logic_vector(108, 8),
39860 => conv_std_logic_vector(108, 8),
39861 => conv_std_logic_vector(109, 8),
39862 => conv_std_logic_vector(110, 8),
39863 => conv_std_logic_vector(110, 8),
39864 => conv_std_logic_vector(111, 8),
39865 => conv_std_logic_vector(112, 8),
39866 => conv_std_logic_vector(112, 8),
39867 => conv_std_logic_vector(113, 8),
39868 => conv_std_logic_vector(113, 8),
39869 => conv_std_logic_vector(114, 8),
39870 => conv_std_logic_vector(115, 8),
39871 => conv_std_logic_vector(115, 8),
39872 => conv_std_logic_vector(116, 8),
39873 => conv_std_logic_vector(116, 8),
39874 => conv_std_logic_vector(117, 8),
39875 => conv_std_logic_vector(118, 8),
39876 => conv_std_logic_vector(118, 8),
39877 => conv_std_logic_vector(119, 8),
39878 => conv_std_logic_vector(119, 8),
39879 => conv_std_logic_vector(120, 8),
39880 => conv_std_logic_vector(121, 8),
39881 => conv_std_logic_vector(121, 8),
39882 => conv_std_logic_vector(122, 8),
39883 => conv_std_logic_vector(122, 8),
39884 => conv_std_logic_vector(123, 8),
39885 => conv_std_logic_vector(124, 8),
39886 => conv_std_logic_vector(124, 8),
39887 => conv_std_logic_vector(125, 8),
39888 => conv_std_logic_vector(125, 8),
39889 => conv_std_logic_vector(126, 8),
39890 => conv_std_logic_vector(127, 8),
39891 => conv_std_logic_vector(127, 8),
39892 => conv_std_logic_vector(128, 8),
39893 => conv_std_logic_vector(128, 8),
39894 => conv_std_logic_vector(129, 8),
39895 => conv_std_logic_vector(130, 8),
39896 => conv_std_logic_vector(130, 8),
39897 => conv_std_logic_vector(131, 8),
39898 => conv_std_logic_vector(131, 8),
39899 => conv_std_logic_vector(132, 8),
39900 => conv_std_logic_vector(133, 8),
39901 => conv_std_logic_vector(133, 8),
39902 => conv_std_logic_vector(134, 8),
39903 => conv_std_logic_vector(135, 8),
39904 => conv_std_logic_vector(135, 8),
39905 => conv_std_logic_vector(136, 8),
39906 => conv_std_logic_vector(136, 8),
39907 => conv_std_logic_vector(137, 8),
39908 => conv_std_logic_vector(138, 8),
39909 => conv_std_logic_vector(138, 8),
39910 => conv_std_logic_vector(139, 8),
39911 => conv_std_logic_vector(139, 8),
39912 => conv_std_logic_vector(140, 8),
39913 => conv_std_logic_vector(141, 8),
39914 => conv_std_logic_vector(141, 8),
39915 => conv_std_logic_vector(142, 8),
39916 => conv_std_logic_vector(142, 8),
39917 => conv_std_logic_vector(143, 8),
39918 => conv_std_logic_vector(144, 8),
39919 => conv_std_logic_vector(144, 8),
39920 => conv_std_logic_vector(145, 8),
39921 => conv_std_logic_vector(145, 8),
39922 => conv_std_logic_vector(146, 8),
39923 => conv_std_logic_vector(147, 8),
39924 => conv_std_logic_vector(147, 8),
39925 => conv_std_logic_vector(148, 8),
39926 => conv_std_logic_vector(148, 8),
39927 => conv_std_logic_vector(149, 8),
39928 => conv_std_logic_vector(150, 8),
39929 => conv_std_logic_vector(150, 8),
39930 => conv_std_logic_vector(151, 8),
39931 => conv_std_logic_vector(151, 8),
39932 => conv_std_logic_vector(152, 8),
39933 => conv_std_logic_vector(153, 8),
39934 => conv_std_logic_vector(153, 8),
39935 => conv_std_logic_vector(154, 8),
39936 => conv_std_logic_vector(0, 8),
39937 => conv_std_logic_vector(0, 8),
39938 => conv_std_logic_vector(1, 8),
39939 => conv_std_logic_vector(1, 8),
39940 => conv_std_logic_vector(2, 8),
39941 => conv_std_logic_vector(3, 8),
39942 => conv_std_logic_vector(3, 8),
39943 => conv_std_logic_vector(4, 8),
39944 => conv_std_logic_vector(4, 8),
39945 => conv_std_logic_vector(5, 8),
39946 => conv_std_logic_vector(6, 8),
39947 => conv_std_logic_vector(6, 8),
39948 => conv_std_logic_vector(7, 8),
39949 => conv_std_logic_vector(7, 8),
39950 => conv_std_logic_vector(8, 8),
39951 => conv_std_logic_vector(9, 8),
39952 => conv_std_logic_vector(9, 8),
39953 => conv_std_logic_vector(10, 8),
39954 => conv_std_logic_vector(10, 8),
39955 => conv_std_logic_vector(11, 8),
39956 => conv_std_logic_vector(12, 8),
39957 => conv_std_logic_vector(12, 8),
39958 => conv_std_logic_vector(13, 8),
39959 => conv_std_logic_vector(14, 8),
39960 => conv_std_logic_vector(14, 8),
39961 => conv_std_logic_vector(15, 8),
39962 => conv_std_logic_vector(15, 8),
39963 => conv_std_logic_vector(16, 8),
39964 => conv_std_logic_vector(17, 8),
39965 => conv_std_logic_vector(17, 8),
39966 => conv_std_logic_vector(18, 8),
39967 => conv_std_logic_vector(18, 8),
39968 => conv_std_logic_vector(19, 8),
39969 => conv_std_logic_vector(20, 8),
39970 => conv_std_logic_vector(20, 8),
39971 => conv_std_logic_vector(21, 8),
39972 => conv_std_logic_vector(21, 8),
39973 => conv_std_logic_vector(22, 8),
39974 => conv_std_logic_vector(23, 8),
39975 => conv_std_logic_vector(23, 8),
39976 => conv_std_logic_vector(24, 8),
39977 => conv_std_logic_vector(24, 8),
39978 => conv_std_logic_vector(25, 8),
39979 => conv_std_logic_vector(26, 8),
39980 => conv_std_logic_vector(26, 8),
39981 => conv_std_logic_vector(27, 8),
39982 => conv_std_logic_vector(28, 8),
39983 => conv_std_logic_vector(28, 8),
39984 => conv_std_logic_vector(29, 8),
39985 => conv_std_logic_vector(29, 8),
39986 => conv_std_logic_vector(30, 8),
39987 => conv_std_logic_vector(31, 8),
39988 => conv_std_logic_vector(31, 8),
39989 => conv_std_logic_vector(32, 8),
39990 => conv_std_logic_vector(32, 8),
39991 => conv_std_logic_vector(33, 8),
39992 => conv_std_logic_vector(34, 8),
39993 => conv_std_logic_vector(34, 8),
39994 => conv_std_logic_vector(35, 8),
39995 => conv_std_logic_vector(35, 8),
39996 => conv_std_logic_vector(36, 8),
39997 => conv_std_logic_vector(37, 8),
39998 => conv_std_logic_vector(37, 8),
39999 => conv_std_logic_vector(38, 8),
40000 => conv_std_logic_vector(39, 8),
40001 => conv_std_logic_vector(39, 8),
40002 => conv_std_logic_vector(40, 8),
40003 => conv_std_logic_vector(40, 8),
40004 => conv_std_logic_vector(41, 8),
40005 => conv_std_logic_vector(42, 8),
40006 => conv_std_logic_vector(42, 8),
40007 => conv_std_logic_vector(43, 8),
40008 => conv_std_logic_vector(43, 8),
40009 => conv_std_logic_vector(44, 8),
40010 => conv_std_logic_vector(45, 8),
40011 => conv_std_logic_vector(45, 8),
40012 => conv_std_logic_vector(46, 8),
40013 => conv_std_logic_vector(46, 8),
40014 => conv_std_logic_vector(47, 8),
40015 => conv_std_logic_vector(48, 8),
40016 => conv_std_logic_vector(48, 8),
40017 => conv_std_logic_vector(49, 8),
40018 => conv_std_logic_vector(49, 8),
40019 => conv_std_logic_vector(50, 8),
40020 => conv_std_logic_vector(51, 8),
40021 => conv_std_logic_vector(51, 8),
40022 => conv_std_logic_vector(52, 8),
40023 => conv_std_logic_vector(53, 8),
40024 => conv_std_logic_vector(53, 8),
40025 => conv_std_logic_vector(54, 8),
40026 => conv_std_logic_vector(54, 8),
40027 => conv_std_logic_vector(55, 8),
40028 => conv_std_logic_vector(56, 8),
40029 => conv_std_logic_vector(56, 8),
40030 => conv_std_logic_vector(57, 8),
40031 => conv_std_logic_vector(57, 8),
40032 => conv_std_logic_vector(58, 8),
40033 => conv_std_logic_vector(59, 8),
40034 => conv_std_logic_vector(59, 8),
40035 => conv_std_logic_vector(60, 8),
40036 => conv_std_logic_vector(60, 8),
40037 => conv_std_logic_vector(61, 8),
40038 => conv_std_logic_vector(62, 8),
40039 => conv_std_logic_vector(62, 8),
40040 => conv_std_logic_vector(63, 8),
40041 => conv_std_logic_vector(63, 8),
40042 => conv_std_logic_vector(64, 8),
40043 => conv_std_logic_vector(65, 8),
40044 => conv_std_logic_vector(65, 8),
40045 => conv_std_logic_vector(66, 8),
40046 => conv_std_logic_vector(67, 8),
40047 => conv_std_logic_vector(67, 8),
40048 => conv_std_logic_vector(68, 8),
40049 => conv_std_logic_vector(68, 8),
40050 => conv_std_logic_vector(69, 8),
40051 => conv_std_logic_vector(70, 8),
40052 => conv_std_logic_vector(70, 8),
40053 => conv_std_logic_vector(71, 8),
40054 => conv_std_logic_vector(71, 8),
40055 => conv_std_logic_vector(72, 8),
40056 => conv_std_logic_vector(73, 8),
40057 => conv_std_logic_vector(73, 8),
40058 => conv_std_logic_vector(74, 8),
40059 => conv_std_logic_vector(74, 8),
40060 => conv_std_logic_vector(75, 8),
40061 => conv_std_logic_vector(76, 8),
40062 => conv_std_logic_vector(76, 8),
40063 => conv_std_logic_vector(77, 8),
40064 => conv_std_logic_vector(78, 8),
40065 => conv_std_logic_vector(78, 8),
40066 => conv_std_logic_vector(79, 8),
40067 => conv_std_logic_vector(79, 8),
40068 => conv_std_logic_vector(80, 8),
40069 => conv_std_logic_vector(81, 8),
40070 => conv_std_logic_vector(81, 8),
40071 => conv_std_logic_vector(82, 8),
40072 => conv_std_logic_vector(82, 8),
40073 => conv_std_logic_vector(83, 8),
40074 => conv_std_logic_vector(84, 8),
40075 => conv_std_logic_vector(84, 8),
40076 => conv_std_logic_vector(85, 8),
40077 => conv_std_logic_vector(85, 8),
40078 => conv_std_logic_vector(86, 8),
40079 => conv_std_logic_vector(87, 8),
40080 => conv_std_logic_vector(87, 8),
40081 => conv_std_logic_vector(88, 8),
40082 => conv_std_logic_vector(88, 8),
40083 => conv_std_logic_vector(89, 8),
40084 => conv_std_logic_vector(90, 8),
40085 => conv_std_logic_vector(90, 8),
40086 => conv_std_logic_vector(91, 8),
40087 => conv_std_logic_vector(92, 8),
40088 => conv_std_logic_vector(92, 8),
40089 => conv_std_logic_vector(93, 8),
40090 => conv_std_logic_vector(93, 8),
40091 => conv_std_logic_vector(94, 8),
40092 => conv_std_logic_vector(95, 8),
40093 => conv_std_logic_vector(95, 8),
40094 => conv_std_logic_vector(96, 8),
40095 => conv_std_logic_vector(96, 8),
40096 => conv_std_logic_vector(97, 8),
40097 => conv_std_logic_vector(98, 8),
40098 => conv_std_logic_vector(98, 8),
40099 => conv_std_logic_vector(99, 8),
40100 => conv_std_logic_vector(99, 8),
40101 => conv_std_logic_vector(100, 8),
40102 => conv_std_logic_vector(101, 8),
40103 => conv_std_logic_vector(101, 8),
40104 => conv_std_logic_vector(102, 8),
40105 => conv_std_logic_vector(102, 8),
40106 => conv_std_logic_vector(103, 8),
40107 => conv_std_logic_vector(104, 8),
40108 => conv_std_logic_vector(104, 8),
40109 => conv_std_logic_vector(105, 8),
40110 => conv_std_logic_vector(106, 8),
40111 => conv_std_logic_vector(106, 8),
40112 => conv_std_logic_vector(107, 8),
40113 => conv_std_logic_vector(107, 8),
40114 => conv_std_logic_vector(108, 8),
40115 => conv_std_logic_vector(109, 8),
40116 => conv_std_logic_vector(109, 8),
40117 => conv_std_logic_vector(110, 8),
40118 => conv_std_logic_vector(110, 8),
40119 => conv_std_logic_vector(111, 8),
40120 => conv_std_logic_vector(112, 8),
40121 => conv_std_logic_vector(112, 8),
40122 => conv_std_logic_vector(113, 8),
40123 => conv_std_logic_vector(113, 8),
40124 => conv_std_logic_vector(114, 8),
40125 => conv_std_logic_vector(115, 8),
40126 => conv_std_logic_vector(115, 8),
40127 => conv_std_logic_vector(116, 8),
40128 => conv_std_logic_vector(117, 8),
40129 => conv_std_logic_vector(117, 8),
40130 => conv_std_logic_vector(118, 8),
40131 => conv_std_logic_vector(118, 8),
40132 => conv_std_logic_vector(119, 8),
40133 => conv_std_logic_vector(120, 8),
40134 => conv_std_logic_vector(120, 8),
40135 => conv_std_logic_vector(121, 8),
40136 => conv_std_logic_vector(121, 8),
40137 => conv_std_logic_vector(122, 8),
40138 => conv_std_logic_vector(123, 8),
40139 => conv_std_logic_vector(123, 8),
40140 => conv_std_logic_vector(124, 8),
40141 => conv_std_logic_vector(124, 8),
40142 => conv_std_logic_vector(125, 8),
40143 => conv_std_logic_vector(126, 8),
40144 => conv_std_logic_vector(126, 8),
40145 => conv_std_logic_vector(127, 8),
40146 => conv_std_logic_vector(127, 8),
40147 => conv_std_logic_vector(128, 8),
40148 => conv_std_logic_vector(129, 8),
40149 => conv_std_logic_vector(129, 8),
40150 => conv_std_logic_vector(130, 8),
40151 => conv_std_logic_vector(131, 8),
40152 => conv_std_logic_vector(131, 8),
40153 => conv_std_logic_vector(132, 8),
40154 => conv_std_logic_vector(132, 8),
40155 => conv_std_logic_vector(133, 8),
40156 => conv_std_logic_vector(134, 8),
40157 => conv_std_logic_vector(134, 8),
40158 => conv_std_logic_vector(135, 8),
40159 => conv_std_logic_vector(135, 8),
40160 => conv_std_logic_vector(136, 8),
40161 => conv_std_logic_vector(137, 8),
40162 => conv_std_logic_vector(137, 8),
40163 => conv_std_logic_vector(138, 8),
40164 => conv_std_logic_vector(138, 8),
40165 => conv_std_logic_vector(139, 8),
40166 => conv_std_logic_vector(140, 8),
40167 => conv_std_logic_vector(140, 8),
40168 => conv_std_logic_vector(141, 8),
40169 => conv_std_logic_vector(141, 8),
40170 => conv_std_logic_vector(142, 8),
40171 => conv_std_logic_vector(143, 8),
40172 => conv_std_logic_vector(143, 8),
40173 => conv_std_logic_vector(144, 8),
40174 => conv_std_logic_vector(145, 8),
40175 => conv_std_logic_vector(145, 8),
40176 => conv_std_logic_vector(146, 8),
40177 => conv_std_logic_vector(146, 8),
40178 => conv_std_logic_vector(147, 8),
40179 => conv_std_logic_vector(148, 8),
40180 => conv_std_logic_vector(148, 8),
40181 => conv_std_logic_vector(149, 8),
40182 => conv_std_logic_vector(149, 8),
40183 => conv_std_logic_vector(150, 8),
40184 => conv_std_logic_vector(151, 8),
40185 => conv_std_logic_vector(151, 8),
40186 => conv_std_logic_vector(152, 8),
40187 => conv_std_logic_vector(152, 8),
40188 => conv_std_logic_vector(153, 8),
40189 => conv_std_logic_vector(154, 8),
40190 => conv_std_logic_vector(154, 8),
40191 => conv_std_logic_vector(155, 8),
40192 => conv_std_logic_vector(0, 8),
40193 => conv_std_logic_vector(0, 8),
40194 => conv_std_logic_vector(1, 8),
40195 => conv_std_logic_vector(1, 8),
40196 => conv_std_logic_vector(2, 8),
40197 => conv_std_logic_vector(3, 8),
40198 => conv_std_logic_vector(3, 8),
40199 => conv_std_logic_vector(4, 8),
40200 => conv_std_logic_vector(4, 8),
40201 => conv_std_logic_vector(5, 8),
40202 => conv_std_logic_vector(6, 8),
40203 => conv_std_logic_vector(6, 8),
40204 => conv_std_logic_vector(7, 8),
40205 => conv_std_logic_vector(7, 8),
40206 => conv_std_logic_vector(8, 8),
40207 => conv_std_logic_vector(9, 8),
40208 => conv_std_logic_vector(9, 8),
40209 => conv_std_logic_vector(10, 8),
40210 => conv_std_logic_vector(11, 8),
40211 => conv_std_logic_vector(11, 8),
40212 => conv_std_logic_vector(12, 8),
40213 => conv_std_logic_vector(12, 8),
40214 => conv_std_logic_vector(13, 8),
40215 => conv_std_logic_vector(14, 8),
40216 => conv_std_logic_vector(14, 8),
40217 => conv_std_logic_vector(15, 8),
40218 => conv_std_logic_vector(15, 8),
40219 => conv_std_logic_vector(16, 8),
40220 => conv_std_logic_vector(17, 8),
40221 => conv_std_logic_vector(17, 8),
40222 => conv_std_logic_vector(18, 8),
40223 => conv_std_logic_vector(19, 8),
40224 => conv_std_logic_vector(19, 8),
40225 => conv_std_logic_vector(20, 8),
40226 => conv_std_logic_vector(20, 8),
40227 => conv_std_logic_vector(21, 8),
40228 => conv_std_logic_vector(22, 8),
40229 => conv_std_logic_vector(22, 8),
40230 => conv_std_logic_vector(23, 8),
40231 => conv_std_logic_vector(23, 8),
40232 => conv_std_logic_vector(24, 8),
40233 => conv_std_logic_vector(25, 8),
40234 => conv_std_logic_vector(25, 8),
40235 => conv_std_logic_vector(26, 8),
40236 => conv_std_logic_vector(26, 8),
40237 => conv_std_logic_vector(27, 8),
40238 => conv_std_logic_vector(28, 8),
40239 => conv_std_logic_vector(28, 8),
40240 => conv_std_logic_vector(29, 8),
40241 => conv_std_logic_vector(30, 8),
40242 => conv_std_logic_vector(30, 8),
40243 => conv_std_logic_vector(31, 8),
40244 => conv_std_logic_vector(31, 8),
40245 => conv_std_logic_vector(32, 8),
40246 => conv_std_logic_vector(33, 8),
40247 => conv_std_logic_vector(33, 8),
40248 => conv_std_logic_vector(34, 8),
40249 => conv_std_logic_vector(34, 8),
40250 => conv_std_logic_vector(35, 8),
40251 => conv_std_logic_vector(36, 8),
40252 => conv_std_logic_vector(36, 8),
40253 => conv_std_logic_vector(37, 8),
40254 => conv_std_logic_vector(38, 8),
40255 => conv_std_logic_vector(38, 8),
40256 => conv_std_logic_vector(39, 8),
40257 => conv_std_logic_vector(39, 8),
40258 => conv_std_logic_vector(40, 8),
40259 => conv_std_logic_vector(41, 8),
40260 => conv_std_logic_vector(41, 8),
40261 => conv_std_logic_vector(42, 8),
40262 => conv_std_logic_vector(42, 8),
40263 => conv_std_logic_vector(43, 8),
40264 => conv_std_logic_vector(44, 8),
40265 => conv_std_logic_vector(44, 8),
40266 => conv_std_logic_vector(45, 8),
40267 => conv_std_logic_vector(45, 8),
40268 => conv_std_logic_vector(46, 8),
40269 => conv_std_logic_vector(47, 8),
40270 => conv_std_logic_vector(47, 8),
40271 => conv_std_logic_vector(48, 8),
40272 => conv_std_logic_vector(49, 8),
40273 => conv_std_logic_vector(49, 8),
40274 => conv_std_logic_vector(50, 8),
40275 => conv_std_logic_vector(50, 8),
40276 => conv_std_logic_vector(51, 8),
40277 => conv_std_logic_vector(52, 8),
40278 => conv_std_logic_vector(52, 8),
40279 => conv_std_logic_vector(53, 8),
40280 => conv_std_logic_vector(53, 8),
40281 => conv_std_logic_vector(54, 8),
40282 => conv_std_logic_vector(55, 8),
40283 => conv_std_logic_vector(55, 8),
40284 => conv_std_logic_vector(56, 8),
40285 => conv_std_logic_vector(57, 8),
40286 => conv_std_logic_vector(57, 8),
40287 => conv_std_logic_vector(58, 8),
40288 => conv_std_logic_vector(58, 8),
40289 => conv_std_logic_vector(59, 8),
40290 => conv_std_logic_vector(60, 8),
40291 => conv_std_logic_vector(60, 8),
40292 => conv_std_logic_vector(61, 8),
40293 => conv_std_logic_vector(61, 8),
40294 => conv_std_logic_vector(62, 8),
40295 => conv_std_logic_vector(63, 8),
40296 => conv_std_logic_vector(63, 8),
40297 => conv_std_logic_vector(64, 8),
40298 => conv_std_logic_vector(65, 8),
40299 => conv_std_logic_vector(65, 8),
40300 => conv_std_logic_vector(66, 8),
40301 => conv_std_logic_vector(66, 8),
40302 => conv_std_logic_vector(67, 8),
40303 => conv_std_logic_vector(68, 8),
40304 => conv_std_logic_vector(68, 8),
40305 => conv_std_logic_vector(69, 8),
40306 => conv_std_logic_vector(69, 8),
40307 => conv_std_logic_vector(70, 8),
40308 => conv_std_logic_vector(71, 8),
40309 => conv_std_logic_vector(71, 8),
40310 => conv_std_logic_vector(72, 8),
40311 => conv_std_logic_vector(72, 8),
40312 => conv_std_logic_vector(73, 8),
40313 => conv_std_logic_vector(74, 8),
40314 => conv_std_logic_vector(74, 8),
40315 => conv_std_logic_vector(75, 8),
40316 => conv_std_logic_vector(76, 8),
40317 => conv_std_logic_vector(76, 8),
40318 => conv_std_logic_vector(77, 8),
40319 => conv_std_logic_vector(77, 8),
40320 => conv_std_logic_vector(78, 8),
40321 => conv_std_logic_vector(79, 8),
40322 => conv_std_logic_vector(79, 8),
40323 => conv_std_logic_vector(80, 8),
40324 => conv_std_logic_vector(80, 8),
40325 => conv_std_logic_vector(81, 8),
40326 => conv_std_logic_vector(82, 8),
40327 => conv_std_logic_vector(82, 8),
40328 => conv_std_logic_vector(83, 8),
40329 => conv_std_logic_vector(84, 8),
40330 => conv_std_logic_vector(84, 8),
40331 => conv_std_logic_vector(85, 8),
40332 => conv_std_logic_vector(85, 8),
40333 => conv_std_logic_vector(86, 8),
40334 => conv_std_logic_vector(87, 8),
40335 => conv_std_logic_vector(87, 8),
40336 => conv_std_logic_vector(88, 8),
40337 => conv_std_logic_vector(88, 8),
40338 => conv_std_logic_vector(89, 8),
40339 => conv_std_logic_vector(90, 8),
40340 => conv_std_logic_vector(90, 8),
40341 => conv_std_logic_vector(91, 8),
40342 => conv_std_logic_vector(91, 8),
40343 => conv_std_logic_vector(92, 8),
40344 => conv_std_logic_vector(93, 8),
40345 => conv_std_logic_vector(93, 8),
40346 => conv_std_logic_vector(94, 8),
40347 => conv_std_logic_vector(95, 8),
40348 => conv_std_logic_vector(95, 8),
40349 => conv_std_logic_vector(96, 8),
40350 => conv_std_logic_vector(96, 8),
40351 => conv_std_logic_vector(97, 8),
40352 => conv_std_logic_vector(98, 8),
40353 => conv_std_logic_vector(98, 8),
40354 => conv_std_logic_vector(99, 8),
40355 => conv_std_logic_vector(99, 8),
40356 => conv_std_logic_vector(100, 8),
40357 => conv_std_logic_vector(101, 8),
40358 => conv_std_logic_vector(101, 8),
40359 => conv_std_logic_vector(102, 8),
40360 => conv_std_logic_vector(103, 8),
40361 => conv_std_logic_vector(103, 8),
40362 => conv_std_logic_vector(104, 8),
40363 => conv_std_logic_vector(104, 8),
40364 => conv_std_logic_vector(105, 8),
40365 => conv_std_logic_vector(106, 8),
40366 => conv_std_logic_vector(106, 8),
40367 => conv_std_logic_vector(107, 8),
40368 => conv_std_logic_vector(107, 8),
40369 => conv_std_logic_vector(108, 8),
40370 => conv_std_logic_vector(109, 8),
40371 => conv_std_logic_vector(109, 8),
40372 => conv_std_logic_vector(110, 8),
40373 => conv_std_logic_vector(111, 8),
40374 => conv_std_logic_vector(111, 8),
40375 => conv_std_logic_vector(112, 8),
40376 => conv_std_logic_vector(112, 8),
40377 => conv_std_logic_vector(113, 8),
40378 => conv_std_logic_vector(114, 8),
40379 => conv_std_logic_vector(114, 8),
40380 => conv_std_logic_vector(115, 8),
40381 => conv_std_logic_vector(115, 8),
40382 => conv_std_logic_vector(116, 8),
40383 => conv_std_logic_vector(117, 8),
40384 => conv_std_logic_vector(117, 8),
40385 => conv_std_logic_vector(118, 8),
40386 => conv_std_logic_vector(118, 8),
40387 => conv_std_logic_vector(119, 8),
40388 => conv_std_logic_vector(120, 8),
40389 => conv_std_logic_vector(120, 8),
40390 => conv_std_logic_vector(121, 8),
40391 => conv_std_logic_vector(122, 8),
40392 => conv_std_logic_vector(122, 8),
40393 => conv_std_logic_vector(123, 8),
40394 => conv_std_logic_vector(123, 8),
40395 => conv_std_logic_vector(124, 8),
40396 => conv_std_logic_vector(125, 8),
40397 => conv_std_logic_vector(125, 8),
40398 => conv_std_logic_vector(126, 8),
40399 => conv_std_logic_vector(126, 8),
40400 => conv_std_logic_vector(127, 8),
40401 => conv_std_logic_vector(128, 8),
40402 => conv_std_logic_vector(128, 8),
40403 => conv_std_logic_vector(129, 8),
40404 => conv_std_logic_vector(130, 8),
40405 => conv_std_logic_vector(130, 8),
40406 => conv_std_logic_vector(131, 8),
40407 => conv_std_logic_vector(131, 8),
40408 => conv_std_logic_vector(132, 8),
40409 => conv_std_logic_vector(133, 8),
40410 => conv_std_logic_vector(133, 8),
40411 => conv_std_logic_vector(134, 8),
40412 => conv_std_logic_vector(134, 8),
40413 => conv_std_logic_vector(135, 8),
40414 => conv_std_logic_vector(136, 8),
40415 => conv_std_logic_vector(136, 8),
40416 => conv_std_logic_vector(137, 8),
40417 => conv_std_logic_vector(137, 8),
40418 => conv_std_logic_vector(138, 8),
40419 => conv_std_logic_vector(139, 8),
40420 => conv_std_logic_vector(139, 8),
40421 => conv_std_logic_vector(140, 8),
40422 => conv_std_logic_vector(141, 8),
40423 => conv_std_logic_vector(141, 8),
40424 => conv_std_logic_vector(142, 8),
40425 => conv_std_logic_vector(142, 8),
40426 => conv_std_logic_vector(143, 8),
40427 => conv_std_logic_vector(144, 8),
40428 => conv_std_logic_vector(144, 8),
40429 => conv_std_logic_vector(145, 8),
40430 => conv_std_logic_vector(145, 8),
40431 => conv_std_logic_vector(146, 8),
40432 => conv_std_logic_vector(147, 8),
40433 => conv_std_logic_vector(147, 8),
40434 => conv_std_logic_vector(148, 8),
40435 => conv_std_logic_vector(149, 8),
40436 => conv_std_logic_vector(149, 8),
40437 => conv_std_logic_vector(150, 8),
40438 => conv_std_logic_vector(150, 8),
40439 => conv_std_logic_vector(151, 8),
40440 => conv_std_logic_vector(152, 8),
40441 => conv_std_logic_vector(152, 8),
40442 => conv_std_logic_vector(153, 8),
40443 => conv_std_logic_vector(153, 8),
40444 => conv_std_logic_vector(154, 8),
40445 => conv_std_logic_vector(155, 8),
40446 => conv_std_logic_vector(155, 8),
40447 => conv_std_logic_vector(156, 8),
40448 => conv_std_logic_vector(0, 8),
40449 => conv_std_logic_vector(0, 8),
40450 => conv_std_logic_vector(1, 8),
40451 => conv_std_logic_vector(1, 8),
40452 => conv_std_logic_vector(2, 8),
40453 => conv_std_logic_vector(3, 8),
40454 => conv_std_logic_vector(3, 8),
40455 => conv_std_logic_vector(4, 8),
40456 => conv_std_logic_vector(4, 8),
40457 => conv_std_logic_vector(5, 8),
40458 => conv_std_logic_vector(6, 8),
40459 => conv_std_logic_vector(6, 8),
40460 => conv_std_logic_vector(7, 8),
40461 => conv_std_logic_vector(8, 8),
40462 => conv_std_logic_vector(8, 8),
40463 => conv_std_logic_vector(9, 8),
40464 => conv_std_logic_vector(9, 8),
40465 => conv_std_logic_vector(10, 8),
40466 => conv_std_logic_vector(11, 8),
40467 => conv_std_logic_vector(11, 8),
40468 => conv_std_logic_vector(12, 8),
40469 => conv_std_logic_vector(12, 8),
40470 => conv_std_logic_vector(13, 8),
40471 => conv_std_logic_vector(14, 8),
40472 => conv_std_logic_vector(14, 8),
40473 => conv_std_logic_vector(15, 8),
40474 => conv_std_logic_vector(16, 8),
40475 => conv_std_logic_vector(16, 8),
40476 => conv_std_logic_vector(17, 8),
40477 => conv_std_logic_vector(17, 8),
40478 => conv_std_logic_vector(18, 8),
40479 => conv_std_logic_vector(19, 8),
40480 => conv_std_logic_vector(19, 8),
40481 => conv_std_logic_vector(20, 8),
40482 => conv_std_logic_vector(20, 8),
40483 => conv_std_logic_vector(21, 8),
40484 => conv_std_logic_vector(22, 8),
40485 => conv_std_logic_vector(22, 8),
40486 => conv_std_logic_vector(23, 8),
40487 => conv_std_logic_vector(24, 8),
40488 => conv_std_logic_vector(24, 8),
40489 => conv_std_logic_vector(25, 8),
40490 => conv_std_logic_vector(25, 8),
40491 => conv_std_logic_vector(26, 8),
40492 => conv_std_logic_vector(27, 8),
40493 => conv_std_logic_vector(27, 8),
40494 => conv_std_logic_vector(28, 8),
40495 => conv_std_logic_vector(29, 8),
40496 => conv_std_logic_vector(29, 8),
40497 => conv_std_logic_vector(30, 8),
40498 => conv_std_logic_vector(30, 8),
40499 => conv_std_logic_vector(31, 8),
40500 => conv_std_logic_vector(32, 8),
40501 => conv_std_logic_vector(32, 8),
40502 => conv_std_logic_vector(33, 8),
40503 => conv_std_logic_vector(33, 8),
40504 => conv_std_logic_vector(34, 8),
40505 => conv_std_logic_vector(35, 8),
40506 => conv_std_logic_vector(35, 8),
40507 => conv_std_logic_vector(36, 8),
40508 => conv_std_logic_vector(37, 8),
40509 => conv_std_logic_vector(37, 8),
40510 => conv_std_logic_vector(38, 8),
40511 => conv_std_logic_vector(38, 8),
40512 => conv_std_logic_vector(39, 8),
40513 => conv_std_logic_vector(40, 8),
40514 => conv_std_logic_vector(40, 8),
40515 => conv_std_logic_vector(41, 8),
40516 => conv_std_logic_vector(41, 8),
40517 => conv_std_logic_vector(42, 8),
40518 => conv_std_logic_vector(43, 8),
40519 => conv_std_logic_vector(43, 8),
40520 => conv_std_logic_vector(44, 8),
40521 => conv_std_logic_vector(45, 8),
40522 => conv_std_logic_vector(45, 8),
40523 => conv_std_logic_vector(46, 8),
40524 => conv_std_logic_vector(46, 8),
40525 => conv_std_logic_vector(47, 8),
40526 => conv_std_logic_vector(48, 8),
40527 => conv_std_logic_vector(48, 8),
40528 => conv_std_logic_vector(49, 8),
40529 => conv_std_logic_vector(49, 8),
40530 => conv_std_logic_vector(50, 8),
40531 => conv_std_logic_vector(51, 8),
40532 => conv_std_logic_vector(51, 8),
40533 => conv_std_logic_vector(52, 8),
40534 => conv_std_logic_vector(53, 8),
40535 => conv_std_logic_vector(53, 8),
40536 => conv_std_logic_vector(54, 8),
40537 => conv_std_logic_vector(54, 8),
40538 => conv_std_logic_vector(55, 8),
40539 => conv_std_logic_vector(56, 8),
40540 => conv_std_logic_vector(56, 8),
40541 => conv_std_logic_vector(57, 8),
40542 => conv_std_logic_vector(58, 8),
40543 => conv_std_logic_vector(58, 8),
40544 => conv_std_logic_vector(59, 8),
40545 => conv_std_logic_vector(59, 8),
40546 => conv_std_logic_vector(60, 8),
40547 => conv_std_logic_vector(61, 8),
40548 => conv_std_logic_vector(61, 8),
40549 => conv_std_logic_vector(62, 8),
40550 => conv_std_logic_vector(62, 8),
40551 => conv_std_logic_vector(63, 8),
40552 => conv_std_logic_vector(64, 8),
40553 => conv_std_logic_vector(64, 8),
40554 => conv_std_logic_vector(65, 8),
40555 => conv_std_logic_vector(66, 8),
40556 => conv_std_logic_vector(66, 8),
40557 => conv_std_logic_vector(67, 8),
40558 => conv_std_logic_vector(67, 8),
40559 => conv_std_logic_vector(68, 8),
40560 => conv_std_logic_vector(69, 8),
40561 => conv_std_logic_vector(69, 8),
40562 => conv_std_logic_vector(70, 8),
40563 => conv_std_logic_vector(70, 8),
40564 => conv_std_logic_vector(71, 8),
40565 => conv_std_logic_vector(72, 8),
40566 => conv_std_logic_vector(72, 8),
40567 => conv_std_logic_vector(73, 8),
40568 => conv_std_logic_vector(74, 8),
40569 => conv_std_logic_vector(74, 8),
40570 => conv_std_logic_vector(75, 8),
40571 => conv_std_logic_vector(75, 8),
40572 => conv_std_logic_vector(76, 8),
40573 => conv_std_logic_vector(77, 8),
40574 => conv_std_logic_vector(77, 8),
40575 => conv_std_logic_vector(78, 8),
40576 => conv_std_logic_vector(79, 8),
40577 => conv_std_logic_vector(79, 8),
40578 => conv_std_logic_vector(80, 8),
40579 => conv_std_logic_vector(80, 8),
40580 => conv_std_logic_vector(81, 8),
40581 => conv_std_logic_vector(82, 8),
40582 => conv_std_logic_vector(82, 8),
40583 => conv_std_logic_vector(83, 8),
40584 => conv_std_logic_vector(83, 8),
40585 => conv_std_logic_vector(84, 8),
40586 => conv_std_logic_vector(85, 8),
40587 => conv_std_logic_vector(85, 8),
40588 => conv_std_logic_vector(86, 8),
40589 => conv_std_logic_vector(87, 8),
40590 => conv_std_logic_vector(87, 8),
40591 => conv_std_logic_vector(88, 8),
40592 => conv_std_logic_vector(88, 8),
40593 => conv_std_logic_vector(89, 8),
40594 => conv_std_logic_vector(90, 8),
40595 => conv_std_logic_vector(90, 8),
40596 => conv_std_logic_vector(91, 8),
40597 => conv_std_logic_vector(91, 8),
40598 => conv_std_logic_vector(92, 8),
40599 => conv_std_logic_vector(93, 8),
40600 => conv_std_logic_vector(93, 8),
40601 => conv_std_logic_vector(94, 8),
40602 => conv_std_logic_vector(95, 8),
40603 => conv_std_logic_vector(95, 8),
40604 => conv_std_logic_vector(96, 8),
40605 => conv_std_logic_vector(96, 8),
40606 => conv_std_logic_vector(97, 8),
40607 => conv_std_logic_vector(98, 8),
40608 => conv_std_logic_vector(98, 8),
40609 => conv_std_logic_vector(99, 8),
40610 => conv_std_logic_vector(99, 8),
40611 => conv_std_logic_vector(100, 8),
40612 => conv_std_logic_vector(101, 8),
40613 => conv_std_logic_vector(101, 8),
40614 => conv_std_logic_vector(102, 8),
40615 => conv_std_logic_vector(103, 8),
40616 => conv_std_logic_vector(103, 8),
40617 => conv_std_logic_vector(104, 8),
40618 => conv_std_logic_vector(104, 8),
40619 => conv_std_logic_vector(105, 8),
40620 => conv_std_logic_vector(106, 8),
40621 => conv_std_logic_vector(106, 8),
40622 => conv_std_logic_vector(107, 8),
40623 => conv_std_logic_vector(108, 8),
40624 => conv_std_logic_vector(108, 8),
40625 => conv_std_logic_vector(109, 8),
40626 => conv_std_logic_vector(109, 8),
40627 => conv_std_logic_vector(110, 8),
40628 => conv_std_logic_vector(111, 8),
40629 => conv_std_logic_vector(111, 8),
40630 => conv_std_logic_vector(112, 8),
40631 => conv_std_logic_vector(112, 8),
40632 => conv_std_logic_vector(113, 8),
40633 => conv_std_logic_vector(114, 8),
40634 => conv_std_logic_vector(114, 8),
40635 => conv_std_logic_vector(115, 8),
40636 => conv_std_logic_vector(116, 8),
40637 => conv_std_logic_vector(116, 8),
40638 => conv_std_logic_vector(117, 8),
40639 => conv_std_logic_vector(117, 8),
40640 => conv_std_logic_vector(118, 8),
40641 => conv_std_logic_vector(119, 8),
40642 => conv_std_logic_vector(119, 8),
40643 => conv_std_logic_vector(120, 8),
40644 => conv_std_logic_vector(120, 8),
40645 => conv_std_logic_vector(121, 8),
40646 => conv_std_logic_vector(122, 8),
40647 => conv_std_logic_vector(122, 8),
40648 => conv_std_logic_vector(123, 8),
40649 => conv_std_logic_vector(124, 8),
40650 => conv_std_logic_vector(124, 8),
40651 => conv_std_logic_vector(125, 8),
40652 => conv_std_logic_vector(125, 8),
40653 => conv_std_logic_vector(126, 8),
40654 => conv_std_logic_vector(127, 8),
40655 => conv_std_logic_vector(127, 8),
40656 => conv_std_logic_vector(128, 8),
40657 => conv_std_logic_vector(128, 8),
40658 => conv_std_logic_vector(129, 8),
40659 => conv_std_logic_vector(130, 8),
40660 => conv_std_logic_vector(130, 8),
40661 => conv_std_logic_vector(131, 8),
40662 => conv_std_logic_vector(132, 8),
40663 => conv_std_logic_vector(132, 8),
40664 => conv_std_logic_vector(133, 8),
40665 => conv_std_logic_vector(133, 8),
40666 => conv_std_logic_vector(134, 8),
40667 => conv_std_logic_vector(135, 8),
40668 => conv_std_logic_vector(135, 8),
40669 => conv_std_logic_vector(136, 8),
40670 => conv_std_logic_vector(137, 8),
40671 => conv_std_logic_vector(137, 8),
40672 => conv_std_logic_vector(138, 8),
40673 => conv_std_logic_vector(138, 8),
40674 => conv_std_logic_vector(139, 8),
40675 => conv_std_logic_vector(140, 8),
40676 => conv_std_logic_vector(140, 8),
40677 => conv_std_logic_vector(141, 8),
40678 => conv_std_logic_vector(141, 8),
40679 => conv_std_logic_vector(142, 8),
40680 => conv_std_logic_vector(143, 8),
40681 => conv_std_logic_vector(143, 8),
40682 => conv_std_logic_vector(144, 8),
40683 => conv_std_logic_vector(145, 8),
40684 => conv_std_logic_vector(145, 8),
40685 => conv_std_logic_vector(146, 8),
40686 => conv_std_logic_vector(146, 8),
40687 => conv_std_logic_vector(147, 8),
40688 => conv_std_logic_vector(148, 8),
40689 => conv_std_logic_vector(148, 8),
40690 => conv_std_logic_vector(149, 8),
40691 => conv_std_logic_vector(149, 8),
40692 => conv_std_logic_vector(150, 8),
40693 => conv_std_logic_vector(151, 8),
40694 => conv_std_logic_vector(151, 8),
40695 => conv_std_logic_vector(152, 8),
40696 => conv_std_logic_vector(153, 8),
40697 => conv_std_logic_vector(153, 8),
40698 => conv_std_logic_vector(154, 8),
40699 => conv_std_logic_vector(154, 8),
40700 => conv_std_logic_vector(155, 8),
40701 => conv_std_logic_vector(156, 8),
40702 => conv_std_logic_vector(156, 8),
40703 => conv_std_logic_vector(157, 8),
40704 => conv_std_logic_vector(0, 8),
40705 => conv_std_logic_vector(0, 8),
40706 => conv_std_logic_vector(1, 8),
40707 => conv_std_logic_vector(1, 8),
40708 => conv_std_logic_vector(2, 8),
40709 => conv_std_logic_vector(3, 8),
40710 => conv_std_logic_vector(3, 8),
40711 => conv_std_logic_vector(4, 8),
40712 => conv_std_logic_vector(4, 8),
40713 => conv_std_logic_vector(5, 8),
40714 => conv_std_logic_vector(6, 8),
40715 => conv_std_logic_vector(6, 8),
40716 => conv_std_logic_vector(7, 8),
40717 => conv_std_logic_vector(8, 8),
40718 => conv_std_logic_vector(8, 8),
40719 => conv_std_logic_vector(9, 8),
40720 => conv_std_logic_vector(9, 8),
40721 => conv_std_logic_vector(10, 8),
40722 => conv_std_logic_vector(11, 8),
40723 => conv_std_logic_vector(11, 8),
40724 => conv_std_logic_vector(12, 8),
40725 => conv_std_logic_vector(13, 8),
40726 => conv_std_logic_vector(13, 8),
40727 => conv_std_logic_vector(14, 8),
40728 => conv_std_logic_vector(14, 8),
40729 => conv_std_logic_vector(15, 8),
40730 => conv_std_logic_vector(16, 8),
40731 => conv_std_logic_vector(16, 8),
40732 => conv_std_logic_vector(17, 8),
40733 => conv_std_logic_vector(18, 8),
40734 => conv_std_logic_vector(18, 8),
40735 => conv_std_logic_vector(19, 8),
40736 => conv_std_logic_vector(19, 8),
40737 => conv_std_logic_vector(20, 8),
40738 => conv_std_logic_vector(21, 8),
40739 => conv_std_logic_vector(21, 8),
40740 => conv_std_logic_vector(22, 8),
40741 => conv_std_logic_vector(22, 8),
40742 => conv_std_logic_vector(23, 8),
40743 => conv_std_logic_vector(24, 8),
40744 => conv_std_logic_vector(24, 8),
40745 => conv_std_logic_vector(25, 8),
40746 => conv_std_logic_vector(26, 8),
40747 => conv_std_logic_vector(26, 8),
40748 => conv_std_logic_vector(27, 8),
40749 => conv_std_logic_vector(27, 8),
40750 => conv_std_logic_vector(28, 8),
40751 => conv_std_logic_vector(29, 8),
40752 => conv_std_logic_vector(29, 8),
40753 => conv_std_logic_vector(30, 8),
40754 => conv_std_logic_vector(31, 8),
40755 => conv_std_logic_vector(31, 8),
40756 => conv_std_logic_vector(32, 8),
40757 => conv_std_logic_vector(32, 8),
40758 => conv_std_logic_vector(33, 8),
40759 => conv_std_logic_vector(34, 8),
40760 => conv_std_logic_vector(34, 8),
40761 => conv_std_logic_vector(35, 8),
40762 => conv_std_logic_vector(36, 8),
40763 => conv_std_logic_vector(36, 8),
40764 => conv_std_logic_vector(37, 8),
40765 => conv_std_logic_vector(37, 8),
40766 => conv_std_logic_vector(38, 8),
40767 => conv_std_logic_vector(39, 8),
40768 => conv_std_logic_vector(39, 8),
40769 => conv_std_logic_vector(40, 8),
40770 => conv_std_logic_vector(40, 8),
40771 => conv_std_logic_vector(41, 8),
40772 => conv_std_logic_vector(42, 8),
40773 => conv_std_logic_vector(42, 8),
40774 => conv_std_logic_vector(43, 8),
40775 => conv_std_logic_vector(44, 8),
40776 => conv_std_logic_vector(44, 8),
40777 => conv_std_logic_vector(45, 8),
40778 => conv_std_logic_vector(45, 8),
40779 => conv_std_logic_vector(46, 8),
40780 => conv_std_logic_vector(47, 8),
40781 => conv_std_logic_vector(47, 8),
40782 => conv_std_logic_vector(48, 8),
40783 => conv_std_logic_vector(49, 8),
40784 => conv_std_logic_vector(49, 8),
40785 => conv_std_logic_vector(50, 8),
40786 => conv_std_logic_vector(50, 8),
40787 => conv_std_logic_vector(51, 8),
40788 => conv_std_logic_vector(52, 8),
40789 => conv_std_logic_vector(52, 8),
40790 => conv_std_logic_vector(53, 8),
40791 => conv_std_logic_vector(54, 8),
40792 => conv_std_logic_vector(54, 8),
40793 => conv_std_logic_vector(55, 8),
40794 => conv_std_logic_vector(55, 8),
40795 => conv_std_logic_vector(56, 8),
40796 => conv_std_logic_vector(57, 8),
40797 => conv_std_logic_vector(57, 8),
40798 => conv_std_logic_vector(58, 8),
40799 => conv_std_logic_vector(59, 8),
40800 => conv_std_logic_vector(59, 8),
40801 => conv_std_logic_vector(60, 8),
40802 => conv_std_logic_vector(60, 8),
40803 => conv_std_logic_vector(61, 8),
40804 => conv_std_logic_vector(62, 8),
40805 => conv_std_logic_vector(62, 8),
40806 => conv_std_logic_vector(63, 8),
40807 => conv_std_logic_vector(63, 8),
40808 => conv_std_logic_vector(64, 8),
40809 => conv_std_logic_vector(65, 8),
40810 => conv_std_logic_vector(65, 8),
40811 => conv_std_logic_vector(66, 8),
40812 => conv_std_logic_vector(67, 8),
40813 => conv_std_logic_vector(67, 8),
40814 => conv_std_logic_vector(68, 8),
40815 => conv_std_logic_vector(68, 8),
40816 => conv_std_logic_vector(69, 8),
40817 => conv_std_logic_vector(70, 8),
40818 => conv_std_logic_vector(70, 8),
40819 => conv_std_logic_vector(71, 8),
40820 => conv_std_logic_vector(72, 8),
40821 => conv_std_logic_vector(72, 8),
40822 => conv_std_logic_vector(73, 8),
40823 => conv_std_logic_vector(73, 8),
40824 => conv_std_logic_vector(74, 8),
40825 => conv_std_logic_vector(75, 8),
40826 => conv_std_logic_vector(75, 8),
40827 => conv_std_logic_vector(76, 8),
40828 => conv_std_logic_vector(77, 8),
40829 => conv_std_logic_vector(77, 8),
40830 => conv_std_logic_vector(78, 8),
40831 => conv_std_logic_vector(78, 8),
40832 => conv_std_logic_vector(79, 8),
40833 => conv_std_logic_vector(80, 8),
40834 => conv_std_logic_vector(80, 8),
40835 => conv_std_logic_vector(81, 8),
40836 => conv_std_logic_vector(81, 8),
40837 => conv_std_logic_vector(82, 8),
40838 => conv_std_logic_vector(83, 8),
40839 => conv_std_logic_vector(83, 8),
40840 => conv_std_logic_vector(84, 8),
40841 => conv_std_logic_vector(85, 8),
40842 => conv_std_logic_vector(85, 8),
40843 => conv_std_logic_vector(86, 8),
40844 => conv_std_logic_vector(86, 8),
40845 => conv_std_logic_vector(87, 8),
40846 => conv_std_logic_vector(88, 8),
40847 => conv_std_logic_vector(88, 8),
40848 => conv_std_logic_vector(89, 8),
40849 => conv_std_logic_vector(90, 8),
40850 => conv_std_logic_vector(90, 8),
40851 => conv_std_logic_vector(91, 8),
40852 => conv_std_logic_vector(91, 8),
40853 => conv_std_logic_vector(92, 8),
40854 => conv_std_logic_vector(93, 8),
40855 => conv_std_logic_vector(93, 8),
40856 => conv_std_logic_vector(94, 8),
40857 => conv_std_logic_vector(95, 8),
40858 => conv_std_logic_vector(95, 8),
40859 => conv_std_logic_vector(96, 8),
40860 => conv_std_logic_vector(96, 8),
40861 => conv_std_logic_vector(97, 8),
40862 => conv_std_logic_vector(98, 8),
40863 => conv_std_logic_vector(98, 8),
40864 => conv_std_logic_vector(99, 8),
40865 => conv_std_logic_vector(99, 8),
40866 => conv_std_logic_vector(100, 8),
40867 => conv_std_logic_vector(101, 8),
40868 => conv_std_logic_vector(101, 8),
40869 => conv_std_logic_vector(102, 8),
40870 => conv_std_logic_vector(103, 8),
40871 => conv_std_logic_vector(103, 8),
40872 => conv_std_logic_vector(104, 8),
40873 => conv_std_logic_vector(104, 8),
40874 => conv_std_logic_vector(105, 8),
40875 => conv_std_logic_vector(106, 8),
40876 => conv_std_logic_vector(106, 8),
40877 => conv_std_logic_vector(107, 8),
40878 => conv_std_logic_vector(108, 8),
40879 => conv_std_logic_vector(108, 8),
40880 => conv_std_logic_vector(109, 8),
40881 => conv_std_logic_vector(109, 8),
40882 => conv_std_logic_vector(110, 8),
40883 => conv_std_logic_vector(111, 8),
40884 => conv_std_logic_vector(111, 8),
40885 => conv_std_logic_vector(112, 8),
40886 => conv_std_logic_vector(113, 8),
40887 => conv_std_logic_vector(113, 8),
40888 => conv_std_logic_vector(114, 8),
40889 => conv_std_logic_vector(114, 8),
40890 => conv_std_logic_vector(115, 8),
40891 => conv_std_logic_vector(116, 8),
40892 => conv_std_logic_vector(116, 8),
40893 => conv_std_logic_vector(117, 8),
40894 => conv_std_logic_vector(118, 8),
40895 => conv_std_logic_vector(118, 8),
40896 => conv_std_logic_vector(119, 8),
40897 => conv_std_logic_vector(119, 8),
40898 => conv_std_logic_vector(120, 8),
40899 => conv_std_logic_vector(121, 8),
40900 => conv_std_logic_vector(121, 8),
40901 => conv_std_logic_vector(122, 8),
40902 => conv_std_logic_vector(122, 8),
40903 => conv_std_logic_vector(123, 8),
40904 => conv_std_logic_vector(124, 8),
40905 => conv_std_logic_vector(124, 8),
40906 => conv_std_logic_vector(125, 8),
40907 => conv_std_logic_vector(126, 8),
40908 => conv_std_logic_vector(126, 8),
40909 => conv_std_logic_vector(127, 8),
40910 => conv_std_logic_vector(127, 8),
40911 => conv_std_logic_vector(128, 8),
40912 => conv_std_logic_vector(129, 8),
40913 => conv_std_logic_vector(129, 8),
40914 => conv_std_logic_vector(130, 8),
40915 => conv_std_logic_vector(131, 8),
40916 => conv_std_logic_vector(131, 8),
40917 => conv_std_logic_vector(132, 8),
40918 => conv_std_logic_vector(132, 8),
40919 => conv_std_logic_vector(133, 8),
40920 => conv_std_logic_vector(134, 8),
40921 => conv_std_logic_vector(134, 8),
40922 => conv_std_logic_vector(135, 8),
40923 => conv_std_logic_vector(136, 8),
40924 => conv_std_logic_vector(136, 8),
40925 => conv_std_logic_vector(137, 8),
40926 => conv_std_logic_vector(137, 8),
40927 => conv_std_logic_vector(138, 8),
40928 => conv_std_logic_vector(139, 8),
40929 => conv_std_logic_vector(139, 8),
40930 => conv_std_logic_vector(140, 8),
40931 => conv_std_logic_vector(140, 8),
40932 => conv_std_logic_vector(141, 8),
40933 => conv_std_logic_vector(142, 8),
40934 => conv_std_logic_vector(142, 8),
40935 => conv_std_logic_vector(143, 8),
40936 => conv_std_logic_vector(144, 8),
40937 => conv_std_logic_vector(144, 8),
40938 => conv_std_logic_vector(145, 8),
40939 => conv_std_logic_vector(145, 8),
40940 => conv_std_logic_vector(146, 8),
40941 => conv_std_logic_vector(147, 8),
40942 => conv_std_logic_vector(147, 8),
40943 => conv_std_logic_vector(148, 8),
40944 => conv_std_logic_vector(149, 8),
40945 => conv_std_logic_vector(149, 8),
40946 => conv_std_logic_vector(150, 8),
40947 => conv_std_logic_vector(150, 8),
40948 => conv_std_logic_vector(151, 8),
40949 => conv_std_logic_vector(152, 8),
40950 => conv_std_logic_vector(152, 8),
40951 => conv_std_logic_vector(153, 8),
40952 => conv_std_logic_vector(154, 8),
40953 => conv_std_logic_vector(154, 8),
40954 => conv_std_logic_vector(155, 8),
40955 => conv_std_logic_vector(155, 8),
40956 => conv_std_logic_vector(156, 8),
40957 => conv_std_logic_vector(157, 8),
40958 => conv_std_logic_vector(157, 8),
40959 => conv_std_logic_vector(158, 8),
40960 => conv_std_logic_vector(0, 8),
40961 => conv_std_logic_vector(0, 8),
40962 => conv_std_logic_vector(1, 8),
40963 => conv_std_logic_vector(1, 8),
40964 => conv_std_logic_vector(2, 8),
40965 => conv_std_logic_vector(3, 8),
40966 => conv_std_logic_vector(3, 8),
40967 => conv_std_logic_vector(4, 8),
40968 => conv_std_logic_vector(5, 8),
40969 => conv_std_logic_vector(5, 8),
40970 => conv_std_logic_vector(6, 8),
40971 => conv_std_logic_vector(6, 8),
40972 => conv_std_logic_vector(7, 8),
40973 => conv_std_logic_vector(8, 8),
40974 => conv_std_logic_vector(8, 8),
40975 => conv_std_logic_vector(9, 8),
40976 => conv_std_logic_vector(10, 8),
40977 => conv_std_logic_vector(10, 8),
40978 => conv_std_logic_vector(11, 8),
40979 => conv_std_logic_vector(11, 8),
40980 => conv_std_logic_vector(12, 8),
40981 => conv_std_logic_vector(13, 8),
40982 => conv_std_logic_vector(13, 8),
40983 => conv_std_logic_vector(14, 8),
40984 => conv_std_logic_vector(15, 8),
40985 => conv_std_logic_vector(15, 8),
40986 => conv_std_logic_vector(16, 8),
40987 => conv_std_logic_vector(16, 8),
40988 => conv_std_logic_vector(17, 8),
40989 => conv_std_logic_vector(18, 8),
40990 => conv_std_logic_vector(18, 8),
40991 => conv_std_logic_vector(19, 8),
40992 => conv_std_logic_vector(20, 8),
40993 => conv_std_logic_vector(20, 8),
40994 => conv_std_logic_vector(21, 8),
40995 => conv_std_logic_vector(21, 8),
40996 => conv_std_logic_vector(22, 8),
40997 => conv_std_logic_vector(23, 8),
40998 => conv_std_logic_vector(23, 8),
40999 => conv_std_logic_vector(24, 8),
41000 => conv_std_logic_vector(25, 8),
41001 => conv_std_logic_vector(25, 8),
41002 => conv_std_logic_vector(26, 8),
41003 => conv_std_logic_vector(26, 8),
41004 => conv_std_logic_vector(27, 8),
41005 => conv_std_logic_vector(28, 8),
41006 => conv_std_logic_vector(28, 8),
41007 => conv_std_logic_vector(29, 8),
41008 => conv_std_logic_vector(30, 8),
41009 => conv_std_logic_vector(30, 8),
41010 => conv_std_logic_vector(31, 8),
41011 => conv_std_logic_vector(31, 8),
41012 => conv_std_logic_vector(32, 8),
41013 => conv_std_logic_vector(33, 8),
41014 => conv_std_logic_vector(33, 8),
41015 => conv_std_logic_vector(34, 8),
41016 => conv_std_logic_vector(35, 8),
41017 => conv_std_logic_vector(35, 8),
41018 => conv_std_logic_vector(36, 8),
41019 => conv_std_logic_vector(36, 8),
41020 => conv_std_logic_vector(37, 8),
41021 => conv_std_logic_vector(38, 8),
41022 => conv_std_logic_vector(38, 8),
41023 => conv_std_logic_vector(39, 8),
41024 => conv_std_logic_vector(40, 8),
41025 => conv_std_logic_vector(40, 8),
41026 => conv_std_logic_vector(41, 8),
41027 => conv_std_logic_vector(41, 8),
41028 => conv_std_logic_vector(42, 8),
41029 => conv_std_logic_vector(43, 8),
41030 => conv_std_logic_vector(43, 8),
41031 => conv_std_logic_vector(44, 8),
41032 => conv_std_logic_vector(45, 8),
41033 => conv_std_logic_vector(45, 8),
41034 => conv_std_logic_vector(46, 8),
41035 => conv_std_logic_vector(46, 8),
41036 => conv_std_logic_vector(47, 8),
41037 => conv_std_logic_vector(48, 8),
41038 => conv_std_logic_vector(48, 8),
41039 => conv_std_logic_vector(49, 8),
41040 => conv_std_logic_vector(50, 8),
41041 => conv_std_logic_vector(50, 8),
41042 => conv_std_logic_vector(51, 8),
41043 => conv_std_logic_vector(51, 8),
41044 => conv_std_logic_vector(52, 8),
41045 => conv_std_logic_vector(53, 8),
41046 => conv_std_logic_vector(53, 8),
41047 => conv_std_logic_vector(54, 8),
41048 => conv_std_logic_vector(55, 8),
41049 => conv_std_logic_vector(55, 8),
41050 => conv_std_logic_vector(56, 8),
41051 => conv_std_logic_vector(56, 8),
41052 => conv_std_logic_vector(57, 8),
41053 => conv_std_logic_vector(58, 8),
41054 => conv_std_logic_vector(58, 8),
41055 => conv_std_logic_vector(59, 8),
41056 => conv_std_logic_vector(60, 8),
41057 => conv_std_logic_vector(60, 8),
41058 => conv_std_logic_vector(61, 8),
41059 => conv_std_logic_vector(61, 8),
41060 => conv_std_logic_vector(62, 8),
41061 => conv_std_logic_vector(63, 8),
41062 => conv_std_logic_vector(63, 8),
41063 => conv_std_logic_vector(64, 8),
41064 => conv_std_logic_vector(65, 8),
41065 => conv_std_logic_vector(65, 8),
41066 => conv_std_logic_vector(66, 8),
41067 => conv_std_logic_vector(66, 8),
41068 => conv_std_logic_vector(67, 8),
41069 => conv_std_logic_vector(68, 8),
41070 => conv_std_logic_vector(68, 8),
41071 => conv_std_logic_vector(69, 8),
41072 => conv_std_logic_vector(70, 8),
41073 => conv_std_logic_vector(70, 8),
41074 => conv_std_logic_vector(71, 8),
41075 => conv_std_logic_vector(71, 8),
41076 => conv_std_logic_vector(72, 8),
41077 => conv_std_logic_vector(73, 8),
41078 => conv_std_logic_vector(73, 8),
41079 => conv_std_logic_vector(74, 8),
41080 => conv_std_logic_vector(75, 8),
41081 => conv_std_logic_vector(75, 8),
41082 => conv_std_logic_vector(76, 8),
41083 => conv_std_logic_vector(76, 8),
41084 => conv_std_logic_vector(77, 8),
41085 => conv_std_logic_vector(78, 8),
41086 => conv_std_logic_vector(78, 8),
41087 => conv_std_logic_vector(79, 8),
41088 => conv_std_logic_vector(80, 8),
41089 => conv_std_logic_vector(80, 8),
41090 => conv_std_logic_vector(81, 8),
41091 => conv_std_logic_vector(81, 8),
41092 => conv_std_logic_vector(82, 8),
41093 => conv_std_logic_vector(83, 8),
41094 => conv_std_logic_vector(83, 8),
41095 => conv_std_logic_vector(84, 8),
41096 => conv_std_logic_vector(85, 8),
41097 => conv_std_logic_vector(85, 8),
41098 => conv_std_logic_vector(86, 8),
41099 => conv_std_logic_vector(86, 8),
41100 => conv_std_logic_vector(87, 8),
41101 => conv_std_logic_vector(88, 8),
41102 => conv_std_logic_vector(88, 8),
41103 => conv_std_logic_vector(89, 8),
41104 => conv_std_logic_vector(90, 8),
41105 => conv_std_logic_vector(90, 8),
41106 => conv_std_logic_vector(91, 8),
41107 => conv_std_logic_vector(91, 8),
41108 => conv_std_logic_vector(92, 8),
41109 => conv_std_logic_vector(93, 8),
41110 => conv_std_logic_vector(93, 8),
41111 => conv_std_logic_vector(94, 8),
41112 => conv_std_logic_vector(95, 8),
41113 => conv_std_logic_vector(95, 8),
41114 => conv_std_logic_vector(96, 8),
41115 => conv_std_logic_vector(96, 8),
41116 => conv_std_logic_vector(97, 8),
41117 => conv_std_logic_vector(98, 8),
41118 => conv_std_logic_vector(98, 8),
41119 => conv_std_logic_vector(99, 8),
41120 => conv_std_logic_vector(100, 8),
41121 => conv_std_logic_vector(100, 8),
41122 => conv_std_logic_vector(101, 8),
41123 => conv_std_logic_vector(101, 8),
41124 => conv_std_logic_vector(102, 8),
41125 => conv_std_logic_vector(103, 8),
41126 => conv_std_logic_vector(103, 8),
41127 => conv_std_logic_vector(104, 8),
41128 => conv_std_logic_vector(105, 8),
41129 => conv_std_logic_vector(105, 8),
41130 => conv_std_logic_vector(106, 8),
41131 => conv_std_logic_vector(106, 8),
41132 => conv_std_logic_vector(107, 8),
41133 => conv_std_logic_vector(108, 8),
41134 => conv_std_logic_vector(108, 8),
41135 => conv_std_logic_vector(109, 8),
41136 => conv_std_logic_vector(110, 8),
41137 => conv_std_logic_vector(110, 8),
41138 => conv_std_logic_vector(111, 8),
41139 => conv_std_logic_vector(111, 8),
41140 => conv_std_logic_vector(112, 8),
41141 => conv_std_logic_vector(113, 8),
41142 => conv_std_logic_vector(113, 8),
41143 => conv_std_logic_vector(114, 8),
41144 => conv_std_logic_vector(115, 8),
41145 => conv_std_logic_vector(115, 8),
41146 => conv_std_logic_vector(116, 8),
41147 => conv_std_logic_vector(116, 8),
41148 => conv_std_logic_vector(117, 8),
41149 => conv_std_logic_vector(118, 8),
41150 => conv_std_logic_vector(118, 8),
41151 => conv_std_logic_vector(119, 8),
41152 => conv_std_logic_vector(120, 8),
41153 => conv_std_logic_vector(120, 8),
41154 => conv_std_logic_vector(121, 8),
41155 => conv_std_logic_vector(121, 8),
41156 => conv_std_logic_vector(122, 8),
41157 => conv_std_logic_vector(123, 8),
41158 => conv_std_logic_vector(123, 8),
41159 => conv_std_logic_vector(124, 8),
41160 => conv_std_logic_vector(125, 8),
41161 => conv_std_logic_vector(125, 8),
41162 => conv_std_logic_vector(126, 8),
41163 => conv_std_logic_vector(126, 8),
41164 => conv_std_logic_vector(127, 8),
41165 => conv_std_logic_vector(128, 8),
41166 => conv_std_logic_vector(128, 8),
41167 => conv_std_logic_vector(129, 8),
41168 => conv_std_logic_vector(130, 8),
41169 => conv_std_logic_vector(130, 8),
41170 => conv_std_logic_vector(131, 8),
41171 => conv_std_logic_vector(131, 8),
41172 => conv_std_logic_vector(132, 8),
41173 => conv_std_logic_vector(133, 8),
41174 => conv_std_logic_vector(133, 8),
41175 => conv_std_logic_vector(134, 8),
41176 => conv_std_logic_vector(135, 8),
41177 => conv_std_logic_vector(135, 8),
41178 => conv_std_logic_vector(136, 8),
41179 => conv_std_logic_vector(136, 8),
41180 => conv_std_logic_vector(137, 8),
41181 => conv_std_logic_vector(138, 8),
41182 => conv_std_logic_vector(138, 8),
41183 => conv_std_logic_vector(139, 8),
41184 => conv_std_logic_vector(140, 8),
41185 => conv_std_logic_vector(140, 8),
41186 => conv_std_logic_vector(141, 8),
41187 => conv_std_logic_vector(141, 8),
41188 => conv_std_logic_vector(142, 8),
41189 => conv_std_logic_vector(143, 8),
41190 => conv_std_logic_vector(143, 8),
41191 => conv_std_logic_vector(144, 8),
41192 => conv_std_logic_vector(145, 8),
41193 => conv_std_logic_vector(145, 8),
41194 => conv_std_logic_vector(146, 8),
41195 => conv_std_logic_vector(146, 8),
41196 => conv_std_logic_vector(147, 8),
41197 => conv_std_logic_vector(148, 8),
41198 => conv_std_logic_vector(148, 8),
41199 => conv_std_logic_vector(149, 8),
41200 => conv_std_logic_vector(150, 8),
41201 => conv_std_logic_vector(150, 8),
41202 => conv_std_logic_vector(151, 8),
41203 => conv_std_logic_vector(151, 8),
41204 => conv_std_logic_vector(152, 8),
41205 => conv_std_logic_vector(153, 8),
41206 => conv_std_logic_vector(153, 8),
41207 => conv_std_logic_vector(154, 8),
41208 => conv_std_logic_vector(155, 8),
41209 => conv_std_logic_vector(155, 8),
41210 => conv_std_logic_vector(156, 8),
41211 => conv_std_logic_vector(156, 8),
41212 => conv_std_logic_vector(157, 8),
41213 => conv_std_logic_vector(158, 8),
41214 => conv_std_logic_vector(158, 8),
41215 => conv_std_logic_vector(159, 8),
41216 => conv_std_logic_vector(0, 8),
41217 => conv_std_logic_vector(0, 8),
41218 => conv_std_logic_vector(1, 8),
41219 => conv_std_logic_vector(1, 8),
41220 => conv_std_logic_vector(2, 8),
41221 => conv_std_logic_vector(3, 8),
41222 => conv_std_logic_vector(3, 8),
41223 => conv_std_logic_vector(4, 8),
41224 => conv_std_logic_vector(5, 8),
41225 => conv_std_logic_vector(5, 8),
41226 => conv_std_logic_vector(6, 8),
41227 => conv_std_logic_vector(6, 8),
41228 => conv_std_logic_vector(7, 8),
41229 => conv_std_logic_vector(8, 8),
41230 => conv_std_logic_vector(8, 8),
41231 => conv_std_logic_vector(9, 8),
41232 => conv_std_logic_vector(10, 8),
41233 => conv_std_logic_vector(10, 8),
41234 => conv_std_logic_vector(11, 8),
41235 => conv_std_logic_vector(11, 8),
41236 => conv_std_logic_vector(12, 8),
41237 => conv_std_logic_vector(13, 8),
41238 => conv_std_logic_vector(13, 8),
41239 => conv_std_logic_vector(14, 8),
41240 => conv_std_logic_vector(15, 8),
41241 => conv_std_logic_vector(15, 8),
41242 => conv_std_logic_vector(16, 8),
41243 => conv_std_logic_vector(16, 8),
41244 => conv_std_logic_vector(17, 8),
41245 => conv_std_logic_vector(18, 8),
41246 => conv_std_logic_vector(18, 8),
41247 => conv_std_logic_vector(19, 8),
41248 => conv_std_logic_vector(20, 8),
41249 => conv_std_logic_vector(20, 8),
41250 => conv_std_logic_vector(21, 8),
41251 => conv_std_logic_vector(22, 8),
41252 => conv_std_logic_vector(22, 8),
41253 => conv_std_logic_vector(23, 8),
41254 => conv_std_logic_vector(23, 8),
41255 => conv_std_logic_vector(24, 8),
41256 => conv_std_logic_vector(25, 8),
41257 => conv_std_logic_vector(25, 8),
41258 => conv_std_logic_vector(26, 8),
41259 => conv_std_logic_vector(27, 8),
41260 => conv_std_logic_vector(27, 8),
41261 => conv_std_logic_vector(28, 8),
41262 => conv_std_logic_vector(28, 8),
41263 => conv_std_logic_vector(29, 8),
41264 => conv_std_logic_vector(30, 8),
41265 => conv_std_logic_vector(30, 8),
41266 => conv_std_logic_vector(31, 8),
41267 => conv_std_logic_vector(32, 8),
41268 => conv_std_logic_vector(32, 8),
41269 => conv_std_logic_vector(33, 8),
41270 => conv_std_logic_vector(33, 8),
41271 => conv_std_logic_vector(34, 8),
41272 => conv_std_logic_vector(35, 8),
41273 => conv_std_logic_vector(35, 8),
41274 => conv_std_logic_vector(36, 8),
41275 => conv_std_logic_vector(37, 8),
41276 => conv_std_logic_vector(37, 8),
41277 => conv_std_logic_vector(38, 8),
41278 => conv_std_logic_vector(38, 8),
41279 => conv_std_logic_vector(39, 8),
41280 => conv_std_logic_vector(40, 8),
41281 => conv_std_logic_vector(40, 8),
41282 => conv_std_logic_vector(41, 8),
41283 => conv_std_logic_vector(42, 8),
41284 => conv_std_logic_vector(42, 8),
41285 => conv_std_logic_vector(43, 8),
41286 => conv_std_logic_vector(44, 8),
41287 => conv_std_logic_vector(44, 8),
41288 => conv_std_logic_vector(45, 8),
41289 => conv_std_logic_vector(45, 8),
41290 => conv_std_logic_vector(46, 8),
41291 => conv_std_logic_vector(47, 8),
41292 => conv_std_logic_vector(47, 8),
41293 => conv_std_logic_vector(48, 8),
41294 => conv_std_logic_vector(49, 8),
41295 => conv_std_logic_vector(49, 8),
41296 => conv_std_logic_vector(50, 8),
41297 => conv_std_logic_vector(50, 8),
41298 => conv_std_logic_vector(51, 8),
41299 => conv_std_logic_vector(52, 8),
41300 => conv_std_logic_vector(52, 8),
41301 => conv_std_logic_vector(53, 8),
41302 => conv_std_logic_vector(54, 8),
41303 => conv_std_logic_vector(54, 8),
41304 => conv_std_logic_vector(55, 8),
41305 => conv_std_logic_vector(55, 8),
41306 => conv_std_logic_vector(56, 8),
41307 => conv_std_logic_vector(57, 8),
41308 => conv_std_logic_vector(57, 8),
41309 => conv_std_logic_vector(58, 8),
41310 => conv_std_logic_vector(59, 8),
41311 => conv_std_logic_vector(59, 8),
41312 => conv_std_logic_vector(60, 8),
41313 => conv_std_logic_vector(61, 8),
41314 => conv_std_logic_vector(61, 8),
41315 => conv_std_logic_vector(62, 8),
41316 => conv_std_logic_vector(62, 8),
41317 => conv_std_logic_vector(63, 8),
41318 => conv_std_logic_vector(64, 8),
41319 => conv_std_logic_vector(64, 8),
41320 => conv_std_logic_vector(65, 8),
41321 => conv_std_logic_vector(66, 8),
41322 => conv_std_logic_vector(66, 8),
41323 => conv_std_logic_vector(67, 8),
41324 => conv_std_logic_vector(67, 8),
41325 => conv_std_logic_vector(68, 8),
41326 => conv_std_logic_vector(69, 8),
41327 => conv_std_logic_vector(69, 8),
41328 => conv_std_logic_vector(70, 8),
41329 => conv_std_logic_vector(71, 8),
41330 => conv_std_logic_vector(71, 8),
41331 => conv_std_logic_vector(72, 8),
41332 => conv_std_logic_vector(72, 8),
41333 => conv_std_logic_vector(73, 8),
41334 => conv_std_logic_vector(74, 8),
41335 => conv_std_logic_vector(74, 8),
41336 => conv_std_logic_vector(75, 8),
41337 => conv_std_logic_vector(76, 8),
41338 => conv_std_logic_vector(76, 8),
41339 => conv_std_logic_vector(77, 8),
41340 => conv_std_logic_vector(77, 8),
41341 => conv_std_logic_vector(78, 8),
41342 => conv_std_logic_vector(79, 8),
41343 => conv_std_logic_vector(79, 8),
41344 => conv_std_logic_vector(80, 8),
41345 => conv_std_logic_vector(81, 8),
41346 => conv_std_logic_vector(81, 8),
41347 => conv_std_logic_vector(82, 8),
41348 => conv_std_logic_vector(83, 8),
41349 => conv_std_logic_vector(83, 8),
41350 => conv_std_logic_vector(84, 8),
41351 => conv_std_logic_vector(84, 8),
41352 => conv_std_logic_vector(85, 8),
41353 => conv_std_logic_vector(86, 8),
41354 => conv_std_logic_vector(86, 8),
41355 => conv_std_logic_vector(87, 8),
41356 => conv_std_logic_vector(88, 8),
41357 => conv_std_logic_vector(88, 8),
41358 => conv_std_logic_vector(89, 8),
41359 => conv_std_logic_vector(89, 8),
41360 => conv_std_logic_vector(90, 8),
41361 => conv_std_logic_vector(91, 8),
41362 => conv_std_logic_vector(91, 8),
41363 => conv_std_logic_vector(92, 8),
41364 => conv_std_logic_vector(93, 8),
41365 => conv_std_logic_vector(93, 8),
41366 => conv_std_logic_vector(94, 8),
41367 => conv_std_logic_vector(94, 8),
41368 => conv_std_logic_vector(95, 8),
41369 => conv_std_logic_vector(96, 8),
41370 => conv_std_logic_vector(96, 8),
41371 => conv_std_logic_vector(97, 8),
41372 => conv_std_logic_vector(98, 8),
41373 => conv_std_logic_vector(98, 8),
41374 => conv_std_logic_vector(99, 8),
41375 => conv_std_logic_vector(99, 8),
41376 => conv_std_logic_vector(100, 8),
41377 => conv_std_logic_vector(101, 8),
41378 => conv_std_logic_vector(101, 8),
41379 => conv_std_logic_vector(102, 8),
41380 => conv_std_logic_vector(103, 8),
41381 => conv_std_logic_vector(103, 8),
41382 => conv_std_logic_vector(104, 8),
41383 => conv_std_logic_vector(105, 8),
41384 => conv_std_logic_vector(105, 8),
41385 => conv_std_logic_vector(106, 8),
41386 => conv_std_logic_vector(106, 8),
41387 => conv_std_logic_vector(107, 8),
41388 => conv_std_logic_vector(108, 8),
41389 => conv_std_logic_vector(108, 8),
41390 => conv_std_logic_vector(109, 8),
41391 => conv_std_logic_vector(110, 8),
41392 => conv_std_logic_vector(110, 8),
41393 => conv_std_logic_vector(111, 8),
41394 => conv_std_logic_vector(111, 8),
41395 => conv_std_logic_vector(112, 8),
41396 => conv_std_logic_vector(113, 8),
41397 => conv_std_logic_vector(113, 8),
41398 => conv_std_logic_vector(114, 8),
41399 => conv_std_logic_vector(115, 8),
41400 => conv_std_logic_vector(115, 8),
41401 => conv_std_logic_vector(116, 8),
41402 => conv_std_logic_vector(116, 8),
41403 => conv_std_logic_vector(117, 8),
41404 => conv_std_logic_vector(118, 8),
41405 => conv_std_logic_vector(118, 8),
41406 => conv_std_logic_vector(119, 8),
41407 => conv_std_logic_vector(120, 8),
41408 => conv_std_logic_vector(120, 8),
41409 => conv_std_logic_vector(121, 8),
41410 => conv_std_logic_vector(122, 8),
41411 => conv_std_logic_vector(122, 8),
41412 => conv_std_logic_vector(123, 8),
41413 => conv_std_logic_vector(123, 8),
41414 => conv_std_logic_vector(124, 8),
41415 => conv_std_logic_vector(125, 8),
41416 => conv_std_logic_vector(125, 8),
41417 => conv_std_logic_vector(126, 8),
41418 => conv_std_logic_vector(127, 8),
41419 => conv_std_logic_vector(127, 8),
41420 => conv_std_logic_vector(128, 8),
41421 => conv_std_logic_vector(128, 8),
41422 => conv_std_logic_vector(129, 8),
41423 => conv_std_logic_vector(130, 8),
41424 => conv_std_logic_vector(130, 8),
41425 => conv_std_logic_vector(131, 8),
41426 => conv_std_logic_vector(132, 8),
41427 => conv_std_logic_vector(132, 8),
41428 => conv_std_logic_vector(133, 8),
41429 => conv_std_logic_vector(133, 8),
41430 => conv_std_logic_vector(134, 8),
41431 => conv_std_logic_vector(135, 8),
41432 => conv_std_logic_vector(135, 8),
41433 => conv_std_logic_vector(136, 8),
41434 => conv_std_logic_vector(137, 8),
41435 => conv_std_logic_vector(137, 8),
41436 => conv_std_logic_vector(138, 8),
41437 => conv_std_logic_vector(138, 8),
41438 => conv_std_logic_vector(139, 8),
41439 => conv_std_logic_vector(140, 8),
41440 => conv_std_logic_vector(140, 8),
41441 => conv_std_logic_vector(141, 8),
41442 => conv_std_logic_vector(142, 8),
41443 => conv_std_logic_vector(142, 8),
41444 => conv_std_logic_vector(143, 8),
41445 => conv_std_logic_vector(144, 8),
41446 => conv_std_logic_vector(144, 8),
41447 => conv_std_logic_vector(145, 8),
41448 => conv_std_logic_vector(145, 8),
41449 => conv_std_logic_vector(146, 8),
41450 => conv_std_logic_vector(147, 8),
41451 => conv_std_logic_vector(147, 8),
41452 => conv_std_logic_vector(148, 8),
41453 => conv_std_logic_vector(149, 8),
41454 => conv_std_logic_vector(149, 8),
41455 => conv_std_logic_vector(150, 8),
41456 => conv_std_logic_vector(150, 8),
41457 => conv_std_logic_vector(151, 8),
41458 => conv_std_logic_vector(152, 8),
41459 => conv_std_logic_vector(152, 8),
41460 => conv_std_logic_vector(153, 8),
41461 => conv_std_logic_vector(154, 8),
41462 => conv_std_logic_vector(154, 8),
41463 => conv_std_logic_vector(155, 8),
41464 => conv_std_logic_vector(155, 8),
41465 => conv_std_logic_vector(156, 8),
41466 => conv_std_logic_vector(157, 8),
41467 => conv_std_logic_vector(157, 8),
41468 => conv_std_logic_vector(158, 8),
41469 => conv_std_logic_vector(159, 8),
41470 => conv_std_logic_vector(159, 8),
41471 => conv_std_logic_vector(160, 8),
41472 => conv_std_logic_vector(0, 8),
41473 => conv_std_logic_vector(0, 8),
41474 => conv_std_logic_vector(1, 8),
41475 => conv_std_logic_vector(1, 8),
41476 => conv_std_logic_vector(2, 8),
41477 => conv_std_logic_vector(3, 8),
41478 => conv_std_logic_vector(3, 8),
41479 => conv_std_logic_vector(4, 8),
41480 => conv_std_logic_vector(5, 8),
41481 => conv_std_logic_vector(5, 8),
41482 => conv_std_logic_vector(6, 8),
41483 => conv_std_logic_vector(6, 8),
41484 => conv_std_logic_vector(7, 8),
41485 => conv_std_logic_vector(8, 8),
41486 => conv_std_logic_vector(8, 8),
41487 => conv_std_logic_vector(9, 8),
41488 => conv_std_logic_vector(10, 8),
41489 => conv_std_logic_vector(10, 8),
41490 => conv_std_logic_vector(11, 8),
41491 => conv_std_logic_vector(12, 8),
41492 => conv_std_logic_vector(12, 8),
41493 => conv_std_logic_vector(13, 8),
41494 => conv_std_logic_vector(13, 8),
41495 => conv_std_logic_vector(14, 8),
41496 => conv_std_logic_vector(15, 8),
41497 => conv_std_logic_vector(15, 8),
41498 => conv_std_logic_vector(16, 8),
41499 => conv_std_logic_vector(17, 8),
41500 => conv_std_logic_vector(17, 8),
41501 => conv_std_logic_vector(18, 8),
41502 => conv_std_logic_vector(18, 8),
41503 => conv_std_logic_vector(19, 8),
41504 => conv_std_logic_vector(20, 8),
41505 => conv_std_logic_vector(20, 8),
41506 => conv_std_logic_vector(21, 8),
41507 => conv_std_logic_vector(22, 8),
41508 => conv_std_logic_vector(22, 8),
41509 => conv_std_logic_vector(23, 8),
41510 => conv_std_logic_vector(24, 8),
41511 => conv_std_logic_vector(24, 8),
41512 => conv_std_logic_vector(25, 8),
41513 => conv_std_logic_vector(25, 8),
41514 => conv_std_logic_vector(26, 8),
41515 => conv_std_logic_vector(27, 8),
41516 => conv_std_logic_vector(27, 8),
41517 => conv_std_logic_vector(28, 8),
41518 => conv_std_logic_vector(29, 8),
41519 => conv_std_logic_vector(29, 8),
41520 => conv_std_logic_vector(30, 8),
41521 => conv_std_logic_vector(31, 8),
41522 => conv_std_logic_vector(31, 8),
41523 => conv_std_logic_vector(32, 8),
41524 => conv_std_logic_vector(32, 8),
41525 => conv_std_logic_vector(33, 8),
41526 => conv_std_logic_vector(34, 8),
41527 => conv_std_logic_vector(34, 8),
41528 => conv_std_logic_vector(35, 8),
41529 => conv_std_logic_vector(36, 8),
41530 => conv_std_logic_vector(36, 8),
41531 => conv_std_logic_vector(37, 8),
41532 => conv_std_logic_vector(37, 8),
41533 => conv_std_logic_vector(38, 8),
41534 => conv_std_logic_vector(39, 8),
41535 => conv_std_logic_vector(39, 8),
41536 => conv_std_logic_vector(40, 8),
41537 => conv_std_logic_vector(41, 8),
41538 => conv_std_logic_vector(41, 8),
41539 => conv_std_logic_vector(42, 8),
41540 => conv_std_logic_vector(43, 8),
41541 => conv_std_logic_vector(43, 8),
41542 => conv_std_logic_vector(44, 8),
41543 => conv_std_logic_vector(44, 8),
41544 => conv_std_logic_vector(45, 8),
41545 => conv_std_logic_vector(46, 8),
41546 => conv_std_logic_vector(46, 8),
41547 => conv_std_logic_vector(47, 8),
41548 => conv_std_logic_vector(48, 8),
41549 => conv_std_logic_vector(48, 8),
41550 => conv_std_logic_vector(49, 8),
41551 => conv_std_logic_vector(49, 8),
41552 => conv_std_logic_vector(50, 8),
41553 => conv_std_logic_vector(51, 8),
41554 => conv_std_logic_vector(51, 8),
41555 => conv_std_logic_vector(52, 8),
41556 => conv_std_logic_vector(53, 8),
41557 => conv_std_logic_vector(53, 8),
41558 => conv_std_logic_vector(54, 8),
41559 => conv_std_logic_vector(55, 8),
41560 => conv_std_logic_vector(55, 8),
41561 => conv_std_logic_vector(56, 8),
41562 => conv_std_logic_vector(56, 8),
41563 => conv_std_logic_vector(57, 8),
41564 => conv_std_logic_vector(58, 8),
41565 => conv_std_logic_vector(58, 8),
41566 => conv_std_logic_vector(59, 8),
41567 => conv_std_logic_vector(60, 8),
41568 => conv_std_logic_vector(60, 8),
41569 => conv_std_logic_vector(61, 8),
41570 => conv_std_logic_vector(62, 8),
41571 => conv_std_logic_vector(62, 8),
41572 => conv_std_logic_vector(63, 8),
41573 => conv_std_logic_vector(63, 8),
41574 => conv_std_logic_vector(64, 8),
41575 => conv_std_logic_vector(65, 8),
41576 => conv_std_logic_vector(65, 8),
41577 => conv_std_logic_vector(66, 8),
41578 => conv_std_logic_vector(67, 8),
41579 => conv_std_logic_vector(67, 8),
41580 => conv_std_logic_vector(68, 8),
41581 => conv_std_logic_vector(68, 8),
41582 => conv_std_logic_vector(69, 8),
41583 => conv_std_logic_vector(70, 8),
41584 => conv_std_logic_vector(70, 8),
41585 => conv_std_logic_vector(71, 8),
41586 => conv_std_logic_vector(72, 8),
41587 => conv_std_logic_vector(72, 8),
41588 => conv_std_logic_vector(73, 8),
41589 => conv_std_logic_vector(74, 8),
41590 => conv_std_logic_vector(74, 8),
41591 => conv_std_logic_vector(75, 8),
41592 => conv_std_logic_vector(75, 8),
41593 => conv_std_logic_vector(76, 8),
41594 => conv_std_logic_vector(77, 8),
41595 => conv_std_logic_vector(77, 8),
41596 => conv_std_logic_vector(78, 8),
41597 => conv_std_logic_vector(79, 8),
41598 => conv_std_logic_vector(79, 8),
41599 => conv_std_logic_vector(80, 8),
41600 => conv_std_logic_vector(81, 8),
41601 => conv_std_logic_vector(81, 8),
41602 => conv_std_logic_vector(82, 8),
41603 => conv_std_logic_vector(82, 8),
41604 => conv_std_logic_vector(83, 8),
41605 => conv_std_logic_vector(84, 8),
41606 => conv_std_logic_vector(84, 8),
41607 => conv_std_logic_vector(85, 8),
41608 => conv_std_logic_vector(86, 8),
41609 => conv_std_logic_vector(86, 8),
41610 => conv_std_logic_vector(87, 8),
41611 => conv_std_logic_vector(87, 8),
41612 => conv_std_logic_vector(88, 8),
41613 => conv_std_logic_vector(89, 8),
41614 => conv_std_logic_vector(89, 8),
41615 => conv_std_logic_vector(90, 8),
41616 => conv_std_logic_vector(91, 8),
41617 => conv_std_logic_vector(91, 8),
41618 => conv_std_logic_vector(92, 8),
41619 => conv_std_logic_vector(93, 8),
41620 => conv_std_logic_vector(93, 8),
41621 => conv_std_logic_vector(94, 8),
41622 => conv_std_logic_vector(94, 8),
41623 => conv_std_logic_vector(95, 8),
41624 => conv_std_logic_vector(96, 8),
41625 => conv_std_logic_vector(96, 8),
41626 => conv_std_logic_vector(97, 8),
41627 => conv_std_logic_vector(98, 8),
41628 => conv_std_logic_vector(98, 8),
41629 => conv_std_logic_vector(99, 8),
41630 => conv_std_logic_vector(99, 8),
41631 => conv_std_logic_vector(100, 8),
41632 => conv_std_logic_vector(101, 8),
41633 => conv_std_logic_vector(101, 8),
41634 => conv_std_logic_vector(102, 8),
41635 => conv_std_logic_vector(103, 8),
41636 => conv_std_logic_vector(103, 8),
41637 => conv_std_logic_vector(104, 8),
41638 => conv_std_logic_vector(105, 8),
41639 => conv_std_logic_vector(105, 8),
41640 => conv_std_logic_vector(106, 8),
41641 => conv_std_logic_vector(106, 8),
41642 => conv_std_logic_vector(107, 8),
41643 => conv_std_logic_vector(108, 8),
41644 => conv_std_logic_vector(108, 8),
41645 => conv_std_logic_vector(109, 8),
41646 => conv_std_logic_vector(110, 8),
41647 => conv_std_logic_vector(110, 8),
41648 => conv_std_logic_vector(111, 8),
41649 => conv_std_logic_vector(112, 8),
41650 => conv_std_logic_vector(112, 8),
41651 => conv_std_logic_vector(113, 8),
41652 => conv_std_logic_vector(113, 8),
41653 => conv_std_logic_vector(114, 8),
41654 => conv_std_logic_vector(115, 8),
41655 => conv_std_logic_vector(115, 8),
41656 => conv_std_logic_vector(116, 8),
41657 => conv_std_logic_vector(117, 8),
41658 => conv_std_logic_vector(117, 8),
41659 => conv_std_logic_vector(118, 8),
41660 => conv_std_logic_vector(118, 8),
41661 => conv_std_logic_vector(119, 8),
41662 => conv_std_logic_vector(120, 8),
41663 => conv_std_logic_vector(120, 8),
41664 => conv_std_logic_vector(121, 8),
41665 => conv_std_logic_vector(122, 8),
41666 => conv_std_logic_vector(122, 8),
41667 => conv_std_logic_vector(123, 8),
41668 => conv_std_logic_vector(124, 8),
41669 => conv_std_logic_vector(124, 8),
41670 => conv_std_logic_vector(125, 8),
41671 => conv_std_logic_vector(125, 8),
41672 => conv_std_logic_vector(126, 8),
41673 => conv_std_logic_vector(127, 8),
41674 => conv_std_logic_vector(127, 8),
41675 => conv_std_logic_vector(128, 8),
41676 => conv_std_logic_vector(129, 8),
41677 => conv_std_logic_vector(129, 8),
41678 => conv_std_logic_vector(130, 8),
41679 => conv_std_logic_vector(130, 8),
41680 => conv_std_logic_vector(131, 8),
41681 => conv_std_logic_vector(132, 8),
41682 => conv_std_logic_vector(132, 8),
41683 => conv_std_logic_vector(133, 8),
41684 => conv_std_logic_vector(134, 8),
41685 => conv_std_logic_vector(134, 8),
41686 => conv_std_logic_vector(135, 8),
41687 => conv_std_logic_vector(136, 8),
41688 => conv_std_logic_vector(136, 8),
41689 => conv_std_logic_vector(137, 8),
41690 => conv_std_logic_vector(137, 8),
41691 => conv_std_logic_vector(138, 8),
41692 => conv_std_logic_vector(139, 8),
41693 => conv_std_logic_vector(139, 8),
41694 => conv_std_logic_vector(140, 8),
41695 => conv_std_logic_vector(141, 8),
41696 => conv_std_logic_vector(141, 8),
41697 => conv_std_logic_vector(142, 8),
41698 => conv_std_logic_vector(143, 8),
41699 => conv_std_logic_vector(143, 8),
41700 => conv_std_logic_vector(144, 8),
41701 => conv_std_logic_vector(144, 8),
41702 => conv_std_logic_vector(145, 8),
41703 => conv_std_logic_vector(146, 8),
41704 => conv_std_logic_vector(146, 8),
41705 => conv_std_logic_vector(147, 8),
41706 => conv_std_logic_vector(148, 8),
41707 => conv_std_logic_vector(148, 8),
41708 => conv_std_logic_vector(149, 8),
41709 => conv_std_logic_vector(149, 8),
41710 => conv_std_logic_vector(150, 8),
41711 => conv_std_logic_vector(151, 8),
41712 => conv_std_logic_vector(151, 8),
41713 => conv_std_logic_vector(152, 8),
41714 => conv_std_logic_vector(153, 8),
41715 => conv_std_logic_vector(153, 8),
41716 => conv_std_logic_vector(154, 8),
41717 => conv_std_logic_vector(155, 8),
41718 => conv_std_logic_vector(155, 8),
41719 => conv_std_logic_vector(156, 8),
41720 => conv_std_logic_vector(156, 8),
41721 => conv_std_logic_vector(157, 8),
41722 => conv_std_logic_vector(158, 8),
41723 => conv_std_logic_vector(158, 8),
41724 => conv_std_logic_vector(159, 8),
41725 => conv_std_logic_vector(160, 8),
41726 => conv_std_logic_vector(160, 8),
41727 => conv_std_logic_vector(161, 8),
41728 => conv_std_logic_vector(0, 8),
41729 => conv_std_logic_vector(0, 8),
41730 => conv_std_logic_vector(1, 8),
41731 => conv_std_logic_vector(1, 8),
41732 => conv_std_logic_vector(2, 8),
41733 => conv_std_logic_vector(3, 8),
41734 => conv_std_logic_vector(3, 8),
41735 => conv_std_logic_vector(4, 8),
41736 => conv_std_logic_vector(5, 8),
41737 => conv_std_logic_vector(5, 8),
41738 => conv_std_logic_vector(6, 8),
41739 => conv_std_logic_vector(7, 8),
41740 => conv_std_logic_vector(7, 8),
41741 => conv_std_logic_vector(8, 8),
41742 => conv_std_logic_vector(8, 8),
41743 => conv_std_logic_vector(9, 8),
41744 => conv_std_logic_vector(10, 8),
41745 => conv_std_logic_vector(10, 8),
41746 => conv_std_logic_vector(11, 8),
41747 => conv_std_logic_vector(12, 8),
41748 => conv_std_logic_vector(12, 8),
41749 => conv_std_logic_vector(13, 8),
41750 => conv_std_logic_vector(14, 8),
41751 => conv_std_logic_vector(14, 8),
41752 => conv_std_logic_vector(15, 8),
41753 => conv_std_logic_vector(15, 8),
41754 => conv_std_logic_vector(16, 8),
41755 => conv_std_logic_vector(17, 8),
41756 => conv_std_logic_vector(17, 8),
41757 => conv_std_logic_vector(18, 8),
41758 => conv_std_logic_vector(19, 8),
41759 => conv_std_logic_vector(19, 8),
41760 => conv_std_logic_vector(20, 8),
41761 => conv_std_logic_vector(21, 8),
41762 => conv_std_logic_vector(21, 8),
41763 => conv_std_logic_vector(22, 8),
41764 => conv_std_logic_vector(22, 8),
41765 => conv_std_logic_vector(23, 8),
41766 => conv_std_logic_vector(24, 8),
41767 => conv_std_logic_vector(24, 8),
41768 => conv_std_logic_vector(25, 8),
41769 => conv_std_logic_vector(26, 8),
41770 => conv_std_logic_vector(26, 8),
41771 => conv_std_logic_vector(27, 8),
41772 => conv_std_logic_vector(28, 8),
41773 => conv_std_logic_vector(28, 8),
41774 => conv_std_logic_vector(29, 8),
41775 => conv_std_logic_vector(29, 8),
41776 => conv_std_logic_vector(30, 8),
41777 => conv_std_logic_vector(31, 8),
41778 => conv_std_logic_vector(31, 8),
41779 => conv_std_logic_vector(32, 8),
41780 => conv_std_logic_vector(33, 8),
41781 => conv_std_logic_vector(33, 8),
41782 => conv_std_logic_vector(34, 8),
41783 => conv_std_logic_vector(35, 8),
41784 => conv_std_logic_vector(35, 8),
41785 => conv_std_logic_vector(36, 8),
41786 => conv_std_logic_vector(36, 8),
41787 => conv_std_logic_vector(37, 8),
41788 => conv_std_logic_vector(38, 8),
41789 => conv_std_logic_vector(38, 8),
41790 => conv_std_logic_vector(39, 8),
41791 => conv_std_logic_vector(40, 8),
41792 => conv_std_logic_vector(40, 8),
41793 => conv_std_logic_vector(41, 8),
41794 => conv_std_logic_vector(42, 8),
41795 => conv_std_logic_vector(42, 8),
41796 => conv_std_logic_vector(43, 8),
41797 => conv_std_logic_vector(43, 8),
41798 => conv_std_logic_vector(44, 8),
41799 => conv_std_logic_vector(45, 8),
41800 => conv_std_logic_vector(45, 8),
41801 => conv_std_logic_vector(46, 8),
41802 => conv_std_logic_vector(47, 8),
41803 => conv_std_logic_vector(47, 8),
41804 => conv_std_logic_vector(48, 8),
41805 => conv_std_logic_vector(49, 8),
41806 => conv_std_logic_vector(49, 8),
41807 => conv_std_logic_vector(50, 8),
41808 => conv_std_logic_vector(50, 8),
41809 => conv_std_logic_vector(51, 8),
41810 => conv_std_logic_vector(52, 8),
41811 => conv_std_logic_vector(52, 8),
41812 => conv_std_logic_vector(53, 8),
41813 => conv_std_logic_vector(54, 8),
41814 => conv_std_logic_vector(54, 8),
41815 => conv_std_logic_vector(55, 8),
41816 => conv_std_logic_vector(56, 8),
41817 => conv_std_logic_vector(56, 8),
41818 => conv_std_logic_vector(57, 8),
41819 => conv_std_logic_vector(57, 8),
41820 => conv_std_logic_vector(58, 8),
41821 => conv_std_logic_vector(59, 8),
41822 => conv_std_logic_vector(59, 8),
41823 => conv_std_logic_vector(60, 8),
41824 => conv_std_logic_vector(61, 8),
41825 => conv_std_logic_vector(61, 8),
41826 => conv_std_logic_vector(62, 8),
41827 => conv_std_logic_vector(63, 8),
41828 => conv_std_logic_vector(63, 8),
41829 => conv_std_logic_vector(64, 8),
41830 => conv_std_logic_vector(64, 8),
41831 => conv_std_logic_vector(65, 8),
41832 => conv_std_logic_vector(66, 8),
41833 => conv_std_logic_vector(66, 8),
41834 => conv_std_logic_vector(67, 8),
41835 => conv_std_logic_vector(68, 8),
41836 => conv_std_logic_vector(68, 8),
41837 => conv_std_logic_vector(69, 8),
41838 => conv_std_logic_vector(70, 8),
41839 => conv_std_logic_vector(70, 8),
41840 => conv_std_logic_vector(71, 8),
41841 => conv_std_logic_vector(71, 8),
41842 => conv_std_logic_vector(72, 8),
41843 => conv_std_logic_vector(73, 8),
41844 => conv_std_logic_vector(73, 8),
41845 => conv_std_logic_vector(74, 8),
41846 => conv_std_logic_vector(75, 8),
41847 => conv_std_logic_vector(75, 8),
41848 => conv_std_logic_vector(76, 8),
41849 => conv_std_logic_vector(77, 8),
41850 => conv_std_logic_vector(77, 8),
41851 => conv_std_logic_vector(78, 8),
41852 => conv_std_logic_vector(78, 8),
41853 => conv_std_logic_vector(79, 8),
41854 => conv_std_logic_vector(80, 8),
41855 => conv_std_logic_vector(80, 8),
41856 => conv_std_logic_vector(81, 8),
41857 => conv_std_logic_vector(82, 8),
41858 => conv_std_logic_vector(82, 8),
41859 => conv_std_logic_vector(83, 8),
41860 => conv_std_logic_vector(84, 8),
41861 => conv_std_logic_vector(84, 8),
41862 => conv_std_logic_vector(85, 8),
41863 => conv_std_logic_vector(85, 8),
41864 => conv_std_logic_vector(86, 8),
41865 => conv_std_logic_vector(87, 8),
41866 => conv_std_logic_vector(87, 8),
41867 => conv_std_logic_vector(88, 8),
41868 => conv_std_logic_vector(89, 8),
41869 => conv_std_logic_vector(89, 8),
41870 => conv_std_logic_vector(90, 8),
41871 => conv_std_logic_vector(91, 8),
41872 => conv_std_logic_vector(91, 8),
41873 => conv_std_logic_vector(92, 8),
41874 => conv_std_logic_vector(92, 8),
41875 => conv_std_logic_vector(93, 8),
41876 => conv_std_logic_vector(94, 8),
41877 => conv_std_logic_vector(94, 8),
41878 => conv_std_logic_vector(95, 8),
41879 => conv_std_logic_vector(96, 8),
41880 => conv_std_logic_vector(96, 8),
41881 => conv_std_logic_vector(97, 8),
41882 => conv_std_logic_vector(98, 8),
41883 => conv_std_logic_vector(98, 8),
41884 => conv_std_logic_vector(99, 8),
41885 => conv_std_logic_vector(99, 8),
41886 => conv_std_logic_vector(100, 8),
41887 => conv_std_logic_vector(101, 8),
41888 => conv_std_logic_vector(101, 8),
41889 => conv_std_logic_vector(102, 8),
41890 => conv_std_logic_vector(103, 8),
41891 => conv_std_logic_vector(103, 8),
41892 => conv_std_logic_vector(104, 8),
41893 => conv_std_logic_vector(105, 8),
41894 => conv_std_logic_vector(105, 8),
41895 => conv_std_logic_vector(106, 8),
41896 => conv_std_logic_vector(106, 8),
41897 => conv_std_logic_vector(107, 8),
41898 => conv_std_logic_vector(108, 8),
41899 => conv_std_logic_vector(108, 8),
41900 => conv_std_logic_vector(109, 8),
41901 => conv_std_logic_vector(110, 8),
41902 => conv_std_logic_vector(110, 8),
41903 => conv_std_logic_vector(111, 8),
41904 => conv_std_logic_vector(112, 8),
41905 => conv_std_logic_vector(112, 8),
41906 => conv_std_logic_vector(113, 8),
41907 => conv_std_logic_vector(113, 8),
41908 => conv_std_logic_vector(114, 8),
41909 => conv_std_logic_vector(115, 8),
41910 => conv_std_logic_vector(115, 8),
41911 => conv_std_logic_vector(116, 8),
41912 => conv_std_logic_vector(117, 8),
41913 => conv_std_logic_vector(117, 8),
41914 => conv_std_logic_vector(118, 8),
41915 => conv_std_logic_vector(119, 8),
41916 => conv_std_logic_vector(119, 8),
41917 => conv_std_logic_vector(120, 8),
41918 => conv_std_logic_vector(120, 8),
41919 => conv_std_logic_vector(121, 8),
41920 => conv_std_logic_vector(122, 8),
41921 => conv_std_logic_vector(122, 8),
41922 => conv_std_logic_vector(123, 8),
41923 => conv_std_logic_vector(124, 8),
41924 => conv_std_logic_vector(124, 8),
41925 => conv_std_logic_vector(125, 8),
41926 => conv_std_logic_vector(126, 8),
41927 => conv_std_logic_vector(126, 8),
41928 => conv_std_logic_vector(127, 8),
41929 => conv_std_logic_vector(127, 8),
41930 => conv_std_logic_vector(128, 8),
41931 => conv_std_logic_vector(129, 8),
41932 => conv_std_logic_vector(129, 8),
41933 => conv_std_logic_vector(130, 8),
41934 => conv_std_logic_vector(131, 8),
41935 => conv_std_logic_vector(131, 8),
41936 => conv_std_logic_vector(132, 8),
41937 => conv_std_logic_vector(133, 8),
41938 => conv_std_logic_vector(133, 8),
41939 => conv_std_logic_vector(134, 8),
41940 => conv_std_logic_vector(134, 8),
41941 => conv_std_logic_vector(135, 8),
41942 => conv_std_logic_vector(136, 8),
41943 => conv_std_logic_vector(136, 8),
41944 => conv_std_logic_vector(137, 8),
41945 => conv_std_logic_vector(138, 8),
41946 => conv_std_logic_vector(138, 8),
41947 => conv_std_logic_vector(139, 8),
41948 => conv_std_logic_vector(140, 8),
41949 => conv_std_logic_vector(140, 8),
41950 => conv_std_logic_vector(141, 8),
41951 => conv_std_logic_vector(141, 8),
41952 => conv_std_logic_vector(142, 8),
41953 => conv_std_logic_vector(143, 8),
41954 => conv_std_logic_vector(143, 8),
41955 => conv_std_logic_vector(144, 8),
41956 => conv_std_logic_vector(145, 8),
41957 => conv_std_logic_vector(145, 8),
41958 => conv_std_logic_vector(146, 8),
41959 => conv_std_logic_vector(147, 8),
41960 => conv_std_logic_vector(147, 8),
41961 => conv_std_logic_vector(148, 8),
41962 => conv_std_logic_vector(148, 8),
41963 => conv_std_logic_vector(149, 8),
41964 => conv_std_logic_vector(150, 8),
41965 => conv_std_logic_vector(150, 8),
41966 => conv_std_logic_vector(151, 8),
41967 => conv_std_logic_vector(152, 8),
41968 => conv_std_logic_vector(152, 8),
41969 => conv_std_logic_vector(153, 8),
41970 => conv_std_logic_vector(154, 8),
41971 => conv_std_logic_vector(154, 8),
41972 => conv_std_logic_vector(155, 8),
41973 => conv_std_logic_vector(155, 8),
41974 => conv_std_logic_vector(156, 8),
41975 => conv_std_logic_vector(157, 8),
41976 => conv_std_logic_vector(157, 8),
41977 => conv_std_logic_vector(158, 8),
41978 => conv_std_logic_vector(159, 8),
41979 => conv_std_logic_vector(159, 8),
41980 => conv_std_logic_vector(160, 8),
41981 => conv_std_logic_vector(161, 8),
41982 => conv_std_logic_vector(161, 8),
41983 => conv_std_logic_vector(162, 8),
41984 => conv_std_logic_vector(0, 8),
41985 => conv_std_logic_vector(0, 8),
41986 => conv_std_logic_vector(1, 8),
41987 => conv_std_logic_vector(1, 8),
41988 => conv_std_logic_vector(2, 8),
41989 => conv_std_logic_vector(3, 8),
41990 => conv_std_logic_vector(3, 8),
41991 => conv_std_logic_vector(4, 8),
41992 => conv_std_logic_vector(5, 8),
41993 => conv_std_logic_vector(5, 8),
41994 => conv_std_logic_vector(6, 8),
41995 => conv_std_logic_vector(7, 8),
41996 => conv_std_logic_vector(7, 8),
41997 => conv_std_logic_vector(8, 8),
41998 => conv_std_logic_vector(8, 8),
41999 => conv_std_logic_vector(9, 8),
42000 => conv_std_logic_vector(10, 8),
42001 => conv_std_logic_vector(10, 8),
42002 => conv_std_logic_vector(11, 8),
42003 => conv_std_logic_vector(12, 8),
42004 => conv_std_logic_vector(12, 8),
42005 => conv_std_logic_vector(13, 8),
42006 => conv_std_logic_vector(14, 8),
42007 => conv_std_logic_vector(14, 8),
42008 => conv_std_logic_vector(15, 8),
42009 => conv_std_logic_vector(16, 8),
42010 => conv_std_logic_vector(16, 8),
42011 => conv_std_logic_vector(17, 8),
42012 => conv_std_logic_vector(17, 8),
42013 => conv_std_logic_vector(18, 8),
42014 => conv_std_logic_vector(19, 8),
42015 => conv_std_logic_vector(19, 8),
42016 => conv_std_logic_vector(20, 8),
42017 => conv_std_logic_vector(21, 8),
42018 => conv_std_logic_vector(21, 8),
42019 => conv_std_logic_vector(22, 8),
42020 => conv_std_logic_vector(23, 8),
42021 => conv_std_logic_vector(23, 8),
42022 => conv_std_logic_vector(24, 8),
42023 => conv_std_logic_vector(24, 8),
42024 => conv_std_logic_vector(25, 8),
42025 => conv_std_logic_vector(26, 8),
42026 => conv_std_logic_vector(26, 8),
42027 => conv_std_logic_vector(27, 8),
42028 => conv_std_logic_vector(28, 8),
42029 => conv_std_logic_vector(28, 8),
42030 => conv_std_logic_vector(29, 8),
42031 => conv_std_logic_vector(30, 8),
42032 => conv_std_logic_vector(30, 8),
42033 => conv_std_logic_vector(31, 8),
42034 => conv_std_logic_vector(32, 8),
42035 => conv_std_logic_vector(32, 8),
42036 => conv_std_logic_vector(33, 8),
42037 => conv_std_logic_vector(33, 8),
42038 => conv_std_logic_vector(34, 8),
42039 => conv_std_logic_vector(35, 8),
42040 => conv_std_logic_vector(35, 8),
42041 => conv_std_logic_vector(36, 8),
42042 => conv_std_logic_vector(37, 8),
42043 => conv_std_logic_vector(37, 8),
42044 => conv_std_logic_vector(38, 8),
42045 => conv_std_logic_vector(39, 8),
42046 => conv_std_logic_vector(39, 8),
42047 => conv_std_logic_vector(40, 8),
42048 => conv_std_logic_vector(41, 8),
42049 => conv_std_logic_vector(41, 8),
42050 => conv_std_logic_vector(42, 8),
42051 => conv_std_logic_vector(42, 8),
42052 => conv_std_logic_vector(43, 8),
42053 => conv_std_logic_vector(44, 8),
42054 => conv_std_logic_vector(44, 8),
42055 => conv_std_logic_vector(45, 8),
42056 => conv_std_logic_vector(46, 8),
42057 => conv_std_logic_vector(46, 8),
42058 => conv_std_logic_vector(47, 8),
42059 => conv_std_logic_vector(48, 8),
42060 => conv_std_logic_vector(48, 8),
42061 => conv_std_logic_vector(49, 8),
42062 => conv_std_logic_vector(49, 8),
42063 => conv_std_logic_vector(50, 8),
42064 => conv_std_logic_vector(51, 8),
42065 => conv_std_logic_vector(51, 8),
42066 => conv_std_logic_vector(52, 8),
42067 => conv_std_logic_vector(53, 8),
42068 => conv_std_logic_vector(53, 8),
42069 => conv_std_logic_vector(54, 8),
42070 => conv_std_logic_vector(55, 8),
42071 => conv_std_logic_vector(55, 8),
42072 => conv_std_logic_vector(56, 8),
42073 => conv_std_logic_vector(57, 8),
42074 => conv_std_logic_vector(57, 8),
42075 => conv_std_logic_vector(58, 8),
42076 => conv_std_logic_vector(58, 8),
42077 => conv_std_logic_vector(59, 8),
42078 => conv_std_logic_vector(60, 8),
42079 => conv_std_logic_vector(60, 8),
42080 => conv_std_logic_vector(61, 8),
42081 => conv_std_logic_vector(62, 8),
42082 => conv_std_logic_vector(62, 8),
42083 => conv_std_logic_vector(63, 8),
42084 => conv_std_logic_vector(64, 8),
42085 => conv_std_logic_vector(64, 8),
42086 => conv_std_logic_vector(65, 8),
42087 => conv_std_logic_vector(65, 8),
42088 => conv_std_logic_vector(66, 8),
42089 => conv_std_logic_vector(67, 8),
42090 => conv_std_logic_vector(67, 8),
42091 => conv_std_logic_vector(68, 8),
42092 => conv_std_logic_vector(69, 8),
42093 => conv_std_logic_vector(69, 8),
42094 => conv_std_logic_vector(70, 8),
42095 => conv_std_logic_vector(71, 8),
42096 => conv_std_logic_vector(71, 8),
42097 => conv_std_logic_vector(72, 8),
42098 => conv_std_logic_vector(73, 8),
42099 => conv_std_logic_vector(73, 8),
42100 => conv_std_logic_vector(74, 8),
42101 => conv_std_logic_vector(74, 8),
42102 => conv_std_logic_vector(75, 8),
42103 => conv_std_logic_vector(76, 8),
42104 => conv_std_logic_vector(76, 8),
42105 => conv_std_logic_vector(77, 8),
42106 => conv_std_logic_vector(78, 8),
42107 => conv_std_logic_vector(78, 8),
42108 => conv_std_logic_vector(79, 8),
42109 => conv_std_logic_vector(80, 8),
42110 => conv_std_logic_vector(80, 8),
42111 => conv_std_logic_vector(81, 8),
42112 => conv_std_logic_vector(82, 8),
42113 => conv_std_logic_vector(82, 8),
42114 => conv_std_logic_vector(83, 8),
42115 => conv_std_logic_vector(83, 8),
42116 => conv_std_logic_vector(84, 8),
42117 => conv_std_logic_vector(85, 8),
42118 => conv_std_logic_vector(85, 8),
42119 => conv_std_logic_vector(86, 8),
42120 => conv_std_logic_vector(87, 8),
42121 => conv_std_logic_vector(87, 8),
42122 => conv_std_logic_vector(88, 8),
42123 => conv_std_logic_vector(89, 8),
42124 => conv_std_logic_vector(89, 8),
42125 => conv_std_logic_vector(90, 8),
42126 => conv_std_logic_vector(90, 8),
42127 => conv_std_logic_vector(91, 8),
42128 => conv_std_logic_vector(92, 8),
42129 => conv_std_logic_vector(92, 8),
42130 => conv_std_logic_vector(93, 8),
42131 => conv_std_logic_vector(94, 8),
42132 => conv_std_logic_vector(94, 8),
42133 => conv_std_logic_vector(95, 8),
42134 => conv_std_logic_vector(96, 8),
42135 => conv_std_logic_vector(96, 8),
42136 => conv_std_logic_vector(97, 8),
42137 => conv_std_logic_vector(98, 8),
42138 => conv_std_logic_vector(98, 8),
42139 => conv_std_logic_vector(99, 8),
42140 => conv_std_logic_vector(99, 8),
42141 => conv_std_logic_vector(100, 8),
42142 => conv_std_logic_vector(101, 8),
42143 => conv_std_logic_vector(101, 8),
42144 => conv_std_logic_vector(102, 8),
42145 => conv_std_logic_vector(103, 8),
42146 => conv_std_logic_vector(103, 8),
42147 => conv_std_logic_vector(104, 8),
42148 => conv_std_logic_vector(105, 8),
42149 => conv_std_logic_vector(105, 8),
42150 => conv_std_logic_vector(106, 8),
42151 => conv_std_logic_vector(106, 8),
42152 => conv_std_logic_vector(107, 8),
42153 => conv_std_logic_vector(108, 8),
42154 => conv_std_logic_vector(108, 8),
42155 => conv_std_logic_vector(109, 8),
42156 => conv_std_logic_vector(110, 8),
42157 => conv_std_logic_vector(110, 8),
42158 => conv_std_logic_vector(111, 8),
42159 => conv_std_logic_vector(112, 8),
42160 => conv_std_logic_vector(112, 8),
42161 => conv_std_logic_vector(113, 8),
42162 => conv_std_logic_vector(114, 8),
42163 => conv_std_logic_vector(114, 8),
42164 => conv_std_logic_vector(115, 8),
42165 => conv_std_logic_vector(115, 8),
42166 => conv_std_logic_vector(116, 8),
42167 => conv_std_logic_vector(117, 8),
42168 => conv_std_logic_vector(117, 8),
42169 => conv_std_logic_vector(118, 8),
42170 => conv_std_logic_vector(119, 8),
42171 => conv_std_logic_vector(119, 8),
42172 => conv_std_logic_vector(120, 8),
42173 => conv_std_logic_vector(121, 8),
42174 => conv_std_logic_vector(121, 8),
42175 => conv_std_logic_vector(122, 8),
42176 => conv_std_logic_vector(123, 8),
42177 => conv_std_logic_vector(123, 8),
42178 => conv_std_logic_vector(124, 8),
42179 => conv_std_logic_vector(124, 8),
42180 => conv_std_logic_vector(125, 8),
42181 => conv_std_logic_vector(126, 8),
42182 => conv_std_logic_vector(126, 8),
42183 => conv_std_logic_vector(127, 8),
42184 => conv_std_logic_vector(128, 8),
42185 => conv_std_logic_vector(128, 8),
42186 => conv_std_logic_vector(129, 8),
42187 => conv_std_logic_vector(130, 8),
42188 => conv_std_logic_vector(130, 8),
42189 => conv_std_logic_vector(131, 8),
42190 => conv_std_logic_vector(131, 8),
42191 => conv_std_logic_vector(132, 8),
42192 => conv_std_logic_vector(133, 8),
42193 => conv_std_logic_vector(133, 8),
42194 => conv_std_logic_vector(134, 8),
42195 => conv_std_logic_vector(135, 8),
42196 => conv_std_logic_vector(135, 8),
42197 => conv_std_logic_vector(136, 8),
42198 => conv_std_logic_vector(137, 8),
42199 => conv_std_logic_vector(137, 8),
42200 => conv_std_logic_vector(138, 8),
42201 => conv_std_logic_vector(139, 8),
42202 => conv_std_logic_vector(139, 8),
42203 => conv_std_logic_vector(140, 8),
42204 => conv_std_logic_vector(140, 8),
42205 => conv_std_logic_vector(141, 8),
42206 => conv_std_logic_vector(142, 8),
42207 => conv_std_logic_vector(142, 8),
42208 => conv_std_logic_vector(143, 8),
42209 => conv_std_logic_vector(144, 8),
42210 => conv_std_logic_vector(144, 8),
42211 => conv_std_logic_vector(145, 8),
42212 => conv_std_logic_vector(146, 8),
42213 => conv_std_logic_vector(146, 8),
42214 => conv_std_logic_vector(147, 8),
42215 => conv_std_logic_vector(147, 8),
42216 => conv_std_logic_vector(148, 8),
42217 => conv_std_logic_vector(149, 8),
42218 => conv_std_logic_vector(149, 8),
42219 => conv_std_logic_vector(150, 8),
42220 => conv_std_logic_vector(151, 8),
42221 => conv_std_logic_vector(151, 8),
42222 => conv_std_logic_vector(152, 8),
42223 => conv_std_logic_vector(153, 8),
42224 => conv_std_logic_vector(153, 8),
42225 => conv_std_logic_vector(154, 8),
42226 => conv_std_logic_vector(155, 8),
42227 => conv_std_logic_vector(155, 8),
42228 => conv_std_logic_vector(156, 8),
42229 => conv_std_logic_vector(156, 8),
42230 => conv_std_logic_vector(157, 8),
42231 => conv_std_logic_vector(158, 8),
42232 => conv_std_logic_vector(158, 8),
42233 => conv_std_logic_vector(159, 8),
42234 => conv_std_logic_vector(160, 8),
42235 => conv_std_logic_vector(160, 8),
42236 => conv_std_logic_vector(161, 8),
42237 => conv_std_logic_vector(162, 8),
42238 => conv_std_logic_vector(162, 8),
42239 => conv_std_logic_vector(163, 8),
42240 => conv_std_logic_vector(0, 8),
42241 => conv_std_logic_vector(0, 8),
42242 => conv_std_logic_vector(1, 8),
42243 => conv_std_logic_vector(1, 8),
42244 => conv_std_logic_vector(2, 8),
42245 => conv_std_logic_vector(3, 8),
42246 => conv_std_logic_vector(3, 8),
42247 => conv_std_logic_vector(4, 8),
42248 => conv_std_logic_vector(5, 8),
42249 => conv_std_logic_vector(5, 8),
42250 => conv_std_logic_vector(6, 8),
42251 => conv_std_logic_vector(7, 8),
42252 => conv_std_logic_vector(7, 8),
42253 => conv_std_logic_vector(8, 8),
42254 => conv_std_logic_vector(9, 8),
42255 => conv_std_logic_vector(9, 8),
42256 => conv_std_logic_vector(10, 8),
42257 => conv_std_logic_vector(10, 8),
42258 => conv_std_logic_vector(11, 8),
42259 => conv_std_logic_vector(12, 8),
42260 => conv_std_logic_vector(12, 8),
42261 => conv_std_logic_vector(13, 8),
42262 => conv_std_logic_vector(14, 8),
42263 => conv_std_logic_vector(14, 8),
42264 => conv_std_logic_vector(15, 8),
42265 => conv_std_logic_vector(16, 8),
42266 => conv_std_logic_vector(16, 8),
42267 => conv_std_logic_vector(17, 8),
42268 => conv_std_logic_vector(18, 8),
42269 => conv_std_logic_vector(18, 8),
42270 => conv_std_logic_vector(19, 8),
42271 => conv_std_logic_vector(19, 8),
42272 => conv_std_logic_vector(20, 8),
42273 => conv_std_logic_vector(21, 8),
42274 => conv_std_logic_vector(21, 8),
42275 => conv_std_logic_vector(22, 8),
42276 => conv_std_logic_vector(23, 8),
42277 => conv_std_logic_vector(23, 8),
42278 => conv_std_logic_vector(24, 8),
42279 => conv_std_logic_vector(25, 8),
42280 => conv_std_logic_vector(25, 8),
42281 => conv_std_logic_vector(26, 8),
42282 => conv_std_logic_vector(27, 8),
42283 => conv_std_logic_vector(27, 8),
42284 => conv_std_logic_vector(28, 8),
42285 => conv_std_logic_vector(29, 8),
42286 => conv_std_logic_vector(29, 8),
42287 => conv_std_logic_vector(30, 8),
42288 => conv_std_logic_vector(30, 8),
42289 => conv_std_logic_vector(31, 8),
42290 => conv_std_logic_vector(32, 8),
42291 => conv_std_logic_vector(32, 8),
42292 => conv_std_logic_vector(33, 8),
42293 => conv_std_logic_vector(34, 8),
42294 => conv_std_logic_vector(34, 8),
42295 => conv_std_logic_vector(35, 8),
42296 => conv_std_logic_vector(36, 8),
42297 => conv_std_logic_vector(36, 8),
42298 => conv_std_logic_vector(37, 8),
42299 => conv_std_logic_vector(38, 8),
42300 => conv_std_logic_vector(38, 8),
42301 => conv_std_logic_vector(39, 8),
42302 => conv_std_logic_vector(39, 8),
42303 => conv_std_logic_vector(40, 8),
42304 => conv_std_logic_vector(41, 8),
42305 => conv_std_logic_vector(41, 8),
42306 => conv_std_logic_vector(42, 8),
42307 => conv_std_logic_vector(43, 8),
42308 => conv_std_logic_vector(43, 8),
42309 => conv_std_logic_vector(44, 8),
42310 => conv_std_logic_vector(45, 8),
42311 => conv_std_logic_vector(45, 8),
42312 => conv_std_logic_vector(46, 8),
42313 => conv_std_logic_vector(47, 8),
42314 => conv_std_logic_vector(47, 8),
42315 => conv_std_logic_vector(48, 8),
42316 => conv_std_logic_vector(48, 8),
42317 => conv_std_logic_vector(49, 8),
42318 => conv_std_logic_vector(50, 8),
42319 => conv_std_logic_vector(50, 8),
42320 => conv_std_logic_vector(51, 8),
42321 => conv_std_logic_vector(52, 8),
42322 => conv_std_logic_vector(52, 8),
42323 => conv_std_logic_vector(53, 8),
42324 => conv_std_logic_vector(54, 8),
42325 => conv_std_logic_vector(54, 8),
42326 => conv_std_logic_vector(55, 8),
42327 => conv_std_logic_vector(56, 8),
42328 => conv_std_logic_vector(56, 8),
42329 => conv_std_logic_vector(57, 8),
42330 => conv_std_logic_vector(58, 8),
42331 => conv_std_logic_vector(58, 8),
42332 => conv_std_logic_vector(59, 8),
42333 => conv_std_logic_vector(59, 8),
42334 => conv_std_logic_vector(60, 8),
42335 => conv_std_logic_vector(61, 8),
42336 => conv_std_logic_vector(61, 8),
42337 => conv_std_logic_vector(62, 8),
42338 => conv_std_logic_vector(63, 8),
42339 => conv_std_logic_vector(63, 8),
42340 => conv_std_logic_vector(64, 8),
42341 => conv_std_logic_vector(65, 8),
42342 => conv_std_logic_vector(65, 8),
42343 => conv_std_logic_vector(66, 8),
42344 => conv_std_logic_vector(67, 8),
42345 => conv_std_logic_vector(67, 8),
42346 => conv_std_logic_vector(68, 8),
42347 => conv_std_logic_vector(68, 8),
42348 => conv_std_logic_vector(69, 8),
42349 => conv_std_logic_vector(70, 8),
42350 => conv_std_logic_vector(70, 8),
42351 => conv_std_logic_vector(71, 8),
42352 => conv_std_logic_vector(72, 8),
42353 => conv_std_logic_vector(72, 8),
42354 => conv_std_logic_vector(73, 8),
42355 => conv_std_logic_vector(74, 8),
42356 => conv_std_logic_vector(74, 8),
42357 => conv_std_logic_vector(75, 8),
42358 => conv_std_logic_vector(76, 8),
42359 => conv_std_logic_vector(76, 8),
42360 => conv_std_logic_vector(77, 8),
42361 => conv_std_logic_vector(77, 8),
42362 => conv_std_logic_vector(78, 8),
42363 => conv_std_logic_vector(79, 8),
42364 => conv_std_logic_vector(79, 8),
42365 => conv_std_logic_vector(80, 8),
42366 => conv_std_logic_vector(81, 8),
42367 => conv_std_logic_vector(81, 8),
42368 => conv_std_logic_vector(82, 8),
42369 => conv_std_logic_vector(83, 8),
42370 => conv_std_logic_vector(83, 8),
42371 => conv_std_logic_vector(84, 8),
42372 => conv_std_logic_vector(85, 8),
42373 => conv_std_logic_vector(85, 8),
42374 => conv_std_logic_vector(86, 8),
42375 => conv_std_logic_vector(87, 8),
42376 => conv_std_logic_vector(87, 8),
42377 => conv_std_logic_vector(88, 8),
42378 => conv_std_logic_vector(88, 8),
42379 => conv_std_logic_vector(89, 8),
42380 => conv_std_logic_vector(90, 8),
42381 => conv_std_logic_vector(90, 8),
42382 => conv_std_logic_vector(91, 8),
42383 => conv_std_logic_vector(92, 8),
42384 => conv_std_logic_vector(92, 8),
42385 => conv_std_logic_vector(93, 8),
42386 => conv_std_logic_vector(94, 8),
42387 => conv_std_logic_vector(94, 8),
42388 => conv_std_logic_vector(95, 8),
42389 => conv_std_logic_vector(96, 8),
42390 => conv_std_logic_vector(96, 8),
42391 => conv_std_logic_vector(97, 8),
42392 => conv_std_logic_vector(97, 8),
42393 => conv_std_logic_vector(98, 8),
42394 => conv_std_logic_vector(99, 8),
42395 => conv_std_logic_vector(99, 8),
42396 => conv_std_logic_vector(100, 8),
42397 => conv_std_logic_vector(101, 8),
42398 => conv_std_logic_vector(101, 8),
42399 => conv_std_logic_vector(102, 8),
42400 => conv_std_logic_vector(103, 8),
42401 => conv_std_logic_vector(103, 8),
42402 => conv_std_logic_vector(104, 8),
42403 => conv_std_logic_vector(105, 8),
42404 => conv_std_logic_vector(105, 8),
42405 => conv_std_logic_vector(106, 8),
42406 => conv_std_logic_vector(106, 8),
42407 => conv_std_logic_vector(107, 8),
42408 => conv_std_logic_vector(108, 8),
42409 => conv_std_logic_vector(108, 8),
42410 => conv_std_logic_vector(109, 8),
42411 => conv_std_logic_vector(110, 8),
42412 => conv_std_logic_vector(110, 8),
42413 => conv_std_logic_vector(111, 8),
42414 => conv_std_logic_vector(112, 8),
42415 => conv_std_logic_vector(112, 8),
42416 => conv_std_logic_vector(113, 8),
42417 => conv_std_logic_vector(114, 8),
42418 => conv_std_logic_vector(114, 8),
42419 => conv_std_logic_vector(115, 8),
42420 => conv_std_logic_vector(116, 8),
42421 => conv_std_logic_vector(116, 8),
42422 => conv_std_logic_vector(117, 8),
42423 => conv_std_logic_vector(117, 8),
42424 => conv_std_logic_vector(118, 8),
42425 => conv_std_logic_vector(119, 8),
42426 => conv_std_logic_vector(119, 8),
42427 => conv_std_logic_vector(120, 8),
42428 => conv_std_logic_vector(121, 8),
42429 => conv_std_logic_vector(121, 8),
42430 => conv_std_logic_vector(122, 8),
42431 => conv_std_logic_vector(123, 8),
42432 => conv_std_logic_vector(123, 8),
42433 => conv_std_logic_vector(124, 8),
42434 => conv_std_logic_vector(125, 8),
42435 => conv_std_logic_vector(125, 8),
42436 => conv_std_logic_vector(126, 8),
42437 => conv_std_logic_vector(126, 8),
42438 => conv_std_logic_vector(127, 8),
42439 => conv_std_logic_vector(128, 8),
42440 => conv_std_logic_vector(128, 8),
42441 => conv_std_logic_vector(129, 8),
42442 => conv_std_logic_vector(130, 8),
42443 => conv_std_logic_vector(130, 8),
42444 => conv_std_logic_vector(131, 8),
42445 => conv_std_logic_vector(132, 8),
42446 => conv_std_logic_vector(132, 8),
42447 => conv_std_logic_vector(133, 8),
42448 => conv_std_logic_vector(134, 8),
42449 => conv_std_logic_vector(134, 8),
42450 => conv_std_logic_vector(135, 8),
42451 => conv_std_logic_vector(135, 8),
42452 => conv_std_logic_vector(136, 8),
42453 => conv_std_logic_vector(137, 8),
42454 => conv_std_logic_vector(137, 8),
42455 => conv_std_logic_vector(138, 8),
42456 => conv_std_logic_vector(139, 8),
42457 => conv_std_logic_vector(139, 8),
42458 => conv_std_logic_vector(140, 8),
42459 => conv_std_logic_vector(141, 8),
42460 => conv_std_logic_vector(141, 8),
42461 => conv_std_logic_vector(142, 8),
42462 => conv_std_logic_vector(143, 8),
42463 => conv_std_logic_vector(143, 8),
42464 => conv_std_logic_vector(144, 8),
42465 => conv_std_logic_vector(145, 8),
42466 => conv_std_logic_vector(145, 8),
42467 => conv_std_logic_vector(146, 8),
42468 => conv_std_logic_vector(146, 8),
42469 => conv_std_logic_vector(147, 8),
42470 => conv_std_logic_vector(148, 8),
42471 => conv_std_logic_vector(148, 8),
42472 => conv_std_logic_vector(149, 8),
42473 => conv_std_logic_vector(150, 8),
42474 => conv_std_logic_vector(150, 8),
42475 => conv_std_logic_vector(151, 8),
42476 => conv_std_logic_vector(152, 8),
42477 => conv_std_logic_vector(152, 8),
42478 => conv_std_logic_vector(153, 8),
42479 => conv_std_logic_vector(154, 8),
42480 => conv_std_logic_vector(154, 8),
42481 => conv_std_logic_vector(155, 8),
42482 => conv_std_logic_vector(155, 8),
42483 => conv_std_logic_vector(156, 8),
42484 => conv_std_logic_vector(157, 8),
42485 => conv_std_logic_vector(157, 8),
42486 => conv_std_logic_vector(158, 8),
42487 => conv_std_logic_vector(159, 8),
42488 => conv_std_logic_vector(159, 8),
42489 => conv_std_logic_vector(160, 8),
42490 => conv_std_logic_vector(161, 8),
42491 => conv_std_logic_vector(161, 8),
42492 => conv_std_logic_vector(162, 8),
42493 => conv_std_logic_vector(163, 8),
42494 => conv_std_logic_vector(163, 8),
42495 => conv_std_logic_vector(164, 8),
42496 => conv_std_logic_vector(0, 8),
42497 => conv_std_logic_vector(0, 8),
42498 => conv_std_logic_vector(1, 8),
42499 => conv_std_logic_vector(1, 8),
42500 => conv_std_logic_vector(2, 8),
42501 => conv_std_logic_vector(3, 8),
42502 => conv_std_logic_vector(3, 8),
42503 => conv_std_logic_vector(4, 8),
42504 => conv_std_logic_vector(5, 8),
42505 => conv_std_logic_vector(5, 8),
42506 => conv_std_logic_vector(6, 8),
42507 => conv_std_logic_vector(7, 8),
42508 => conv_std_logic_vector(7, 8),
42509 => conv_std_logic_vector(8, 8),
42510 => conv_std_logic_vector(9, 8),
42511 => conv_std_logic_vector(9, 8),
42512 => conv_std_logic_vector(10, 8),
42513 => conv_std_logic_vector(11, 8),
42514 => conv_std_logic_vector(11, 8),
42515 => conv_std_logic_vector(12, 8),
42516 => conv_std_logic_vector(12, 8),
42517 => conv_std_logic_vector(13, 8),
42518 => conv_std_logic_vector(14, 8),
42519 => conv_std_logic_vector(14, 8),
42520 => conv_std_logic_vector(15, 8),
42521 => conv_std_logic_vector(16, 8),
42522 => conv_std_logic_vector(16, 8),
42523 => conv_std_logic_vector(17, 8),
42524 => conv_std_logic_vector(18, 8),
42525 => conv_std_logic_vector(18, 8),
42526 => conv_std_logic_vector(19, 8),
42527 => conv_std_logic_vector(20, 8),
42528 => conv_std_logic_vector(20, 8),
42529 => conv_std_logic_vector(21, 8),
42530 => conv_std_logic_vector(22, 8),
42531 => conv_std_logic_vector(22, 8),
42532 => conv_std_logic_vector(23, 8),
42533 => conv_std_logic_vector(23, 8),
42534 => conv_std_logic_vector(24, 8),
42535 => conv_std_logic_vector(25, 8),
42536 => conv_std_logic_vector(25, 8),
42537 => conv_std_logic_vector(26, 8),
42538 => conv_std_logic_vector(27, 8),
42539 => conv_std_logic_vector(27, 8),
42540 => conv_std_logic_vector(28, 8),
42541 => conv_std_logic_vector(29, 8),
42542 => conv_std_logic_vector(29, 8),
42543 => conv_std_logic_vector(30, 8),
42544 => conv_std_logic_vector(31, 8),
42545 => conv_std_logic_vector(31, 8),
42546 => conv_std_logic_vector(32, 8),
42547 => conv_std_logic_vector(33, 8),
42548 => conv_std_logic_vector(33, 8),
42549 => conv_std_logic_vector(34, 8),
42550 => conv_std_logic_vector(35, 8),
42551 => conv_std_logic_vector(35, 8),
42552 => conv_std_logic_vector(36, 8),
42553 => conv_std_logic_vector(36, 8),
42554 => conv_std_logic_vector(37, 8),
42555 => conv_std_logic_vector(38, 8),
42556 => conv_std_logic_vector(38, 8),
42557 => conv_std_logic_vector(39, 8),
42558 => conv_std_logic_vector(40, 8),
42559 => conv_std_logic_vector(40, 8),
42560 => conv_std_logic_vector(41, 8),
42561 => conv_std_logic_vector(42, 8),
42562 => conv_std_logic_vector(42, 8),
42563 => conv_std_logic_vector(43, 8),
42564 => conv_std_logic_vector(44, 8),
42565 => conv_std_logic_vector(44, 8),
42566 => conv_std_logic_vector(45, 8),
42567 => conv_std_logic_vector(46, 8),
42568 => conv_std_logic_vector(46, 8),
42569 => conv_std_logic_vector(47, 8),
42570 => conv_std_logic_vector(47, 8),
42571 => conv_std_logic_vector(48, 8),
42572 => conv_std_logic_vector(49, 8),
42573 => conv_std_logic_vector(49, 8),
42574 => conv_std_logic_vector(50, 8),
42575 => conv_std_logic_vector(51, 8),
42576 => conv_std_logic_vector(51, 8),
42577 => conv_std_logic_vector(52, 8),
42578 => conv_std_logic_vector(53, 8),
42579 => conv_std_logic_vector(53, 8),
42580 => conv_std_logic_vector(54, 8),
42581 => conv_std_logic_vector(55, 8),
42582 => conv_std_logic_vector(55, 8),
42583 => conv_std_logic_vector(56, 8),
42584 => conv_std_logic_vector(57, 8),
42585 => conv_std_logic_vector(57, 8),
42586 => conv_std_logic_vector(58, 8),
42587 => conv_std_logic_vector(59, 8),
42588 => conv_std_logic_vector(59, 8),
42589 => conv_std_logic_vector(60, 8),
42590 => conv_std_logic_vector(60, 8),
42591 => conv_std_logic_vector(61, 8),
42592 => conv_std_logic_vector(62, 8),
42593 => conv_std_logic_vector(62, 8),
42594 => conv_std_logic_vector(63, 8),
42595 => conv_std_logic_vector(64, 8),
42596 => conv_std_logic_vector(64, 8),
42597 => conv_std_logic_vector(65, 8),
42598 => conv_std_logic_vector(66, 8),
42599 => conv_std_logic_vector(66, 8),
42600 => conv_std_logic_vector(67, 8),
42601 => conv_std_logic_vector(68, 8),
42602 => conv_std_logic_vector(68, 8),
42603 => conv_std_logic_vector(69, 8),
42604 => conv_std_logic_vector(70, 8),
42605 => conv_std_logic_vector(70, 8),
42606 => conv_std_logic_vector(71, 8),
42607 => conv_std_logic_vector(71, 8),
42608 => conv_std_logic_vector(72, 8),
42609 => conv_std_logic_vector(73, 8),
42610 => conv_std_logic_vector(73, 8),
42611 => conv_std_logic_vector(74, 8),
42612 => conv_std_logic_vector(75, 8),
42613 => conv_std_logic_vector(75, 8),
42614 => conv_std_logic_vector(76, 8),
42615 => conv_std_logic_vector(77, 8),
42616 => conv_std_logic_vector(77, 8),
42617 => conv_std_logic_vector(78, 8),
42618 => conv_std_logic_vector(79, 8),
42619 => conv_std_logic_vector(79, 8),
42620 => conv_std_logic_vector(80, 8),
42621 => conv_std_logic_vector(81, 8),
42622 => conv_std_logic_vector(81, 8),
42623 => conv_std_logic_vector(82, 8),
42624 => conv_std_logic_vector(83, 8),
42625 => conv_std_logic_vector(83, 8),
42626 => conv_std_logic_vector(84, 8),
42627 => conv_std_logic_vector(84, 8),
42628 => conv_std_logic_vector(85, 8),
42629 => conv_std_logic_vector(86, 8),
42630 => conv_std_logic_vector(86, 8),
42631 => conv_std_logic_vector(87, 8),
42632 => conv_std_logic_vector(88, 8),
42633 => conv_std_logic_vector(88, 8),
42634 => conv_std_logic_vector(89, 8),
42635 => conv_std_logic_vector(90, 8),
42636 => conv_std_logic_vector(90, 8),
42637 => conv_std_logic_vector(91, 8),
42638 => conv_std_logic_vector(92, 8),
42639 => conv_std_logic_vector(92, 8),
42640 => conv_std_logic_vector(93, 8),
42641 => conv_std_logic_vector(94, 8),
42642 => conv_std_logic_vector(94, 8),
42643 => conv_std_logic_vector(95, 8),
42644 => conv_std_logic_vector(95, 8),
42645 => conv_std_logic_vector(96, 8),
42646 => conv_std_logic_vector(97, 8),
42647 => conv_std_logic_vector(97, 8),
42648 => conv_std_logic_vector(98, 8),
42649 => conv_std_logic_vector(99, 8),
42650 => conv_std_logic_vector(99, 8),
42651 => conv_std_logic_vector(100, 8),
42652 => conv_std_logic_vector(101, 8),
42653 => conv_std_logic_vector(101, 8),
42654 => conv_std_logic_vector(102, 8),
42655 => conv_std_logic_vector(103, 8),
42656 => conv_std_logic_vector(103, 8),
42657 => conv_std_logic_vector(104, 8),
42658 => conv_std_logic_vector(105, 8),
42659 => conv_std_logic_vector(105, 8),
42660 => conv_std_logic_vector(106, 8),
42661 => conv_std_logic_vector(106, 8),
42662 => conv_std_logic_vector(107, 8),
42663 => conv_std_logic_vector(108, 8),
42664 => conv_std_logic_vector(108, 8),
42665 => conv_std_logic_vector(109, 8),
42666 => conv_std_logic_vector(110, 8),
42667 => conv_std_logic_vector(110, 8),
42668 => conv_std_logic_vector(111, 8),
42669 => conv_std_logic_vector(112, 8),
42670 => conv_std_logic_vector(112, 8),
42671 => conv_std_logic_vector(113, 8),
42672 => conv_std_logic_vector(114, 8),
42673 => conv_std_logic_vector(114, 8),
42674 => conv_std_logic_vector(115, 8),
42675 => conv_std_logic_vector(116, 8),
42676 => conv_std_logic_vector(116, 8),
42677 => conv_std_logic_vector(117, 8),
42678 => conv_std_logic_vector(118, 8),
42679 => conv_std_logic_vector(118, 8),
42680 => conv_std_logic_vector(119, 8),
42681 => conv_std_logic_vector(119, 8),
42682 => conv_std_logic_vector(120, 8),
42683 => conv_std_logic_vector(121, 8),
42684 => conv_std_logic_vector(121, 8),
42685 => conv_std_logic_vector(122, 8),
42686 => conv_std_logic_vector(123, 8),
42687 => conv_std_logic_vector(123, 8),
42688 => conv_std_logic_vector(124, 8),
42689 => conv_std_logic_vector(125, 8),
42690 => conv_std_logic_vector(125, 8),
42691 => conv_std_logic_vector(126, 8),
42692 => conv_std_logic_vector(127, 8),
42693 => conv_std_logic_vector(127, 8),
42694 => conv_std_logic_vector(128, 8),
42695 => conv_std_logic_vector(129, 8),
42696 => conv_std_logic_vector(129, 8),
42697 => conv_std_logic_vector(130, 8),
42698 => conv_std_logic_vector(130, 8),
42699 => conv_std_logic_vector(131, 8),
42700 => conv_std_logic_vector(132, 8),
42701 => conv_std_logic_vector(132, 8),
42702 => conv_std_logic_vector(133, 8),
42703 => conv_std_logic_vector(134, 8),
42704 => conv_std_logic_vector(134, 8),
42705 => conv_std_logic_vector(135, 8),
42706 => conv_std_logic_vector(136, 8),
42707 => conv_std_logic_vector(136, 8),
42708 => conv_std_logic_vector(137, 8),
42709 => conv_std_logic_vector(138, 8),
42710 => conv_std_logic_vector(138, 8),
42711 => conv_std_logic_vector(139, 8),
42712 => conv_std_logic_vector(140, 8),
42713 => conv_std_logic_vector(140, 8),
42714 => conv_std_logic_vector(141, 8),
42715 => conv_std_logic_vector(142, 8),
42716 => conv_std_logic_vector(142, 8),
42717 => conv_std_logic_vector(143, 8),
42718 => conv_std_logic_vector(143, 8),
42719 => conv_std_logic_vector(144, 8),
42720 => conv_std_logic_vector(145, 8),
42721 => conv_std_logic_vector(145, 8),
42722 => conv_std_logic_vector(146, 8),
42723 => conv_std_logic_vector(147, 8),
42724 => conv_std_logic_vector(147, 8),
42725 => conv_std_logic_vector(148, 8),
42726 => conv_std_logic_vector(149, 8),
42727 => conv_std_logic_vector(149, 8),
42728 => conv_std_logic_vector(150, 8),
42729 => conv_std_logic_vector(151, 8),
42730 => conv_std_logic_vector(151, 8),
42731 => conv_std_logic_vector(152, 8),
42732 => conv_std_logic_vector(153, 8),
42733 => conv_std_logic_vector(153, 8),
42734 => conv_std_logic_vector(154, 8),
42735 => conv_std_logic_vector(154, 8),
42736 => conv_std_logic_vector(155, 8),
42737 => conv_std_logic_vector(156, 8),
42738 => conv_std_logic_vector(156, 8),
42739 => conv_std_logic_vector(157, 8),
42740 => conv_std_logic_vector(158, 8),
42741 => conv_std_logic_vector(158, 8),
42742 => conv_std_logic_vector(159, 8),
42743 => conv_std_logic_vector(160, 8),
42744 => conv_std_logic_vector(160, 8),
42745 => conv_std_logic_vector(161, 8),
42746 => conv_std_logic_vector(162, 8),
42747 => conv_std_logic_vector(162, 8),
42748 => conv_std_logic_vector(163, 8),
42749 => conv_std_logic_vector(164, 8),
42750 => conv_std_logic_vector(164, 8),
42751 => conv_std_logic_vector(165, 8),
42752 => conv_std_logic_vector(0, 8),
42753 => conv_std_logic_vector(0, 8),
42754 => conv_std_logic_vector(1, 8),
42755 => conv_std_logic_vector(1, 8),
42756 => conv_std_logic_vector(2, 8),
42757 => conv_std_logic_vector(3, 8),
42758 => conv_std_logic_vector(3, 8),
42759 => conv_std_logic_vector(4, 8),
42760 => conv_std_logic_vector(5, 8),
42761 => conv_std_logic_vector(5, 8),
42762 => conv_std_logic_vector(6, 8),
42763 => conv_std_logic_vector(7, 8),
42764 => conv_std_logic_vector(7, 8),
42765 => conv_std_logic_vector(8, 8),
42766 => conv_std_logic_vector(9, 8),
42767 => conv_std_logic_vector(9, 8),
42768 => conv_std_logic_vector(10, 8),
42769 => conv_std_logic_vector(11, 8),
42770 => conv_std_logic_vector(11, 8),
42771 => conv_std_logic_vector(12, 8),
42772 => conv_std_logic_vector(13, 8),
42773 => conv_std_logic_vector(13, 8),
42774 => conv_std_logic_vector(14, 8),
42775 => conv_std_logic_vector(15, 8),
42776 => conv_std_logic_vector(15, 8),
42777 => conv_std_logic_vector(16, 8),
42778 => conv_std_logic_vector(16, 8),
42779 => conv_std_logic_vector(17, 8),
42780 => conv_std_logic_vector(18, 8),
42781 => conv_std_logic_vector(18, 8),
42782 => conv_std_logic_vector(19, 8),
42783 => conv_std_logic_vector(20, 8),
42784 => conv_std_logic_vector(20, 8),
42785 => conv_std_logic_vector(21, 8),
42786 => conv_std_logic_vector(22, 8),
42787 => conv_std_logic_vector(22, 8),
42788 => conv_std_logic_vector(23, 8),
42789 => conv_std_logic_vector(24, 8),
42790 => conv_std_logic_vector(24, 8),
42791 => conv_std_logic_vector(25, 8),
42792 => conv_std_logic_vector(26, 8),
42793 => conv_std_logic_vector(26, 8),
42794 => conv_std_logic_vector(27, 8),
42795 => conv_std_logic_vector(28, 8),
42796 => conv_std_logic_vector(28, 8),
42797 => conv_std_logic_vector(29, 8),
42798 => conv_std_logic_vector(30, 8),
42799 => conv_std_logic_vector(30, 8),
42800 => conv_std_logic_vector(31, 8),
42801 => conv_std_logic_vector(31, 8),
42802 => conv_std_logic_vector(32, 8),
42803 => conv_std_logic_vector(33, 8),
42804 => conv_std_logic_vector(33, 8),
42805 => conv_std_logic_vector(34, 8),
42806 => conv_std_logic_vector(35, 8),
42807 => conv_std_logic_vector(35, 8),
42808 => conv_std_logic_vector(36, 8),
42809 => conv_std_logic_vector(37, 8),
42810 => conv_std_logic_vector(37, 8),
42811 => conv_std_logic_vector(38, 8),
42812 => conv_std_logic_vector(39, 8),
42813 => conv_std_logic_vector(39, 8),
42814 => conv_std_logic_vector(40, 8),
42815 => conv_std_logic_vector(41, 8),
42816 => conv_std_logic_vector(41, 8),
42817 => conv_std_logic_vector(42, 8),
42818 => conv_std_logic_vector(43, 8),
42819 => conv_std_logic_vector(43, 8),
42820 => conv_std_logic_vector(44, 8),
42821 => conv_std_logic_vector(45, 8),
42822 => conv_std_logic_vector(45, 8),
42823 => conv_std_logic_vector(46, 8),
42824 => conv_std_logic_vector(46, 8),
42825 => conv_std_logic_vector(47, 8),
42826 => conv_std_logic_vector(48, 8),
42827 => conv_std_logic_vector(48, 8),
42828 => conv_std_logic_vector(49, 8),
42829 => conv_std_logic_vector(50, 8),
42830 => conv_std_logic_vector(50, 8),
42831 => conv_std_logic_vector(51, 8),
42832 => conv_std_logic_vector(52, 8),
42833 => conv_std_logic_vector(52, 8),
42834 => conv_std_logic_vector(53, 8),
42835 => conv_std_logic_vector(54, 8),
42836 => conv_std_logic_vector(54, 8),
42837 => conv_std_logic_vector(55, 8),
42838 => conv_std_logic_vector(56, 8),
42839 => conv_std_logic_vector(56, 8),
42840 => conv_std_logic_vector(57, 8),
42841 => conv_std_logic_vector(58, 8),
42842 => conv_std_logic_vector(58, 8),
42843 => conv_std_logic_vector(59, 8),
42844 => conv_std_logic_vector(60, 8),
42845 => conv_std_logic_vector(60, 8),
42846 => conv_std_logic_vector(61, 8),
42847 => conv_std_logic_vector(61, 8),
42848 => conv_std_logic_vector(62, 8),
42849 => conv_std_logic_vector(63, 8),
42850 => conv_std_logic_vector(63, 8),
42851 => conv_std_logic_vector(64, 8),
42852 => conv_std_logic_vector(65, 8),
42853 => conv_std_logic_vector(65, 8),
42854 => conv_std_logic_vector(66, 8),
42855 => conv_std_logic_vector(67, 8),
42856 => conv_std_logic_vector(67, 8),
42857 => conv_std_logic_vector(68, 8),
42858 => conv_std_logic_vector(69, 8),
42859 => conv_std_logic_vector(69, 8),
42860 => conv_std_logic_vector(70, 8),
42861 => conv_std_logic_vector(71, 8),
42862 => conv_std_logic_vector(71, 8),
42863 => conv_std_logic_vector(72, 8),
42864 => conv_std_logic_vector(73, 8),
42865 => conv_std_logic_vector(73, 8),
42866 => conv_std_logic_vector(74, 8),
42867 => conv_std_logic_vector(75, 8),
42868 => conv_std_logic_vector(75, 8),
42869 => conv_std_logic_vector(76, 8),
42870 => conv_std_logic_vector(76, 8),
42871 => conv_std_logic_vector(77, 8),
42872 => conv_std_logic_vector(78, 8),
42873 => conv_std_logic_vector(78, 8),
42874 => conv_std_logic_vector(79, 8),
42875 => conv_std_logic_vector(80, 8),
42876 => conv_std_logic_vector(80, 8),
42877 => conv_std_logic_vector(81, 8),
42878 => conv_std_logic_vector(82, 8),
42879 => conv_std_logic_vector(82, 8),
42880 => conv_std_logic_vector(83, 8),
42881 => conv_std_logic_vector(84, 8),
42882 => conv_std_logic_vector(84, 8),
42883 => conv_std_logic_vector(85, 8),
42884 => conv_std_logic_vector(86, 8),
42885 => conv_std_logic_vector(86, 8),
42886 => conv_std_logic_vector(87, 8),
42887 => conv_std_logic_vector(88, 8),
42888 => conv_std_logic_vector(88, 8),
42889 => conv_std_logic_vector(89, 8),
42890 => conv_std_logic_vector(90, 8),
42891 => conv_std_logic_vector(90, 8),
42892 => conv_std_logic_vector(91, 8),
42893 => conv_std_logic_vector(91, 8),
42894 => conv_std_logic_vector(92, 8),
42895 => conv_std_logic_vector(93, 8),
42896 => conv_std_logic_vector(93, 8),
42897 => conv_std_logic_vector(94, 8),
42898 => conv_std_logic_vector(95, 8),
42899 => conv_std_logic_vector(95, 8),
42900 => conv_std_logic_vector(96, 8),
42901 => conv_std_logic_vector(97, 8),
42902 => conv_std_logic_vector(97, 8),
42903 => conv_std_logic_vector(98, 8),
42904 => conv_std_logic_vector(99, 8),
42905 => conv_std_logic_vector(99, 8),
42906 => conv_std_logic_vector(100, 8),
42907 => conv_std_logic_vector(101, 8),
42908 => conv_std_logic_vector(101, 8),
42909 => conv_std_logic_vector(102, 8),
42910 => conv_std_logic_vector(103, 8),
42911 => conv_std_logic_vector(103, 8),
42912 => conv_std_logic_vector(104, 8),
42913 => conv_std_logic_vector(105, 8),
42914 => conv_std_logic_vector(105, 8),
42915 => conv_std_logic_vector(106, 8),
42916 => conv_std_logic_vector(106, 8),
42917 => conv_std_logic_vector(107, 8),
42918 => conv_std_logic_vector(108, 8),
42919 => conv_std_logic_vector(108, 8),
42920 => conv_std_logic_vector(109, 8),
42921 => conv_std_logic_vector(110, 8),
42922 => conv_std_logic_vector(110, 8),
42923 => conv_std_logic_vector(111, 8),
42924 => conv_std_logic_vector(112, 8),
42925 => conv_std_logic_vector(112, 8),
42926 => conv_std_logic_vector(113, 8),
42927 => conv_std_logic_vector(114, 8),
42928 => conv_std_logic_vector(114, 8),
42929 => conv_std_logic_vector(115, 8),
42930 => conv_std_logic_vector(116, 8),
42931 => conv_std_logic_vector(116, 8),
42932 => conv_std_logic_vector(117, 8),
42933 => conv_std_logic_vector(118, 8),
42934 => conv_std_logic_vector(118, 8),
42935 => conv_std_logic_vector(119, 8),
42936 => conv_std_logic_vector(120, 8),
42937 => conv_std_logic_vector(120, 8),
42938 => conv_std_logic_vector(121, 8),
42939 => conv_std_logic_vector(121, 8),
42940 => conv_std_logic_vector(122, 8),
42941 => conv_std_logic_vector(123, 8),
42942 => conv_std_logic_vector(123, 8),
42943 => conv_std_logic_vector(124, 8),
42944 => conv_std_logic_vector(125, 8),
42945 => conv_std_logic_vector(125, 8),
42946 => conv_std_logic_vector(126, 8),
42947 => conv_std_logic_vector(127, 8),
42948 => conv_std_logic_vector(127, 8),
42949 => conv_std_logic_vector(128, 8),
42950 => conv_std_logic_vector(129, 8),
42951 => conv_std_logic_vector(129, 8),
42952 => conv_std_logic_vector(130, 8),
42953 => conv_std_logic_vector(131, 8),
42954 => conv_std_logic_vector(131, 8),
42955 => conv_std_logic_vector(132, 8),
42956 => conv_std_logic_vector(133, 8),
42957 => conv_std_logic_vector(133, 8),
42958 => conv_std_logic_vector(134, 8),
42959 => conv_std_logic_vector(135, 8),
42960 => conv_std_logic_vector(135, 8),
42961 => conv_std_logic_vector(136, 8),
42962 => conv_std_logic_vector(136, 8),
42963 => conv_std_logic_vector(137, 8),
42964 => conv_std_logic_vector(138, 8),
42965 => conv_std_logic_vector(138, 8),
42966 => conv_std_logic_vector(139, 8),
42967 => conv_std_logic_vector(140, 8),
42968 => conv_std_logic_vector(140, 8),
42969 => conv_std_logic_vector(141, 8),
42970 => conv_std_logic_vector(142, 8),
42971 => conv_std_logic_vector(142, 8),
42972 => conv_std_logic_vector(143, 8),
42973 => conv_std_logic_vector(144, 8),
42974 => conv_std_logic_vector(144, 8),
42975 => conv_std_logic_vector(145, 8),
42976 => conv_std_logic_vector(146, 8),
42977 => conv_std_logic_vector(146, 8),
42978 => conv_std_logic_vector(147, 8),
42979 => conv_std_logic_vector(148, 8),
42980 => conv_std_logic_vector(148, 8),
42981 => conv_std_logic_vector(149, 8),
42982 => conv_std_logic_vector(150, 8),
42983 => conv_std_logic_vector(150, 8),
42984 => conv_std_logic_vector(151, 8),
42985 => conv_std_logic_vector(151, 8),
42986 => conv_std_logic_vector(152, 8),
42987 => conv_std_logic_vector(153, 8),
42988 => conv_std_logic_vector(153, 8),
42989 => conv_std_logic_vector(154, 8),
42990 => conv_std_logic_vector(155, 8),
42991 => conv_std_logic_vector(155, 8),
42992 => conv_std_logic_vector(156, 8),
42993 => conv_std_logic_vector(157, 8),
42994 => conv_std_logic_vector(157, 8),
42995 => conv_std_logic_vector(158, 8),
42996 => conv_std_logic_vector(159, 8),
42997 => conv_std_logic_vector(159, 8),
42998 => conv_std_logic_vector(160, 8),
42999 => conv_std_logic_vector(161, 8),
43000 => conv_std_logic_vector(161, 8),
43001 => conv_std_logic_vector(162, 8),
43002 => conv_std_logic_vector(163, 8),
43003 => conv_std_logic_vector(163, 8),
43004 => conv_std_logic_vector(164, 8),
43005 => conv_std_logic_vector(165, 8),
43006 => conv_std_logic_vector(165, 8),
43007 => conv_std_logic_vector(166, 8),
43008 => conv_std_logic_vector(0, 8),
43009 => conv_std_logic_vector(0, 8),
43010 => conv_std_logic_vector(1, 8),
43011 => conv_std_logic_vector(1, 8),
43012 => conv_std_logic_vector(2, 8),
43013 => conv_std_logic_vector(3, 8),
43014 => conv_std_logic_vector(3, 8),
43015 => conv_std_logic_vector(4, 8),
43016 => conv_std_logic_vector(5, 8),
43017 => conv_std_logic_vector(5, 8),
43018 => conv_std_logic_vector(6, 8),
43019 => conv_std_logic_vector(7, 8),
43020 => conv_std_logic_vector(7, 8),
43021 => conv_std_logic_vector(8, 8),
43022 => conv_std_logic_vector(9, 8),
43023 => conv_std_logic_vector(9, 8),
43024 => conv_std_logic_vector(10, 8),
43025 => conv_std_logic_vector(11, 8),
43026 => conv_std_logic_vector(11, 8),
43027 => conv_std_logic_vector(12, 8),
43028 => conv_std_logic_vector(13, 8),
43029 => conv_std_logic_vector(13, 8),
43030 => conv_std_logic_vector(14, 8),
43031 => conv_std_logic_vector(15, 8),
43032 => conv_std_logic_vector(15, 8),
43033 => conv_std_logic_vector(16, 8),
43034 => conv_std_logic_vector(17, 8),
43035 => conv_std_logic_vector(17, 8),
43036 => conv_std_logic_vector(18, 8),
43037 => conv_std_logic_vector(19, 8),
43038 => conv_std_logic_vector(19, 8),
43039 => conv_std_logic_vector(20, 8),
43040 => conv_std_logic_vector(21, 8),
43041 => conv_std_logic_vector(21, 8),
43042 => conv_std_logic_vector(22, 8),
43043 => conv_std_logic_vector(22, 8),
43044 => conv_std_logic_vector(23, 8),
43045 => conv_std_logic_vector(24, 8),
43046 => conv_std_logic_vector(24, 8),
43047 => conv_std_logic_vector(25, 8),
43048 => conv_std_logic_vector(26, 8),
43049 => conv_std_logic_vector(26, 8),
43050 => conv_std_logic_vector(27, 8),
43051 => conv_std_logic_vector(28, 8),
43052 => conv_std_logic_vector(28, 8),
43053 => conv_std_logic_vector(29, 8),
43054 => conv_std_logic_vector(30, 8),
43055 => conv_std_logic_vector(30, 8),
43056 => conv_std_logic_vector(31, 8),
43057 => conv_std_logic_vector(32, 8),
43058 => conv_std_logic_vector(32, 8),
43059 => conv_std_logic_vector(33, 8),
43060 => conv_std_logic_vector(34, 8),
43061 => conv_std_logic_vector(34, 8),
43062 => conv_std_logic_vector(35, 8),
43063 => conv_std_logic_vector(36, 8),
43064 => conv_std_logic_vector(36, 8),
43065 => conv_std_logic_vector(37, 8),
43066 => conv_std_logic_vector(38, 8),
43067 => conv_std_logic_vector(38, 8),
43068 => conv_std_logic_vector(39, 8),
43069 => conv_std_logic_vector(40, 8),
43070 => conv_std_logic_vector(40, 8),
43071 => conv_std_logic_vector(41, 8),
43072 => conv_std_logic_vector(42, 8),
43073 => conv_std_logic_vector(42, 8),
43074 => conv_std_logic_vector(43, 8),
43075 => conv_std_logic_vector(43, 8),
43076 => conv_std_logic_vector(44, 8),
43077 => conv_std_logic_vector(45, 8),
43078 => conv_std_logic_vector(45, 8),
43079 => conv_std_logic_vector(46, 8),
43080 => conv_std_logic_vector(47, 8),
43081 => conv_std_logic_vector(47, 8),
43082 => conv_std_logic_vector(48, 8),
43083 => conv_std_logic_vector(49, 8),
43084 => conv_std_logic_vector(49, 8),
43085 => conv_std_logic_vector(50, 8),
43086 => conv_std_logic_vector(51, 8),
43087 => conv_std_logic_vector(51, 8),
43088 => conv_std_logic_vector(52, 8),
43089 => conv_std_logic_vector(53, 8),
43090 => conv_std_logic_vector(53, 8),
43091 => conv_std_logic_vector(54, 8),
43092 => conv_std_logic_vector(55, 8),
43093 => conv_std_logic_vector(55, 8),
43094 => conv_std_logic_vector(56, 8),
43095 => conv_std_logic_vector(57, 8),
43096 => conv_std_logic_vector(57, 8),
43097 => conv_std_logic_vector(58, 8),
43098 => conv_std_logic_vector(59, 8),
43099 => conv_std_logic_vector(59, 8),
43100 => conv_std_logic_vector(60, 8),
43101 => conv_std_logic_vector(61, 8),
43102 => conv_std_logic_vector(61, 8),
43103 => conv_std_logic_vector(62, 8),
43104 => conv_std_logic_vector(63, 8),
43105 => conv_std_logic_vector(63, 8),
43106 => conv_std_logic_vector(64, 8),
43107 => conv_std_logic_vector(64, 8),
43108 => conv_std_logic_vector(65, 8),
43109 => conv_std_logic_vector(66, 8),
43110 => conv_std_logic_vector(66, 8),
43111 => conv_std_logic_vector(67, 8),
43112 => conv_std_logic_vector(68, 8),
43113 => conv_std_logic_vector(68, 8),
43114 => conv_std_logic_vector(69, 8),
43115 => conv_std_logic_vector(70, 8),
43116 => conv_std_logic_vector(70, 8),
43117 => conv_std_logic_vector(71, 8),
43118 => conv_std_logic_vector(72, 8),
43119 => conv_std_logic_vector(72, 8),
43120 => conv_std_logic_vector(73, 8),
43121 => conv_std_logic_vector(74, 8),
43122 => conv_std_logic_vector(74, 8),
43123 => conv_std_logic_vector(75, 8),
43124 => conv_std_logic_vector(76, 8),
43125 => conv_std_logic_vector(76, 8),
43126 => conv_std_logic_vector(77, 8),
43127 => conv_std_logic_vector(78, 8),
43128 => conv_std_logic_vector(78, 8),
43129 => conv_std_logic_vector(79, 8),
43130 => conv_std_logic_vector(80, 8),
43131 => conv_std_logic_vector(80, 8),
43132 => conv_std_logic_vector(81, 8),
43133 => conv_std_logic_vector(82, 8),
43134 => conv_std_logic_vector(82, 8),
43135 => conv_std_logic_vector(83, 8),
43136 => conv_std_logic_vector(84, 8),
43137 => conv_std_logic_vector(84, 8),
43138 => conv_std_logic_vector(85, 8),
43139 => conv_std_logic_vector(85, 8),
43140 => conv_std_logic_vector(86, 8),
43141 => conv_std_logic_vector(87, 8),
43142 => conv_std_logic_vector(87, 8),
43143 => conv_std_logic_vector(88, 8),
43144 => conv_std_logic_vector(89, 8),
43145 => conv_std_logic_vector(89, 8),
43146 => conv_std_logic_vector(90, 8),
43147 => conv_std_logic_vector(91, 8),
43148 => conv_std_logic_vector(91, 8),
43149 => conv_std_logic_vector(92, 8),
43150 => conv_std_logic_vector(93, 8),
43151 => conv_std_logic_vector(93, 8),
43152 => conv_std_logic_vector(94, 8),
43153 => conv_std_logic_vector(95, 8),
43154 => conv_std_logic_vector(95, 8),
43155 => conv_std_logic_vector(96, 8),
43156 => conv_std_logic_vector(97, 8),
43157 => conv_std_logic_vector(97, 8),
43158 => conv_std_logic_vector(98, 8),
43159 => conv_std_logic_vector(99, 8),
43160 => conv_std_logic_vector(99, 8),
43161 => conv_std_logic_vector(100, 8),
43162 => conv_std_logic_vector(101, 8),
43163 => conv_std_logic_vector(101, 8),
43164 => conv_std_logic_vector(102, 8),
43165 => conv_std_logic_vector(103, 8),
43166 => conv_std_logic_vector(103, 8),
43167 => conv_std_logic_vector(104, 8),
43168 => conv_std_logic_vector(105, 8),
43169 => conv_std_logic_vector(105, 8),
43170 => conv_std_logic_vector(106, 8),
43171 => conv_std_logic_vector(106, 8),
43172 => conv_std_logic_vector(107, 8),
43173 => conv_std_logic_vector(108, 8),
43174 => conv_std_logic_vector(108, 8),
43175 => conv_std_logic_vector(109, 8),
43176 => conv_std_logic_vector(110, 8),
43177 => conv_std_logic_vector(110, 8),
43178 => conv_std_logic_vector(111, 8),
43179 => conv_std_logic_vector(112, 8),
43180 => conv_std_logic_vector(112, 8),
43181 => conv_std_logic_vector(113, 8),
43182 => conv_std_logic_vector(114, 8),
43183 => conv_std_logic_vector(114, 8),
43184 => conv_std_logic_vector(115, 8),
43185 => conv_std_logic_vector(116, 8),
43186 => conv_std_logic_vector(116, 8),
43187 => conv_std_logic_vector(117, 8),
43188 => conv_std_logic_vector(118, 8),
43189 => conv_std_logic_vector(118, 8),
43190 => conv_std_logic_vector(119, 8),
43191 => conv_std_logic_vector(120, 8),
43192 => conv_std_logic_vector(120, 8),
43193 => conv_std_logic_vector(121, 8),
43194 => conv_std_logic_vector(122, 8),
43195 => conv_std_logic_vector(122, 8),
43196 => conv_std_logic_vector(123, 8),
43197 => conv_std_logic_vector(124, 8),
43198 => conv_std_logic_vector(124, 8),
43199 => conv_std_logic_vector(125, 8),
43200 => conv_std_logic_vector(126, 8),
43201 => conv_std_logic_vector(126, 8),
43202 => conv_std_logic_vector(127, 8),
43203 => conv_std_logic_vector(127, 8),
43204 => conv_std_logic_vector(128, 8),
43205 => conv_std_logic_vector(129, 8),
43206 => conv_std_logic_vector(129, 8),
43207 => conv_std_logic_vector(130, 8),
43208 => conv_std_logic_vector(131, 8),
43209 => conv_std_logic_vector(131, 8),
43210 => conv_std_logic_vector(132, 8),
43211 => conv_std_logic_vector(133, 8),
43212 => conv_std_logic_vector(133, 8),
43213 => conv_std_logic_vector(134, 8),
43214 => conv_std_logic_vector(135, 8),
43215 => conv_std_logic_vector(135, 8),
43216 => conv_std_logic_vector(136, 8),
43217 => conv_std_logic_vector(137, 8),
43218 => conv_std_logic_vector(137, 8),
43219 => conv_std_logic_vector(138, 8),
43220 => conv_std_logic_vector(139, 8),
43221 => conv_std_logic_vector(139, 8),
43222 => conv_std_logic_vector(140, 8),
43223 => conv_std_logic_vector(141, 8),
43224 => conv_std_logic_vector(141, 8),
43225 => conv_std_logic_vector(142, 8),
43226 => conv_std_logic_vector(143, 8),
43227 => conv_std_logic_vector(143, 8),
43228 => conv_std_logic_vector(144, 8),
43229 => conv_std_logic_vector(145, 8),
43230 => conv_std_logic_vector(145, 8),
43231 => conv_std_logic_vector(146, 8),
43232 => conv_std_logic_vector(147, 8),
43233 => conv_std_logic_vector(147, 8),
43234 => conv_std_logic_vector(148, 8),
43235 => conv_std_logic_vector(148, 8),
43236 => conv_std_logic_vector(149, 8),
43237 => conv_std_logic_vector(150, 8),
43238 => conv_std_logic_vector(150, 8),
43239 => conv_std_logic_vector(151, 8),
43240 => conv_std_logic_vector(152, 8),
43241 => conv_std_logic_vector(152, 8),
43242 => conv_std_logic_vector(153, 8),
43243 => conv_std_logic_vector(154, 8),
43244 => conv_std_logic_vector(154, 8),
43245 => conv_std_logic_vector(155, 8),
43246 => conv_std_logic_vector(156, 8),
43247 => conv_std_logic_vector(156, 8),
43248 => conv_std_logic_vector(157, 8),
43249 => conv_std_logic_vector(158, 8),
43250 => conv_std_logic_vector(158, 8),
43251 => conv_std_logic_vector(159, 8),
43252 => conv_std_logic_vector(160, 8),
43253 => conv_std_logic_vector(160, 8),
43254 => conv_std_logic_vector(161, 8),
43255 => conv_std_logic_vector(162, 8),
43256 => conv_std_logic_vector(162, 8),
43257 => conv_std_logic_vector(163, 8),
43258 => conv_std_logic_vector(164, 8),
43259 => conv_std_logic_vector(164, 8),
43260 => conv_std_logic_vector(165, 8),
43261 => conv_std_logic_vector(166, 8),
43262 => conv_std_logic_vector(166, 8),
43263 => conv_std_logic_vector(167, 8),
43264 => conv_std_logic_vector(0, 8),
43265 => conv_std_logic_vector(0, 8),
43266 => conv_std_logic_vector(1, 8),
43267 => conv_std_logic_vector(1, 8),
43268 => conv_std_logic_vector(2, 8),
43269 => conv_std_logic_vector(3, 8),
43270 => conv_std_logic_vector(3, 8),
43271 => conv_std_logic_vector(4, 8),
43272 => conv_std_logic_vector(5, 8),
43273 => conv_std_logic_vector(5, 8),
43274 => conv_std_logic_vector(6, 8),
43275 => conv_std_logic_vector(7, 8),
43276 => conv_std_logic_vector(7, 8),
43277 => conv_std_logic_vector(8, 8),
43278 => conv_std_logic_vector(9, 8),
43279 => conv_std_logic_vector(9, 8),
43280 => conv_std_logic_vector(10, 8),
43281 => conv_std_logic_vector(11, 8),
43282 => conv_std_logic_vector(11, 8),
43283 => conv_std_logic_vector(12, 8),
43284 => conv_std_logic_vector(13, 8),
43285 => conv_std_logic_vector(13, 8),
43286 => conv_std_logic_vector(14, 8),
43287 => conv_std_logic_vector(15, 8),
43288 => conv_std_logic_vector(15, 8),
43289 => conv_std_logic_vector(16, 8),
43290 => conv_std_logic_vector(17, 8),
43291 => conv_std_logic_vector(17, 8),
43292 => conv_std_logic_vector(18, 8),
43293 => conv_std_logic_vector(19, 8),
43294 => conv_std_logic_vector(19, 8),
43295 => conv_std_logic_vector(20, 8),
43296 => conv_std_logic_vector(21, 8),
43297 => conv_std_logic_vector(21, 8),
43298 => conv_std_logic_vector(22, 8),
43299 => conv_std_logic_vector(23, 8),
43300 => conv_std_logic_vector(23, 8),
43301 => conv_std_logic_vector(24, 8),
43302 => conv_std_logic_vector(25, 8),
43303 => conv_std_logic_vector(25, 8),
43304 => conv_std_logic_vector(26, 8),
43305 => conv_std_logic_vector(27, 8),
43306 => conv_std_logic_vector(27, 8),
43307 => conv_std_logic_vector(28, 8),
43308 => conv_std_logic_vector(29, 8),
43309 => conv_std_logic_vector(29, 8),
43310 => conv_std_logic_vector(30, 8),
43311 => conv_std_logic_vector(31, 8),
43312 => conv_std_logic_vector(31, 8),
43313 => conv_std_logic_vector(32, 8),
43314 => conv_std_logic_vector(33, 8),
43315 => conv_std_logic_vector(33, 8),
43316 => conv_std_logic_vector(34, 8),
43317 => conv_std_logic_vector(34, 8),
43318 => conv_std_logic_vector(35, 8),
43319 => conv_std_logic_vector(36, 8),
43320 => conv_std_logic_vector(36, 8),
43321 => conv_std_logic_vector(37, 8),
43322 => conv_std_logic_vector(38, 8),
43323 => conv_std_logic_vector(38, 8),
43324 => conv_std_logic_vector(39, 8),
43325 => conv_std_logic_vector(40, 8),
43326 => conv_std_logic_vector(40, 8),
43327 => conv_std_logic_vector(41, 8),
43328 => conv_std_logic_vector(42, 8),
43329 => conv_std_logic_vector(42, 8),
43330 => conv_std_logic_vector(43, 8),
43331 => conv_std_logic_vector(44, 8),
43332 => conv_std_logic_vector(44, 8),
43333 => conv_std_logic_vector(45, 8),
43334 => conv_std_logic_vector(46, 8),
43335 => conv_std_logic_vector(46, 8),
43336 => conv_std_logic_vector(47, 8),
43337 => conv_std_logic_vector(48, 8),
43338 => conv_std_logic_vector(48, 8),
43339 => conv_std_logic_vector(49, 8),
43340 => conv_std_logic_vector(50, 8),
43341 => conv_std_logic_vector(50, 8),
43342 => conv_std_logic_vector(51, 8),
43343 => conv_std_logic_vector(52, 8),
43344 => conv_std_logic_vector(52, 8),
43345 => conv_std_logic_vector(53, 8),
43346 => conv_std_logic_vector(54, 8),
43347 => conv_std_logic_vector(54, 8),
43348 => conv_std_logic_vector(55, 8),
43349 => conv_std_logic_vector(56, 8),
43350 => conv_std_logic_vector(56, 8),
43351 => conv_std_logic_vector(57, 8),
43352 => conv_std_logic_vector(58, 8),
43353 => conv_std_logic_vector(58, 8),
43354 => conv_std_logic_vector(59, 8),
43355 => conv_std_logic_vector(60, 8),
43356 => conv_std_logic_vector(60, 8),
43357 => conv_std_logic_vector(61, 8),
43358 => conv_std_logic_vector(62, 8),
43359 => conv_std_logic_vector(62, 8),
43360 => conv_std_logic_vector(63, 8),
43361 => conv_std_logic_vector(64, 8),
43362 => conv_std_logic_vector(64, 8),
43363 => conv_std_logic_vector(65, 8),
43364 => conv_std_logic_vector(66, 8),
43365 => conv_std_logic_vector(66, 8),
43366 => conv_std_logic_vector(67, 8),
43367 => conv_std_logic_vector(67, 8),
43368 => conv_std_logic_vector(68, 8),
43369 => conv_std_logic_vector(69, 8),
43370 => conv_std_logic_vector(69, 8),
43371 => conv_std_logic_vector(70, 8),
43372 => conv_std_logic_vector(71, 8),
43373 => conv_std_logic_vector(71, 8),
43374 => conv_std_logic_vector(72, 8),
43375 => conv_std_logic_vector(73, 8),
43376 => conv_std_logic_vector(73, 8),
43377 => conv_std_logic_vector(74, 8),
43378 => conv_std_logic_vector(75, 8),
43379 => conv_std_logic_vector(75, 8),
43380 => conv_std_logic_vector(76, 8),
43381 => conv_std_logic_vector(77, 8),
43382 => conv_std_logic_vector(77, 8),
43383 => conv_std_logic_vector(78, 8),
43384 => conv_std_logic_vector(79, 8),
43385 => conv_std_logic_vector(79, 8),
43386 => conv_std_logic_vector(80, 8),
43387 => conv_std_logic_vector(81, 8),
43388 => conv_std_logic_vector(81, 8),
43389 => conv_std_logic_vector(82, 8),
43390 => conv_std_logic_vector(83, 8),
43391 => conv_std_logic_vector(83, 8),
43392 => conv_std_logic_vector(84, 8),
43393 => conv_std_logic_vector(85, 8),
43394 => conv_std_logic_vector(85, 8),
43395 => conv_std_logic_vector(86, 8),
43396 => conv_std_logic_vector(87, 8),
43397 => conv_std_logic_vector(87, 8),
43398 => conv_std_logic_vector(88, 8),
43399 => conv_std_logic_vector(89, 8),
43400 => conv_std_logic_vector(89, 8),
43401 => conv_std_logic_vector(90, 8),
43402 => conv_std_logic_vector(91, 8),
43403 => conv_std_logic_vector(91, 8),
43404 => conv_std_logic_vector(92, 8),
43405 => conv_std_logic_vector(93, 8),
43406 => conv_std_logic_vector(93, 8),
43407 => conv_std_logic_vector(94, 8),
43408 => conv_std_logic_vector(95, 8),
43409 => conv_std_logic_vector(95, 8),
43410 => conv_std_logic_vector(96, 8),
43411 => conv_std_logic_vector(97, 8),
43412 => conv_std_logic_vector(97, 8),
43413 => conv_std_logic_vector(98, 8),
43414 => conv_std_logic_vector(99, 8),
43415 => conv_std_logic_vector(99, 8),
43416 => conv_std_logic_vector(100, 8),
43417 => conv_std_logic_vector(101, 8),
43418 => conv_std_logic_vector(101, 8),
43419 => conv_std_logic_vector(102, 8),
43420 => conv_std_logic_vector(102, 8),
43421 => conv_std_logic_vector(103, 8),
43422 => conv_std_logic_vector(104, 8),
43423 => conv_std_logic_vector(104, 8),
43424 => conv_std_logic_vector(105, 8),
43425 => conv_std_logic_vector(106, 8),
43426 => conv_std_logic_vector(106, 8),
43427 => conv_std_logic_vector(107, 8),
43428 => conv_std_logic_vector(108, 8),
43429 => conv_std_logic_vector(108, 8),
43430 => conv_std_logic_vector(109, 8),
43431 => conv_std_logic_vector(110, 8),
43432 => conv_std_logic_vector(110, 8),
43433 => conv_std_logic_vector(111, 8),
43434 => conv_std_logic_vector(112, 8),
43435 => conv_std_logic_vector(112, 8),
43436 => conv_std_logic_vector(113, 8),
43437 => conv_std_logic_vector(114, 8),
43438 => conv_std_logic_vector(114, 8),
43439 => conv_std_logic_vector(115, 8),
43440 => conv_std_logic_vector(116, 8),
43441 => conv_std_logic_vector(116, 8),
43442 => conv_std_logic_vector(117, 8),
43443 => conv_std_logic_vector(118, 8),
43444 => conv_std_logic_vector(118, 8),
43445 => conv_std_logic_vector(119, 8),
43446 => conv_std_logic_vector(120, 8),
43447 => conv_std_logic_vector(120, 8),
43448 => conv_std_logic_vector(121, 8),
43449 => conv_std_logic_vector(122, 8),
43450 => conv_std_logic_vector(122, 8),
43451 => conv_std_logic_vector(123, 8),
43452 => conv_std_logic_vector(124, 8),
43453 => conv_std_logic_vector(124, 8),
43454 => conv_std_logic_vector(125, 8),
43455 => conv_std_logic_vector(126, 8),
43456 => conv_std_logic_vector(126, 8),
43457 => conv_std_logic_vector(127, 8),
43458 => conv_std_logic_vector(128, 8),
43459 => conv_std_logic_vector(128, 8),
43460 => conv_std_logic_vector(129, 8),
43461 => conv_std_logic_vector(130, 8),
43462 => conv_std_logic_vector(130, 8),
43463 => conv_std_logic_vector(131, 8),
43464 => conv_std_logic_vector(132, 8),
43465 => conv_std_logic_vector(132, 8),
43466 => conv_std_logic_vector(133, 8),
43467 => conv_std_logic_vector(134, 8),
43468 => conv_std_logic_vector(134, 8),
43469 => conv_std_logic_vector(135, 8),
43470 => conv_std_logic_vector(135, 8),
43471 => conv_std_logic_vector(136, 8),
43472 => conv_std_logic_vector(137, 8),
43473 => conv_std_logic_vector(137, 8),
43474 => conv_std_logic_vector(138, 8),
43475 => conv_std_logic_vector(139, 8),
43476 => conv_std_logic_vector(139, 8),
43477 => conv_std_logic_vector(140, 8),
43478 => conv_std_logic_vector(141, 8),
43479 => conv_std_logic_vector(141, 8),
43480 => conv_std_logic_vector(142, 8),
43481 => conv_std_logic_vector(143, 8),
43482 => conv_std_logic_vector(143, 8),
43483 => conv_std_logic_vector(144, 8),
43484 => conv_std_logic_vector(145, 8),
43485 => conv_std_logic_vector(145, 8),
43486 => conv_std_logic_vector(146, 8),
43487 => conv_std_logic_vector(147, 8),
43488 => conv_std_logic_vector(147, 8),
43489 => conv_std_logic_vector(148, 8),
43490 => conv_std_logic_vector(149, 8),
43491 => conv_std_logic_vector(149, 8),
43492 => conv_std_logic_vector(150, 8),
43493 => conv_std_logic_vector(151, 8),
43494 => conv_std_logic_vector(151, 8),
43495 => conv_std_logic_vector(152, 8),
43496 => conv_std_logic_vector(153, 8),
43497 => conv_std_logic_vector(153, 8),
43498 => conv_std_logic_vector(154, 8),
43499 => conv_std_logic_vector(155, 8),
43500 => conv_std_logic_vector(155, 8),
43501 => conv_std_logic_vector(156, 8),
43502 => conv_std_logic_vector(157, 8),
43503 => conv_std_logic_vector(157, 8),
43504 => conv_std_logic_vector(158, 8),
43505 => conv_std_logic_vector(159, 8),
43506 => conv_std_logic_vector(159, 8),
43507 => conv_std_logic_vector(160, 8),
43508 => conv_std_logic_vector(161, 8),
43509 => conv_std_logic_vector(161, 8),
43510 => conv_std_logic_vector(162, 8),
43511 => conv_std_logic_vector(163, 8),
43512 => conv_std_logic_vector(163, 8),
43513 => conv_std_logic_vector(164, 8),
43514 => conv_std_logic_vector(165, 8),
43515 => conv_std_logic_vector(165, 8),
43516 => conv_std_logic_vector(166, 8),
43517 => conv_std_logic_vector(167, 8),
43518 => conv_std_logic_vector(167, 8),
43519 => conv_std_logic_vector(168, 8),
43520 => conv_std_logic_vector(0, 8),
43521 => conv_std_logic_vector(0, 8),
43522 => conv_std_logic_vector(1, 8),
43523 => conv_std_logic_vector(1, 8),
43524 => conv_std_logic_vector(2, 8),
43525 => conv_std_logic_vector(3, 8),
43526 => conv_std_logic_vector(3, 8),
43527 => conv_std_logic_vector(4, 8),
43528 => conv_std_logic_vector(5, 8),
43529 => conv_std_logic_vector(5, 8),
43530 => conv_std_logic_vector(6, 8),
43531 => conv_std_logic_vector(7, 8),
43532 => conv_std_logic_vector(7, 8),
43533 => conv_std_logic_vector(8, 8),
43534 => conv_std_logic_vector(9, 8),
43535 => conv_std_logic_vector(9, 8),
43536 => conv_std_logic_vector(10, 8),
43537 => conv_std_logic_vector(11, 8),
43538 => conv_std_logic_vector(11, 8),
43539 => conv_std_logic_vector(12, 8),
43540 => conv_std_logic_vector(13, 8),
43541 => conv_std_logic_vector(13, 8),
43542 => conv_std_logic_vector(14, 8),
43543 => conv_std_logic_vector(15, 8),
43544 => conv_std_logic_vector(15, 8),
43545 => conv_std_logic_vector(16, 8),
43546 => conv_std_logic_vector(17, 8),
43547 => conv_std_logic_vector(17, 8),
43548 => conv_std_logic_vector(18, 8),
43549 => conv_std_logic_vector(19, 8),
43550 => conv_std_logic_vector(19, 8),
43551 => conv_std_logic_vector(20, 8),
43552 => conv_std_logic_vector(21, 8),
43553 => conv_std_logic_vector(21, 8),
43554 => conv_std_logic_vector(22, 8),
43555 => conv_std_logic_vector(23, 8),
43556 => conv_std_logic_vector(23, 8),
43557 => conv_std_logic_vector(24, 8),
43558 => conv_std_logic_vector(25, 8),
43559 => conv_std_logic_vector(25, 8),
43560 => conv_std_logic_vector(26, 8),
43561 => conv_std_logic_vector(27, 8),
43562 => conv_std_logic_vector(27, 8),
43563 => conv_std_logic_vector(28, 8),
43564 => conv_std_logic_vector(29, 8),
43565 => conv_std_logic_vector(29, 8),
43566 => conv_std_logic_vector(30, 8),
43567 => conv_std_logic_vector(31, 8),
43568 => conv_std_logic_vector(31, 8),
43569 => conv_std_logic_vector(32, 8),
43570 => conv_std_logic_vector(33, 8),
43571 => conv_std_logic_vector(33, 8),
43572 => conv_std_logic_vector(34, 8),
43573 => conv_std_logic_vector(35, 8),
43574 => conv_std_logic_vector(35, 8),
43575 => conv_std_logic_vector(36, 8),
43576 => conv_std_logic_vector(37, 8),
43577 => conv_std_logic_vector(37, 8),
43578 => conv_std_logic_vector(38, 8),
43579 => conv_std_logic_vector(39, 8),
43580 => conv_std_logic_vector(39, 8),
43581 => conv_std_logic_vector(40, 8),
43582 => conv_std_logic_vector(41, 8),
43583 => conv_std_logic_vector(41, 8),
43584 => conv_std_logic_vector(42, 8),
43585 => conv_std_logic_vector(43, 8),
43586 => conv_std_logic_vector(43, 8),
43587 => conv_std_logic_vector(44, 8),
43588 => conv_std_logic_vector(45, 8),
43589 => conv_std_logic_vector(45, 8),
43590 => conv_std_logic_vector(46, 8),
43591 => conv_std_logic_vector(47, 8),
43592 => conv_std_logic_vector(47, 8),
43593 => conv_std_logic_vector(48, 8),
43594 => conv_std_logic_vector(49, 8),
43595 => conv_std_logic_vector(49, 8),
43596 => conv_std_logic_vector(50, 8),
43597 => conv_std_logic_vector(51, 8),
43598 => conv_std_logic_vector(51, 8),
43599 => conv_std_logic_vector(52, 8),
43600 => conv_std_logic_vector(53, 8),
43601 => conv_std_logic_vector(53, 8),
43602 => conv_std_logic_vector(54, 8),
43603 => conv_std_logic_vector(55, 8),
43604 => conv_std_logic_vector(55, 8),
43605 => conv_std_logic_vector(56, 8),
43606 => conv_std_logic_vector(57, 8),
43607 => conv_std_logic_vector(57, 8),
43608 => conv_std_logic_vector(58, 8),
43609 => conv_std_logic_vector(59, 8),
43610 => conv_std_logic_vector(59, 8),
43611 => conv_std_logic_vector(60, 8),
43612 => conv_std_logic_vector(61, 8),
43613 => conv_std_logic_vector(61, 8),
43614 => conv_std_logic_vector(62, 8),
43615 => conv_std_logic_vector(63, 8),
43616 => conv_std_logic_vector(63, 8),
43617 => conv_std_logic_vector(64, 8),
43618 => conv_std_logic_vector(65, 8),
43619 => conv_std_logic_vector(65, 8),
43620 => conv_std_logic_vector(66, 8),
43621 => conv_std_logic_vector(67, 8),
43622 => conv_std_logic_vector(67, 8),
43623 => conv_std_logic_vector(68, 8),
43624 => conv_std_logic_vector(69, 8),
43625 => conv_std_logic_vector(69, 8),
43626 => conv_std_logic_vector(70, 8),
43627 => conv_std_logic_vector(71, 8),
43628 => conv_std_logic_vector(71, 8),
43629 => conv_std_logic_vector(72, 8),
43630 => conv_std_logic_vector(73, 8),
43631 => conv_std_logic_vector(73, 8),
43632 => conv_std_logic_vector(74, 8),
43633 => conv_std_logic_vector(75, 8),
43634 => conv_std_logic_vector(75, 8),
43635 => conv_std_logic_vector(76, 8),
43636 => conv_std_logic_vector(77, 8),
43637 => conv_std_logic_vector(77, 8),
43638 => conv_std_logic_vector(78, 8),
43639 => conv_std_logic_vector(79, 8),
43640 => conv_std_logic_vector(79, 8),
43641 => conv_std_logic_vector(80, 8),
43642 => conv_std_logic_vector(81, 8),
43643 => conv_std_logic_vector(81, 8),
43644 => conv_std_logic_vector(82, 8),
43645 => conv_std_logic_vector(83, 8),
43646 => conv_std_logic_vector(83, 8),
43647 => conv_std_logic_vector(84, 8),
43648 => conv_std_logic_vector(85, 8),
43649 => conv_std_logic_vector(85, 8),
43650 => conv_std_logic_vector(86, 8),
43651 => conv_std_logic_vector(86, 8),
43652 => conv_std_logic_vector(87, 8),
43653 => conv_std_logic_vector(88, 8),
43654 => conv_std_logic_vector(88, 8),
43655 => conv_std_logic_vector(89, 8),
43656 => conv_std_logic_vector(90, 8),
43657 => conv_std_logic_vector(90, 8),
43658 => conv_std_logic_vector(91, 8),
43659 => conv_std_logic_vector(92, 8),
43660 => conv_std_logic_vector(92, 8),
43661 => conv_std_logic_vector(93, 8),
43662 => conv_std_logic_vector(94, 8),
43663 => conv_std_logic_vector(94, 8),
43664 => conv_std_logic_vector(95, 8),
43665 => conv_std_logic_vector(96, 8),
43666 => conv_std_logic_vector(96, 8),
43667 => conv_std_logic_vector(97, 8),
43668 => conv_std_logic_vector(98, 8),
43669 => conv_std_logic_vector(98, 8),
43670 => conv_std_logic_vector(99, 8),
43671 => conv_std_logic_vector(100, 8),
43672 => conv_std_logic_vector(100, 8),
43673 => conv_std_logic_vector(101, 8),
43674 => conv_std_logic_vector(102, 8),
43675 => conv_std_logic_vector(102, 8),
43676 => conv_std_logic_vector(103, 8),
43677 => conv_std_logic_vector(104, 8),
43678 => conv_std_logic_vector(104, 8),
43679 => conv_std_logic_vector(105, 8),
43680 => conv_std_logic_vector(106, 8),
43681 => conv_std_logic_vector(106, 8),
43682 => conv_std_logic_vector(107, 8),
43683 => conv_std_logic_vector(108, 8),
43684 => conv_std_logic_vector(108, 8),
43685 => conv_std_logic_vector(109, 8),
43686 => conv_std_logic_vector(110, 8),
43687 => conv_std_logic_vector(110, 8),
43688 => conv_std_logic_vector(111, 8),
43689 => conv_std_logic_vector(112, 8),
43690 => conv_std_logic_vector(112, 8),
43691 => conv_std_logic_vector(113, 8),
43692 => conv_std_logic_vector(114, 8),
43693 => conv_std_logic_vector(114, 8),
43694 => conv_std_logic_vector(115, 8),
43695 => conv_std_logic_vector(116, 8),
43696 => conv_std_logic_vector(116, 8),
43697 => conv_std_logic_vector(117, 8),
43698 => conv_std_logic_vector(118, 8),
43699 => conv_std_logic_vector(118, 8),
43700 => conv_std_logic_vector(119, 8),
43701 => conv_std_logic_vector(120, 8),
43702 => conv_std_logic_vector(120, 8),
43703 => conv_std_logic_vector(121, 8),
43704 => conv_std_logic_vector(122, 8),
43705 => conv_std_logic_vector(122, 8),
43706 => conv_std_logic_vector(123, 8),
43707 => conv_std_logic_vector(124, 8),
43708 => conv_std_logic_vector(124, 8),
43709 => conv_std_logic_vector(125, 8),
43710 => conv_std_logic_vector(126, 8),
43711 => conv_std_logic_vector(126, 8),
43712 => conv_std_logic_vector(127, 8),
43713 => conv_std_logic_vector(128, 8),
43714 => conv_std_logic_vector(128, 8),
43715 => conv_std_logic_vector(129, 8),
43716 => conv_std_logic_vector(130, 8),
43717 => conv_std_logic_vector(130, 8),
43718 => conv_std_logic_vector(131, 8),
43719 => conv_std_logic_vector(132, 8),
43720 => conv_std_logic_vector(132, 8),
43721 => conv_std_logic_vector(133, 8),
43722 => conv_std_logic_vector(134, 8),
43723 => conv_std_logic_vector(134, 8),
43724 => conv_std_logic_vector(135, 8),
43725 => conv_std_logic_vector(136, 8),
43726 => conv_std_logic_vector(136, 8),
43727 => conv_std_logic_vector(137, 8),
43728 => conv_std_logic_vector(138, 8),
43729 => conv_std_logic_vector(138, 8),
43730 => conv_std_logic_vector(139, 8),
43731 => conv_std_logic_vector(140, 8),
43732 => conv_std_logic_vector(140, 8),
43733 => conv_std_logic_vector(141, 8),
43734 => conv_std_logic_vector(142, 8),
43735 => conv_std_logic_vector(142, 8),
43736 => conv_std_logic_vector(143, 8),
43737 => conv_std_logic_vector(144, 8),
43738 => conv_std_logic_vector(144, 8),
43739 => conv_std_logic_vector(145, 8),
43740 => conv_std_logic_vector(146, 8),
43741 => conv_std_logic_vector(146, 8),
43742 => conv_std_logic_vector(147, 8),
43743 => conv_std_logic_vector(148, 8),
43744 => conv_std_logic_vector(148, 8),
43745 => conv_std_logic_vector(149, 8),
43746 => conv_std_logic_vector(150, 8),
43747 => conv_std_logic_vector(150, 8),
43748 => conv_std_logic_vector(151, 8),
43749 => conv_std_logic_vector(152, 8),
43750 => conv_std_logic_vector(152, 8),
43751 => conv_std_logic_vector(153, 8),
43752 => conv_std_logic_vector(154, 8),
43753 => conv_std_logic_vector(154, 8),
43754 => conv_std_logic_vector(155, 8),
43755 => conv_std_logic_vector(156, 8),
43756 => conv_std_logic_vector(156, 8),
43757 => conv_std_logic_vector(157, 8),
43758 => conv_std_logic_vector(158, 8),
43759 => conv_std_logic_vector(158, 8),
43760 => conv_std_logic_vector(159, 8),
43761 => conv_std_logic_vector(160, 8),
43762 => conv_std_logic_vector(160, 8),
43763 => conv_std_logic_vector(161, 8),
43764 => conv_std_logic_vector(162, 8),
43765 => conv_std_logic_vector(162, 8),
43766 => conv_std_logic_vector(163, 8),
43767 => conv_std_logic_vector(164, 8),
43768 => conv_std_logic_vector(164, 8),
43769 => conv_std_logic_vector(165, 8),
43770 => conv_std_logic_vector(166, 8),
43771 => conv_std_logic_vector(166, 8),
43772 => conv_std_logic_vector(167, 8),
43773 => conv_std_logic_vector(168, 8),
43774 => conv_std_logic_vector(168, 8),
43775 => conv_std_logic_vector(169, 8),
43776 => conv_std_logic_vector(0, 8),
43777 => conv_std_logic_vector(0, 8),
43778 => conv_std_logic_vector(1, 8),
43779 => conv_std_logic_vector(2, 8),
43780 => conv_std_logic_vector(2, 8),
43781 => conv_std_logic_vector(3, 8),
43782 => conv_std_logic_vector(4, 8),
43783 => conv_std_logic_vector(4, 8),
43784 => conv_std_logic_vector(5, 8),
43785 => conv_std_logic_vector(6, 8),
43786 => conv_std_logic_vector(6, 8),
43787 => conv_std_logic_vector(7, 8),
43788 => conv_std_logic_vector(8, 8),
43789 => conv_std_logic_vector(8, 8),
43790 => conv_std_logic_vector(9, 8),
43791 => conv_std_logic_vector(10, 8),
43792 => conv_std_logic_vector(10, 8),
43793 => conv_std_logic_vector(11, 8),
43794 => conv_std_logic_vector(12, 8),
43795 => conv_std_logic_vector(12, 8),
43796 => conv_std_logic_vector(13, 8),
43797 => conv_std_logic_vector(14, 8),
43798 => conv_std_logic_vector(14, 8),
43799 => conv_std_logic_vector(15, 8),
43800 => conv_std_logic_vector(16, 8),
43801 => conv_std_logic_vector(16, 8),
43802 => conv_std_logic_vector(17, 8),
43803 => conv_std_logic_vector(18, 8),
43804 => conv_std_logic_vector(18, 8),
43805 => conv_std_logic_vector(19, 8),
43806 => conv_std_logic_vector(20, 8),
43807 => conv_std_logic_vector(20, 8),
43808 => conv_std_logic_vector(21, 8),
43809 => conv_std_logic_vector(22, 8),
43810 => conv_std_logic_vector(22, 8),
43811 => conv_std_logic_vector(23, 8),
43812 => conv_std_logic_vector(24, 8),
43813 => conv_std_logic_vector(24, 8),
43814 => conv_std_logic_vector(25, 8),
43815 => conv_std_logic_vector(26, 8),
43816 => conv_std_logic_vector(26, 8),
43817 => conv_std_logic_vector(27, 8),
43818 => conv_std_logic_vector(28, 8),
43819 => conv_std_logic_vector(28, 8),
43820 => conv_std_logic_vector(29, 8),
43821 => conv_std_logic_vector(30, 8),
43822 => conv_std_logic_vector(30, 8),
43823 => conv_std_logic_vector(31, 8),
43824 => conv_std_logic_vector(32, 8),
43825 => conv_std_logic_vector(32, 8),
43826 => conv_std_logic_vector(33, 8),
43827 => conv_std_logic_vector(34, 8),
43828 => conv_std_logic_vector(34, 8),
43829 => conv_std_logic_vector(35, 8),
43830 => conv_std_logic_vector(36, 8),
43831 => conv_std_logic_vector(36, 8),
43832 => conv_std_logic_vector(37, 8),
43833 => conv_std_logic_vector(38, 8),
43834 => conv_std_logic_vector(38, 8),
43835 => conv_std_logic_vector(39, 8),
43836 => conv_std_logic_vector(40, 8),
43837 => conv_std_logic_vector(40, 8),
43838 => conv_std_logic_vector(41, 8),
43839 => conv_std_logic_vector(42, 8),
43840 => conv_std_logic_vector(42, 8),
43841 => conv_std_logic_vector(43, 8),
43842 => conv_std_logic_vector(44, 8),
43843 => conv_std_logic_vector(44, 8),
43844 => conv_std_logic_vector(45, 8),
43845 => conv_std_logic_vector(46, 8),
43846 => conv_std_logic_vector(46, 8),
43847 => conv_std_logic_vector(47, 8),
43848 => conv_std_logic_vector(48, 8),
43849 => conv_std_logic_vector(48, 8),
43850 => conv_std_logic_vector(49, 8),
43851 => conv_std_logic_vector(50, 8),
43852 => conv_std_logic_vector(50, 8),
43853 => conv_std_logic_vector(51, 8),
43854 => conv_std_logic_vector(52, 8),
43855 => conv_std_logic_vector(52, 8),
43856 => conv_std_logic_vector(53, 8),
43857 => conv_std_logic_vector(54, 8),
43858 => conv_std_logic_vector(54, 8),
43859 => conv_std_logic_vector(55, 8),
43860 => conv_std_logic_vector(56, 8),
43861 => conv_std_logic_vector(56, 8),
43862 => conv_std_logic_vector(57, 8),
43863 => conv_std_logic_vector(58, 8),
43864 => conv_std_logic_vector(58, 8),
43865 => conv_std_logic_vector(59, 8),
43866 => conv_std_logic_vector(60, 8),
43867 => conv_std_logic_vector(60, 8),
43868 => conv_std_logic_vector(61, 8),
43869 => conv_std_logic_vector(62, 8),
43870 => conv_std_logic_vector(62, 8),
43871 => conv_std_logic_vector(63, 8),
43872 => conv_std_logic_vector(64, 8),
43873 => conv_std_logic_vector(64, 8),
43874 => conv_std_logic_vector(65, 8),
43875 => conv_std_logic_vector(66, 8),
43876 => conv_std_logic_vector(66, 8),
43877 => conv_std_logic_vector(67, 8),
43878 => conv_std_logic_vector(68, 8),
43879 => conv_std_logic_vector(68, 8),
43880 => conv_std_logic_vector(69, 8),
43881 => conv_std_logic_vector(70, 8),
43882 => conv_std_logic_vector(70, 8),
43883 => conv_std_logic_vector(71, 8),
43884 => conv_std_logic_vector(72, 8),
43885 => conv_std_logic_vector(72, 8),
43886 => conv_std_logic_vector(73, 8),
43887 => conv_std_logic_vector(74, 8),
43888 => conv_std_logic_vector(74, 8),
43889 => conv_std_logic_vector(75, 8),
43890 => conv_std_logic_vector(76, 8),
43891 => conv_std_logic_vector(76, 8),
43892 => conv_std_logic_vector(77, 8),
43893 => conv_std_logic_vector(78, 8),
43894 => conv_std_logic_vector(78, 8),
43895 => conv_std_logic_vector(79, 8),
43896 => conv_std_logic_vector(80, 8),
43897 => conv_std_logic_vector(80, 8),
43898 => conv_std_logic_vector(81, 8),
43899 => conv_std_logic_vector(82, 8),
43900 => conv_std_logic_vector(82, 8),
43901 => conv_std_logic_vector(83, 8),
43902 => conv_std_logic_vector(84, 8),
43903 => conv_std_logic_vector(84, 8),
43904 => conv_std_logic_vector(85, 8),
43905 => conv_std_logic_vector(86, 8),
43906 => conv_std_logic_vector(86, 8),
43907 => conv_std_logic_vector(87, 8),
43908 => conv_std_logic_vector(88, 8),
43909 => conv_std_logic_vector(88, 8),
43910 => conv_std_logic_vector(89, 8),
43911 => conv_std_logic_vector(90, 8),
43912 => conv_std_logic_vector(90, 8),
43913 => conv_std_logic_vector(91, 8),
43914 => conv_std_logic_vector(92, 8),
43915 => conv_std_logic_vector(92, 8),
43916 => conv_std_logic_vector(93, 8),
43917 => conv_std_logic_vector(94, 8),
43918 => conv_std_logic_vector(94, 8),
43919 => conv_std_logic_vector(95, 8),
43920 => conv_std_logic_vector(96, 8),
43921 => conv_std_logic_vector(96, 8),
43922 => conv_std_logic_vector(97, 8),
43923 => conv_std_logic_vector(98, 8),
43924 => conv_std_logic_vector(98, 8),
43925 => conv_std_logic_vector(99, 8),
43926 => conv_std_logic_vector(100, 8),
43927 => conv_std_logic_vector(100, 8),
43928 => conv_std_logic_vector(101, 8),
43929 => conv_std_logic_vector(102, 8),
43930 => conv_std_logic_vector(102, 8),
43931 => conv_std_logic_vector(103, 8),
43932 => conv_std_logic_vector(104, 8),
43933 => conv_std_logic_vector(104, 8),
43934 => conv_std_logic_vector(105, 8),
43935 => conv_std_logic_vector(106, 8),
43936 => conv_std_logic_vector(106, 8),
43937 => conv_std_logic_vector(107, 8),
43938 => conv_std_logic_vector(108, 8),
43939 => conv_std_logic_vector(108, 8),
43940 => conv_std_logic_vector(109, 8),
43941 => conv_std_logic_vector(110, 8),
43942 => conv_std_logic_vector(110, 8),
43943 => conv_std_logic_vector(111, 8),
43944 => conv_std_logic_vector(112, 8),
43945 => conv_std_logic_vector(112, 8),
43946 => conv_std_logic_vector(113, 8),
43947 => conv_std_logic_vector(114, 8),
43948 => conv_std_logic_vector(114, 8),
43949 => conv_std_logic_vector(115, 8),
43950 => conv_std_logic_vector(116, 8),
43951 => conv_std_logic_vector(116, 8),
43952 => conv_std_logic_vector(117, 8),
43953 => conv_std_logic_vector(118, 8),
43954 => conv_std_logic_vector(118, 8),
43955 => conv_std_logic_vector(119, 8),
43956 => conv_std_logic_vector(120, 8),
43957 => conv_std_logic_vector(120, 8),
43958 => conv_std_logic_vector(121, 8),
43959 => conv_std_logic_vector(122, 8),
43960 => conv_std_logic_vector(122, 8),
43961 => conv_std_logic_vector(123, 8),
43962 => conv_std_logic_vector(124, 8),
43963 => conv_std_logic_vector(124, 8),
43964 => conv_std_logic_vector(125, 8),
43965 => conv_std_logic_vector(126, 8),
43966 => conv_std_logic_vector(126, 8),
43967 => conv_std_logic_vector(127, 8),
43968 => conv_std_logic_vector(128, 8),
43969 => conv_std_logic_vector(128, 8),
43970 => conv_std_logic_vector(129, 8),
43971 => conv_std_logic_vector(130, 8),
43972 => conv_std_logic_vector(130, 8),
43973 => conv_std_logic_vector(131, 8),
43974 => conv_std_logic_vector(132, 8),
43975 => conv_std_logic_vector(132, 8),
43976 => conv_std_logic_vector(133, 8),
43977 => conv_std_logic_vector(134, 8),
43978 => conv_std_logic_vector(134, 8),
43979 => conv_std_logic_vector(135, 8),
43980 => conv_std_logic_vector(136, 8),
43981 => conv_std_logic_vector(136, 8),
43982 => conv_std_logic_vector(137, 8),
43983 => conv_std_logic_vector(138, 8),
43984 => conv_std_logic_vector(138, 8),
43985 => conv_std_logic_vector(139, 8),
43986 => conv_std_logic_vector(140, 8),
43987 => conv_std_logic_vector(140, 8),
43988 => conv_std_logic_vector(141, 8),
43989 => conv_std_logic_vector(142, 8),
43990 => conv_std_logic_vector(142, 8),
43991 => conv_std_logic_vector(143, 8),
43992 => conv_std_logic_vector(144, 8),
43993 => conv_std_logic_vector(144, 8),
43994 => conv_std_logic_vector(145, 8),
43995 => conv_std_logic_vector(146, 8),
43996 => conv_std_logic_vector(146, 8),
43997 => conv_std_logic_vector(147, 8),
43998 => conv_std_logic_vector(148, 8),
43999 => conv_std_logic_vector(148, 8),
44000 => conv_std_logic_vector(149, 8),
44001 => conv_std_logic_vector(150, 8),
44002 => conv_std_logic_vector(150, 8),
44003 => conv_std_logic_vector(151, 8),
44004 => conv_std_logic_vector(152, 8),
44005 => conv_std_logic_vector(152, 8),
44006 => conv_std_logic_vector(153, 8),
44007 => conv_std_logic_vector(154, 8),
44008 => conv_std_logic_vector(154, 8),
44009 => conv_std_logic_vector(155, 8),
44010 => conv_std_logic_vector(156, 8),
44011 => conv_std_logic_vector(156, 8),
44012 => conv_std_logic_vector(157, 8),
44013 => conv_std_logic_vector(158, 8),
44014 => conv_std_logic_vector(158, 8),
44015 => conv_std_logic_vector(159, 8),
44016 => conv_std_logic_vector(160, 8),
44017 => conv_std_logic_vector(160, 8),
44018 => conv_std_logic_vector(161, 8),
44019 => conv_std_logic_vector(162, 8),
44020 => conv_std_logic_vector(162, 8),
44021 => conv_std_logic_vector(163, 8),
44022 => conv_std_logic_vector(164, 8),
44023 => conv_std_logic_vector(164, 8),
44024 => conv_std_logic_vector(165, 8),
44025 => conv_std_logic_vector(166, 8),
44026 => conv_std_logic_vector(166, 8),
44027 => conv_std_logic_vector(167, 8),
44028 => conv_std_logic_vector(168, 8),
44029 => conv_std_logic_vector(168, 8),
44030 => conv_std_logic_vector(169, 8),
44031 => conv_std_logic_vector(170, 8),
44032 => conv_std_logic_vector(0, 8),
44033 => conv_std_logic_vector(0, 8),
44034 => conv_std_logic_vector(1, 8),
44035 => conv_std_logic_vector(2, 8),
44036 => conv_std_logic_vector(2, 8),
44037 => conv_std_logic_vector(3, 8),
44038 => conv_std_logic_vector(4, 8),
44039 => conv_std_logic_vector(4, 8),
44040 => conv_std_logic_vector(5, 8),
44041 => conv_std_logic_vector(6, 8),
44042 => conv_std_logic_vector(6, 8),
44043 => conv_std_logic_vector(7, 8),
44044 => conv_std_logic_vector(8, 8),
44045 => conv_std_logic_vector(8, 8),
44046 => conv_std_logic_vector(9, 8),
44047 => conv_std_logic_vector(10, 8),
44048 => conv_std_logic_vector(10, 8),
44049 => conv_std_logic_vector(11, 8),
44050 => conv_std_logic_vector(12, 8),
44051 => conv_std_logic_vector(12, 8),
44052 => conv_std_logic_vector(13, 8),
44053 => conv_std_logic_vector(14, 8),
44054 => conv_std_logic_vector(14, 8),
44055 => conv_std_logic_vector(15, 8),
44056 => conv_std_logic_vector(16, 8),
44057 => conv_std_logic_vector(16, 8),
44058 => conv_std_logic_vector(17, 8),
44059 => conv_std_logic_vector(18, 8),
44060 => conv_std_logic_vector(18, 8),
44061 => conv_std_logic_vector(19, 8),
44062 => conv_std_logic_vector(20, 8),
44063 => conv_std_logic_vector(20, 8),
44064 => conv_std_logic_vector(21, 8),
44065 => conv_std_logic_vector(22, 8),
44066 => conv_std_logic_vector(22, 8),
44067 => conv_std_logic_vector(23, 8),
44068 => conv_std_logic_vector(24, 8),
44069 => conv_std_logic_vector(24, 8),
44070 => conv_std_logic_vector(25, 8),
44071 => conv_std_logic_vector(26, 8),
44072 => conv_std_logic_vector(26, 8),
44073 => conv_std_logic_vector(27, 8),
44074 => conv_std_logic_vector(28, 8),
44075 => conv_std_logic_vector(28, 8),
44076 => conv_std_logic_vector(29, 8),
44077 => conv_std_logic_vector(30, 8),
44078 => conv_std_logic_vector(30, 8),
44079 => conv_std_logic_vector(31, 8),
44080 => conv_std_logic_vector(32, 8),
44081 => conv_std_logic_vector(32, 8),
44082 => conv_std_logic_vector(33, 8),
44083 => conv_std_logic_vector(34, 8),
44084 => conv_std_logic_vector(34, 8),
44085 => conv_std_logic_vector(35, 8),
44086 => conv_std_logic_vector(36, 8),
44087 => conv_std_logic_vector(36, 8),
44088 => conv_std_logic_vector(37, 8),
44089 => conv_std_logic_vector(38, 8),
44090 => conv_std_logic_vector(38, 8),
44091 => conv_std_logic_vector(39, 8),
44092 => conv_std_logic_vector(40, 8),
44093 => conv_std_logic_vector(40, 8),
44094 => conv_std_logic_vector(41, 8),
44095 => conv_std_logic_vector(42, 8),
44096 => conv_std_logic_vector(43, 8),
44097 => conv_std_logic_vector(43, 8),
44098 => conv_std_logic_vector(44, 8),
44099 => conv_std_logic_vector(45, 8),
44100 => conv_std_logic_vector(45, 8),
44101 => conv_std_logic_vector(46, 8),
44102 => conv_std_logic_vector(47, 8),
44103 => conv_std_logic_vector(47, 8),
44104 => conv_std_logic_vector(48, 8),
44105 => conv_std_logic_vector(49, 8),
44106 => conv_std_logic_vector(49, 8),
44107 => conv_std_logic_vector(50, 8),
44108 => conv_std_logic_vector(51, 8),
44109 => conv_std_logic_vector(51, 8),
44110 => conv_std_logic_vector(52, 8),
44111 => conv_std_logic_vector(53, 8),
44112 => conv_std_logic_vector(53, 8),
44113 => conv_std_logic_vector(54, 8),
44114 => conv_std_logic_vector(55, 8),
44115 => conv_std_logic_vector(55, 8),
44116 => conv_std_logic_vector(56, 8),
44117 => conv_std_logic_vector(57, 8),
44118 => conv_std_logic_vector(57, 8),
44119 => conv_std_logic_vector(58, 8),
44120 => conv_std_logic_vector(59, 8),
44121 => conv_std_logic_vector(59, 8),
44122 => conv_std_logic_vector(60, 8),
44123 => conv_std_logic_vector(61, 8),
44124 => conv_std_logic_vector(61, 8),
44125 => conv_std_logic_vector(62, 8),
44126 => conv_std_logic_vector(63, 8),
44127 => conv_std_logic_vector(63, 8),
44128 => conv_std_logic_vector(64, 8),
44129 => conv_std_logic_vector(65, 8),
44130 => conv_std_logic_vector(65, 8),
44131 => conv_std_logic_vector(66, 8),
44132 => conv_std_logic_vector(67, 8),
44133 => conv_std_logic_vector(67, 8),
44134 => conv_std_logic_vector(68, 8),
44135 => conv_std_logic_vector(69, 8),
44136 => conv_std_logic_vector(69, 8),
44137 => conv_std_logic_vector(70, 8),
44138 => conv_std_logic_vector(71, 8),
44139 => conv_std_logic_vector(71, 8),
44140 => conv_std_logic_vector(72, 8),
44141 => conv_std_logic_vector(73, 8),
44142 => conv_std_logic_vector(73, 8),
44143 => conv_std_logic_vector(74, 8),
44144 => conv_std_logic_vector(75, 8),
44145 => conv_std_logic_vector(75, 8),
44146 => conv_std_logic_vector(76, 8),
44147 => conv_std_logic_vector(77, 8),
44148 => conv_std_logic_vector(77, 8),
44149 => conv_std_logic_vector(78, 8),
44150 => conv_std_logic_vector(79, 8),
44151 => conv_std_logic_vector(79, 8),
44152 => conv_std_logic_vector(80, 8),
44153 => conv_std_logic_vector(81, 8),
44154 => conv_std_logic_vector(81, 8),
44155 => conv_std_logic_vector(82, 8),
44156 => conv_std_logic_vector(83, 8),
44157 => conv_std_logic_vector(83, 8),
44158 => conv_std_logic_vector(84, 8),
44159 => conv_std_logic_vector(85, 8),
44160 => conv_std_logic_vector(86, 8),
44161 => conv_std_logic_vector(86, 8),
44162 => conv_std_logic_vector(87, 8),
44163 => conv_std_logic_vector(88, 8),
44164 => conv_std_logic_vector(88, 8),
44165 => conv_std_logic_vector(89, 8),
44166 => conv_std_logic_vector(90, 8),
44167 => conv_std_logic_vector(90, 8),
44168 => conv_std_logic_vector(91, 8),
44169 => conv_std_logic_vector(92, 8),
44170 => conv_std_logic_vector(92, 8),
44171 => conv_std_logic_vector(93, 8),
44172 => conv_std_logic_vector(94, 8),
44173 => conv_std_logic_vector(94, 8),
44174 => conv_std_logic_vector(95, 8),
44175 => conv_std_logic_vector(96, 8),
44176 => conv_std_logic_vector(96, 8),
44177 => conv_std_logic_vector(97, 8),
44178 => conv_std_logic_vector(98, 8),
44179 => conv_std_logic_vector(98, 8),
44180 => conv_std_logic_vector(99, 8),
44181 => conv_std_logic_vector(100, 8),
44182 => conv_std_logic_vector(100, 8),
44183 => conv_std_logic_vector(101, 8),
44184 => conv_std_logic_vector(102, 8),
44185 => conv_std_logic_vector(102, 8),
44186 => conv_std_logic_vector(103, 8),
44187 => conv_std_logic_vector(104, 8),
44188 => conv_std_logic_vector(104, 8),
44189 => conv_std_logic_vector(105, 8),
44190 => conv_std_logic_vector(106, 8),
44191 => conv_std_logic_vector(106, 8),
44192 => conv_std_logic_vector(107, 8),
44193 => conv_std_logic_vector(108, 8),
44194 => conv_std_logic_vector(108, 8),
44195 => conv_std_logic_vector(109, 8),
44196 => conv_std_logic_vector(110, 8),
44197 => conv_std_logic_vector(110, 8),
44198 => conv_std_logic_vector(111, 8),
44199 => conv_std_logic_vector(112, 8),
44200 => conv_std_logic_vector(112, 8),
44201 => conv_std_logic_vector(113, 8),
44202 => conv_std_logic_vector(114, 8),
44203 => conv_std_logic_vector(114, 8),
44204 => conv_std_logic_vector(115, 8),
44205 => conv_std_logic_vector(116, 8),
44206 => conv_std_logic_vector(116, 8),
44207 => conv_std_logic_vector(117, 8),
44208 => conv_std_logic_vector(118, 8),
44209 => conv_std_logic_vector(118, 8),
44210 => conv_std_logic_vector(119, 8),
44211 => conv_std_logic_vector(120, 8),
44212 => conv_std_logic_vector(120, 8),
44213 => conv_std_logic_vector(121, 8),
44214 => conv_std_logic_vector(122, 8),
44215 => conv_std_logic_vector(122, 8),
44216 => conv_std_logic_vector(123, 8),
44217 => conv_std_logic_vector(124, 8),
44218 => conv_std_logic_vector(124, 8),
44219 => conv_std_logic_vector(125, 8),
44220 => conv_std_logic_vector(126, 8),
44221 => conv_std_logic_vector(126, 8),
44222 => conv_std_logic_vector(127, 8),
44223 => conv_std_logic_vector(128, 8),
44224 => conv_std_logic_vector(129, 8),
44225 => conv_std_logic_vector(129, 8),
44226 => conv_std_logic_vector(130, 8),
44227 => conv_std_logic_vector(131, 8),
44228 => conv_std_logic_vector(131, 8),
44229 => conv_std_logic_vector(132, 8),
44230 => conv_std_logic_vector(133, 8),
44231 => conv_std_logic_vector(133, 8),
44232 => conv_std_logic_vector(134, 8),
44233 => conv_std_logic_vector(135, 8),
44234 => conv_std_logic_vector(135, 8),
44235 => conv_std_logic_vector(136, 8),
44236 => conv_std_logic_vector(137, 8),
44237 => conv_std_logic_vector(137, 8),
44238 => conv_std_logic_vector(138, 8),
44239 => conv_std_logic_vector(139, 8),
44240 => conv_std_logic_vector(139, 8),
44241 => conv_std_logic_vector(140, 8),
44242 => conv_std_logic_vector(141, 8),
44243 => conv_std_logic_vector(141, 8),
44244 => conv_std_logic_vector(142, 8),
44245 => conv_std_logic_vector(143, 8),
44246 => conv_std_logic_vector(143, 8),
44247 => conv_std_logic_vector(144, 8),
44248 => conv_std_logic_vector(145, 8),
44249 => conv_std_logic_vector(145, 8),
44250 => conv_std_logic_vector(146, 8),
44251 => conv_std_logic_vector(147, 8),
44252 => conv_std_logic_vector(147, 8),
44253 => conv_std_logic_vector(148, 8),
44254 => conv_std_logic_vector(149, 8),
44255 => conv_std_logic_vector(149, 8),
44256 => conv_std_logic_vector(150, 8),
44257 => conv_std_logic_vector(151, 8),
44258 => conv_std_logic_vector(151, 8),
44259 => conv_std_logic_vector(152, 8),
44260 => conv_std_logic_vector(153, 8),
44261 => conv_std_logic_vector(153, 8),
44262 => conv_std_logic_vector(154, 8),
44263 => conv_std_logic_vector(155, 8),
44264 => conv_std_logic_vector(155, 8),
44265 => conv_std_logic_vector(156, 8),
44266 => conv_std_logic_vector(157, 8),
44267 => conv_std_logic_vector(157, 8),
44268 => conv_std_logic_vector(158, 8),
44269 => conv_std_logic_vector(159, 8),
44270 => conv_std_logic_vector(159, 8),
44271 => conv_std_logic_vector(160, 8),
44272 => conv_std_logic_vector(161, 8),
44273 => conv_std_logic_vector(161, 8),
44274 => conv_std_logic_vector(162, 8),
44275 => conv_std_logic_vector(163, 8),
44276 => conv_std_logic_vector(163, 8),
44277 => conv_std_logic_vector(164, 8),
44278 => conv_std_logic_vector(165, 8),
44279 => conv_std_logic_vector(165, 8),
44280 => conv_std_logic_vector(166, 8),
44281 => conv_std_logic_vector(167, 8),
44282 => conv_std_logic_vector(167, 8),
44283 => conv_std_logic_vector(168, 8),
44284 => conv_std_logic_vector(169, 8),
44285 => conv_std_logic_vector(169, 8),
44286 => conv_std_logic_vector(170, 8),
44287 => conv_std_logic_vector(171, 8),
44288 => conv_std_logic_vector(0, 8),
44289 => conv_std_logic_vector(0, 8),
44290 => conv_std_logic_vector(1, 8),
44291 => conv_std_logic_vector(2, 8),
44292 => conv_std_logic_vector(2, 8),
44293 => conv_std_logic_vector(3, 8),
44294 => conv_std_logic_vector(4, 8),
44295 => conv_std_logic_vector(4, 8),
44296 => conv_std_logic_vector(5, 8),
44297 => conv_std_logic_vector(6, 8),
44298 => conv_std_logic_vector(6, 8),
44299 => conv_std_logic_vector(7, 8),
44300 => conv_std_logic_vector(8, 8),
44301 => conv_std_logic_vector(8, 8),
44302 => conv_std_logic_vector(9, 8),
44303 => conv_std_logic_vector(10, 8),
44304 => conv_std_logic_vector(10, 8),
44305 => conv_std_logic_vector(11, 8),
44306 => conv_std_logic_vector(12, 8),
44307 => conv_std_logic_vector(12, 8),
44308 => conv_std_logic_vector(13, 8),
44309 => conv_std_logic_vector(14, 8),
44310 => conv_std_logic_vector(14, 8),
44311 => conv_std_logic_vector(15, 8),
44312 => conv_std_logic_vector(16, 8),
44313 => conv_std_logic_vector(16, 8),
44314 => conv_std_logic_vector(17, 8),
44315 => conv_std_logic_vector(18, 8),
44316 => conv_std_logic_vector(18, 8),
44317 => conv_std_logic_vector(19, 8),
44318 => conv_std_logic_vector(20, 8),
44319 => conv_std_logic_vector(20, 8),
44320 => conv_std_logic_vector(21, 8),
44321 => conv_std_logic_vector(22, 8),
44322 => conv_std_logic_vector(22, 8),
44323 => conv_std_logic_vector(23, 8),
44324 => conv_std_logic_vector(24, 8),
44325 => conv_std_logic_vector(25, 8),
44326 => conv_std_logic_vector(25, 8),
44327 => conv_std_logic_vector(26, 8),
44328 => conv_std_logic_vector(27, 8),
44329 => conv_std_logic_vector(27, 8),
44330 => conv_std_logic_vector(28, 8),
44331 => conv_std_logic_vector(29, 8),
44332 => conv_std_logic_vector(29, 8),
44333 => conv_std_logic_vector(30, 8),
44334 => conv_std_logic_vector(31, 8),
44335 => conv_std_logic_vector(31, 8),
44336 => conv_std_logic_vector(32, 8),
44337 => conv_std_logic_vector(33, 8),
44338 => conv_std_logic_vector(33, 8),
44339 => conv_std_logic_vector(34, 8),
44340 => conv_std_logic_vector(35, 8),
44341 => conv_std_logic_vector(35, 8),
44342 => conv_std_logic_vector(36, 8),
44343 => conv_std_logic_vector(37, 8),
44344 => conv_std_logic_vector(37, 8),
44345 => conv_std_logic_vector(38, 8),
44346 => conv_std_logic_vector(39, 8),
44347 => conv_std_logic_vector(39, 8),
44348 => conv_std_logic_vector(40, 8),
44349 => conv_std_logic_vector(41, 8),
44350 => conv_std_logic_vector(41, 8),
44351 => conv_std_logic_vector(42, 8),
44352 => conv_std_logic_vector(43, 8),
44353 => conv_std_logic_vector(43, 8),
44354 => conv_std_logic_vector(44, 8),
44355 => conv_std_logic_vector(45, 8),
44356 => conv_std_logic_vector(45, 8),
44357 => conv_std_logic_vector(46, 8),
44358 => conv_std_logic_vector(47, 8),
44359 => conv_std_logic_vector(47, 8),
44360 => conv_std_logic_vector(48, 8),
44361 => conv_std_logic_vector(49, 8),
44362 => conv_std_logic_vector(50, 8),
44363 => conv_std_logic_vector(50, 8),
44364 => conv_std_logic_vector(51, 8),
44365 => conv_std_logic_vector(52, 8),
44366 => conv_std_logic_vector(52, 8),
44367 => conv_std_logic_vector(53, 8),
44368 => conv_std_logic_vector(54, 8),
44369 => conv_std_logic_vector(54, 8),
44370 => conv_std_logic_vector(55, 8),
44371 => conv_std_logic_vector(56, 8),
44372 => conv_std_logic_vector(56, 8),
44373 => conv_std_logic_vector(57, 8),
44374 => conv_std_logic_vector(58, 8),
44375 => conv_std_logic_vector(58, 8),
44376 => conv_std_logic_vector(59, 8),
44377 => conv_std_logic_vector(60, 8),
44378 => conv_std_logic_vector(60, 8),
44379 => conv_std_logic_vector(61, 8),
44380 => conv_std_logic_vector(62, 8),
44381 => conv_std_logic_vector(62, 8),
44382 => conv_std_logic_vector(63, 8),
44383 => conv_std_logic_vector(64, 8),
44384 => conv_std_logic_vector(64, 8),
44385 => conv_std_logic_vector(65, 8),
44386 => conv_std_logic_vector(66, 8),
44387 => conv_std_logic_vector(66, 8),
44388 => conv_std_logic_vector(67, 8),
44389 => conv_std_logic_vector(68, 8),
44390 => conv_std_logic_vector(68, 8),
44391 => conv_std_logic_vector(69, 8),
44392 => conv_std_logic_vector(70, 8),
44393 => conv_std_logic_vector(70, 8),
44394 => conv_std_logic_vector(71, 8),
44395 => conv_std_logic_vector(72, 8),
44396 => conv_std_logic_vector(72, 8),
44397 => conv_std_logic_vector(73, 8),
44398 => conv_std_logic_vector(74, 8),
44399 => conv_std_logic_vector(75, 8),
44400 => conv_std_logic_vector(75, 8),
44401 => conv_std_logic_vector(76, 8),
44402 => conv_std_logic_vector(77, 8),
44403 => conv_std_logic_vector(77, 8),
44404 => conv_std_logic_vector(78, 8),
44405 => conv_std_logic_vector(79, 8),
44406 => conv_std_logic_vector(79, 8),
44407 => conv_std_logic_vector(80, 8),
44408 => conv_std_logic_vector(81, 8),
44409 => conv_std_logic_vector(81, 8),
44410 => conv_std_logic_vector(82, 8),
44411 => conv_std_logic_vector(83, 8),
44412 => conv_std_logic_vector(83, 8),
44413 => conv_std_logic_vector(84, 8),
44414 => conv_std_logic_vector(85, 8),
44415 => conv_std_logic_vector(85, 8),
44416 => conv_std_logic_vector(86, 8),
44417 => conv_std_logic_vector(87, 8),
44418 => conv_std_logic_vector(87, 8),
44419 => conv_std_logic_vector(88, 8),
44420 => conv_std_logic_vector(89, 8),
44421 => conv_std_logic_vector(89, 8),
44422 => conv_std_logic_vector(90, 8),
44423 => conv_std_logic_vector(91, 8),
44424 => conv_std_logic_vector(91, 8),
44425 => conv_std_logic_vector(92, 8),
44426 => conv_std_logic_vector(93, 8),
44427 => conv_std_logic_vector(93, 8),
44428 => conv_std_logic_vector(94, 8),
44429 => conv_std_logic_vector(95, 8),
44430 => conv_std_logic_vector(95, 8),
44431 => conv_std_logic_vector(96, 8),
44432 => conv_std_logic_vector(97, 8),
44433 => conv_std_logic_vector(97, 8),
44434 => conv_std_logic_vector(98, 8),
44435 => conv_std_logic_vector(99, 8),
44436 => conv_std_logic_vector(100, 8),
44437 => conv_std_logic_vector(100, 8),
44438 => conv_std_logic_vector(101, 8),
44439 => conv_std_logic_vector(102, 8),
44440 => conv_std_logic_vector(102, 8),
44441 => conv_std_logic_vector(103, 8),
44442 => conv_std_logic_vector(104, 8),
44443 => conv_std_logic_vector(104, 8),
44444 => conv_std_logic_vector(105, 8),
44445 => conv_std_logic_vector(106, 8),
44446 => conv_std_logic_vector(106, 8),
44447 => conv_std_logic_vector(107, 8),
44448 => conv_std_logic_vector(108, 8),
44449 => conv_std_logic_vector(108, 8),
44450 => conv_std_logic_vector(109, 8),
44451 => conv_std_logic_vector(110, 8),
44452 => conv_std_logic_vector(110, 8),
44453 => conv_std_logic_vector(111, 8),
44454 => conv_std_logic_vector(112, 8),
44455 => conv_std_logic_vector(112, 8),
44456 => conv_std_logic_vector(113, 8),
44457 => conv_std_logic_vector(114, 8),
44458 => conv_std_logic_vector(114, 8),
44459 => conv_std_logic_vector(115, 8),
44460 => conv_std_logic_vector(116, 8),
44461 => conv_std_logic_vector(116, 8),
44462 => conv_std_logic_vector(117, 8),
44463 => conv_std_logic_vector(118, 8),
44464 => conv_std_logic_vector(118, 8),
44465 => conv_std_logic_vector(119, 8),
44466 => conv_std_logic_vector(120, 8),
44467 => conv_std_logic_vector(120, 8),
44468 => conv_std_logic_vector(121, 8),
44469 => conv_std_logic_vector(122, 8),
44470 => conv_std_logic_vector(122, 8),
44471 => conv_std_logic_vector(123, 8),
44472 => conv_std_logic_vector(124, 8),
44473 => conv_std_logic_vector(125, 8),
44474 => conv_std_logic_vector(125, 8),
44475 => conv_std_logic_vector(126, 8),
44476 => conv_std_logic_vector(127, 8),
44477 => conv_std_logic_vector(127, 8),
44478 => conv_std_logic_vector(128, 8),
44479 => conv_std_logic_vector(129, 8),
44480 => conv_std_logic_vector(129, 8),
44481 => conv_std_logic_vector(130, 8),
44482 => conv_std_logic_vector(131, 8),
44483 => conv_std_logic_vector(131, 8),
44484 => conv_std_logic_vector(132, 8),
44485 => conv_std_logic_vector(133, 8),
44486 => conv_std_logic_vector(133, 8),
44487 => conv_std_logic_vector(134, 8),
44488 => conv_std_logic_vector(135, 8),
44489 => conv_std_logic_vector(135, 8),
44490 => conv_std_logic_vector(136, 8),
44491 => conv_std_logic_vector(137, 8),
44492 => conv_std_logic_vector(137, 8),
44493 => conv_std_logic_vector(138, 8),
44494 => conv_std_logic_vector(139, 8),
44495 => conv_std_logic_vector(139, 8),
44496 => conv_std_logic_vector(140, 8),
44497 => conv_std_logic_vector(141, 8),
44498 => conv_std_logic_vector(141, 8),
44499 => conv_std_logic_vector(142, 8),
44500 => conv_std_logic_vector(143, 8),
44501 => conv_std_logic_vector(143, 8),
44502 => conv_std_logic_vector(144, 8),
44503 => conv_std_logic_vector(145, 8),
44504 => conv_std_logic_vector(145, 8),
44505 => conv_std_logic_vector(146, 8),
44506 => conv_std_logic_vector(147, 8),
44507 => conv_std_logic_vector(147, 8),
44508 => conv_std_logic_vector(148, 8),
44509 => conv_std_logic_vector(149, 8),
44510 => conv_std_logic_vector(150, 8),
44511 => conv_std_logic_vector(150, 8),
44512 => conv_std_logic_vector(151, 8),
44513 => conv_std_logic_vector(152, 8),
44514 => conv_std_logic_vector(152, 8),
44515 => conv_std_logic_vector(153, 8),
44516 => conv_std_logic_vector(154, 8),
44517 => conv_std_logic_vector(154, 8),
44518 => conv_std_logic_vector(155, 8),
44519 => conv_std_logic_vector(156, 8),
44520 => conv_std_logic_vector(156, 8),
44521 => conv_std_logic_vector(157, 8),
44522 => conv_std_logic_vector(158, 8),
44523 => conv_std_logic_vector(158, 8),
44524 => conv_std_logic_vector(159, 8),
44525 => conv_std_logic_vector(160, 8),
44526 => conv_std_logic_vector(160, 8),
44527 => conv_std_logic_vector(161, 8),
44528 => conv_std_logic_vector(162, 8),
44529 => conv_std_logic_vector(162, 8),
44530 => conv_std_logic_vector(163, 8),
44531 => conv_std_logic_vector(164, 8),
44532 => conv_std_logic_vector(164, 8),
44533 => conv_std_logic_vector(165, 8),
44534 => conv_std_logic_vector(166, 8),
44535 => conv_std_logic_vector(166, 8),
44536 => conv_std_logic_vector(167, 8),
44537 => conv_std_logic_vector(168, 8),
44538 => conv_std_logic_vector(168, 8),
44539 => conv_std_logic_vector(169, 8),
44540 => conv_std_logic_vector(170, 8),
44541 => conv_std_logic_vector(170, 8),
44542 => conv_std_logic_vector(171, 8),
44543 => conv_std_logic_vector(172, 8),
44544 => conv_std_logic_vector(0, 8),
44545 => conv_std_logic_vector(0, 8),
44546 => conv_std_logic_vector(1, 8),
44547 => conv_std_logic_vector(2, 8),
44548 => conv_std_logic_vector(2, 8),
44549 => conv_std_logic_vector(3, 8),
44550 => conv_std_logic_vector(4, 8),
44551 => conv_std_logic_vector(4, 8),
44552 => conv_std_logic_vector(5, 8),
44553 => conv_std_logic_vector(6, 8),
44554 => conv_std_logic_vector(6, 8),
44555 => conv_std_logic_vector(7, 8),
44556 => conv_std_logic_vector(8, 8),
44557 => conv_std_logic_vector(8, 8),
44558 => conv_std_logic_vector(9, 8),
44559 => conv_std_logic_vector(10, 8),
44560 => conv_std_logic_vector(10, 8),
44561 => conv_std_logic_vector(11, 8),
44562 => conv_std_logic_vector(12, 8),
44563 => conv_std_logic_vector(12, 8),
44564 => conv_std_logic_vector(13, 8),
44565 => conv_std_logic_vector(14, 8),
44566 => conv_std_logic_vector(14, 8),
44567 => conv_std_logic_vector(15, 8),
44568 => conv_std_logic_vector(16, 8),
44569 => conv_std_logic_vector(16, 8),
44570 => conv_std_logic_vector(17, 8),
44571 => conv_std_logic_vector(18, 8),
44572 => conv_std_logic_vector(19, 8),
44573 => conv_std_logic_vector(19, 8),
44574 => conv_std_logic_vector(20, 8),
44575 => conv_std_logic_vector(21, 8),
44576 => conv_std_logic_vector(21, 8),
44577 => conv_std_logic_vector(22, 8),
44578 => conv_std_logic_vector(23, 8),
44579 => conv_std_logic_vector(23, 8),
44580 => conv_std_logic_vector(24, 8),
44581 => conv_std_logic_vector(25, 8),
44582 => conv_std_logic_vector(25, 8),
44583 => conv_std_logic_vector(26, 8),
44584 => conv_std_logic_vector(27, 8),
44585 => conv_std_logic_vector(27, 8),
44586 => conv_std_logic_vector(28, 8),
44587 => conv_std_logic_vector(29, 8),
44588 => conv_std_logic_vector(29, 8),
44589 => conv_std_logic_vector(30, 8),
44590 => conv_std_logic_vector(31, 8),
44591 => conv_std_logic_vector(31, 8),
44592 => conv_std_logic_vector(32, 8),
44593 => conv_std_logic_vector(33, 8),
44594 => conv_std_logic_vector(33, 8),
44595 => conv_std_logic_vector(34, 8),
44596 => conv_std_logic_vector(35, 8),
44597 => conv_std_logic_vector(36, 8),
44598 => conv_std_logic_vector(36, 8),
44599 => conv_std_logic_vector(37, 8),
44600 => conv_std_logic_vector(38, 8),
44601 => conv_std_logic_vector(38, 8),
44602 => conv_std_logic_vector(39, 8),
44603 => conv_std_logic_vector(40, 8),
44604 => conv_std_logic_vector(40, 8),
44605 => conv_std_logic_vector(41, 8),
44606 => conv_std_logic_vector(42, 8),
44607 => conv_std_logic_vector(42, 8),
44608 => conv_std_logic_vector(43, 8),
44609 => conv_std_logic_vector(44, 8),
44610 => conv_std_logic_vector(44, 8),
44611 => conv_std_logic_vector(45, 8),
44612 => conv_std_logic_vector(46, 8),
44613 => conv_std_logic_vector(46, 8),
44614 => conv_std_logic_vector(47, 8),
44615 => conv_std_logic_vector(48, 8),
44616 => conv_std_logic_vector(48, 8),
44617 => conv_std_logic_vector(49, 8),
44618 => conv_std_logic_vector(50, 8),
44619 => conv_std_logic_vector(50, 8),
44620 => conv_std_logic_vector(51, 8),
44621 => conv_std_logic_vector(52, 8),
44622 => conv_std_logic_vector(53, 8),
44623 => conv_std_logic_vector(53, 8),
44624 => conv_std_logic_vector(54, 8),
44625 => conv_std_logic_vector(55, 8),
44626 => conv_std_logic_vector(55, 8),
44627 => conv_std_logic_vector(56, 8),
44628 => conv_std_logic_vector(57, 8),
44629 => conv_std_logic_vector(57, 8),
44630 => conv_std_logic_vector(58, 8),
44631 => conv_std_logic_vector(59, 8),
44632 => conv_std_logic_vector(59, 8),
44633 => conv_std_logic_vector(60, 8),
44634 => conv_std_logic_vector(61, 8),
44635 => conv_std_logic_vector(61, 8),
44636 => conv_std_logic_vector(62, 8),
44637 => conv_std_logic_vector(63, 8),
44638 => conv_std_logic_vector(63, 8),
44639 => conv_std_logic_vector(64, 8),
44640 => conv_std_logic_vector(65, 8),
44641 => conv_std_logic_vector(65, 8),
44642 => conv_std_logic_vector(66, 8),
44643 => conv_std_logic_vector(67, 8),
44644 => conv_std_logic_vector(67, 8),
44645 => conv_std_logic_vector(68, 8),
44646 => conv_std_logic_vector(69, 8),
44647 => conv_std_logic_vector(70, 8),
44648 => conv_std_logic_vector(70, 8),
44649 => conv_std_logic_vector(71, 8),
44650 => conv_std_logic_vector(72, 8),
44651 => conv_std_logic_vector(72, 8),
44652 => conv_std_logic_vector(73, 8),
44653 => conv_std_logic_vector(74, 8),
44654 => conv_std_logic_vector(74, 8),
44655 => conv_std_logic_vector(75, 8),
44656 => conv_std_logic_vector(76, 8),
44657 => conv_std_logic_vector(76, 8),
44658 => conv_std_logic_vector(77, 8),
44659 => conv_std_logic_vector(78, 8),
44660 => conv_std_logic_vector(78, 8),
44661 => conv_std_logic_vector(79, 8),
44662 => conv_std_logic_vector(80, 8),
44663 => conv_std_logic_vector(80, 8),
44664 => conv_std_logic_vector(81, 8),
44665 => conv_std_logic_vector(82, 8),
44666 => conv_std_logic_vector(82, 8),
44667 => conv_std_logic_vector(83, 8),
44668 => conv_std_logic_vector(84, 8),
44669 => conv_std_logic_vector(84, 8),
44670 => conv_std_logic_vector(85, 8),
44671 => conv_std_logic_vector(86, 8),
44672 => conv_std_logic_vector(87, 8),
44673 => conv_std_logic_vector(87, 8),
44674 => conv_std_logic_vector(88, 8),
44675 => conv_std_logic_vector(89, 8),
44676 => conv_std_logic_vector(89, 8),
44677 => conv_std_logic_vector(90, 8),
44678 => conv_std_logic_vector(91, 8),
44679 => conv_std_logic_vector(91, 8),
44680 => conv_std_logic_vector(92, 8),
44681 => conv_std_logic_vector(93, 8),
44682 => conv_std_logic_vector(93, 8),
44683 => conv_std_logic_vector(94, 8),
44684 => conv_std_logic_vector(95, 8),
44685 => conv_std_logic_vector(95, 8),
44686 => conv_std_logic_vector(96, 8),
44687 => conv_std_logic_vector(97, 8),
44688 => conv_std_logic_vector(97, 8),
44689 => conv_std_logic_vector(98, 8),
44690 => conv_std_logic_vector(99, 8),
44691 => conv_std_logic_vector(99, 8),
44692 => conv_std_logic_vector(100, 8),
44693 => conv_std_logic_vector(101, 8),
44694 => conv_std_logic_vector(101, 8),
44695 => conv_std_logic_vector(102, 8),
44696 => conv_std_logic_vector(103, 8),
44697 => conv_std_logic_vector(103, 8),
44698 => conv_std_logic_vector(104, 8),
44699 => conv_std_logic_vector(105, 8),
44700 => conv_std_logic_vector(106, 8),
44701 => conv_std_logic_vector(106, 8),
44702 => conv_std_logic_vector(107, 8),
44703 => conv_std_logic_vector(108, 8),
44704 => conv_std_logic_vector(108, 8),
44705 => conv_std_logic_vector(109, 8),
44706 => conv_std_logic_vector(110, 8),
44707 => conv_std_logic_vector(110, 8),
44708 => conv_std_logic_vector(111, 8),
44709 => conv_std_logic_vector(112, 8),
44710 => conv_std_logic_vector(112, 8),
44711 => conv_std_logic_vector(113, 8),
44712 => conv_std_logic_vector(114, 8),
44713 => conv_std_logic_vector(114, 8),
44714 => conv_std_logic_vector(115, 8),
44715 => conv_std_logic_vector(116, 8),
44716 => conv_std_logic_vector(116, 8),
44717 => conv_std_logic_vector(117, 8),
44718 => conv_std_logic_vector(118, 8),
44719 => conv_std_logic_vector(118, 8),
44720 => conv_std_logic_vector(119, 8),
44721 => conv_std_logic_vector(120, 8),
44722 => conv_std_logic_vector(120, 8),
44723 => conv_std_logic_vector(121, 8),
44724 => conv_std_logic_vector(122, 8),
44725 => conv_std_logic_vector(123, 8),
44726 => conv_std_logic_vector(123, 8),
44727 => conv_std_logic_vector(124, 8),
44728 => conv_std_logic_vector(125, 8),
44729 => conv_std_logic_vector(125, 8),
44730 => conv_std_logic_vector(126, 8),
44731 => conv_std_logic_vector(127, 8),
44732 => conv_std_logic_vector(127, 8),
44733 => conv_std_logic_vector(128, 8),
44734 => conv_std_logic_vector(129, 8),
44735 => conv_std_logic_vector(129, 8),
44736 => conv_std_logic_vector(130, 8),
44737 => conv_std_logic_vector(131, 8),
44738 => conv_std_logic_vector(131, 8),
44739 => conv_std_logic_vector(132, 8),
44740 => conv_std_logic_vector(133, 8),
44741 => conv_std_logic_vector(133, 8),
44742 => conv_std_logic_vector(134, 8),
44743 => conv_std_logic_vector(135, 8),
44744 => conv_std_logic_vector(135, 8),
44745 => conv_std_logic_vector(136, 8),
44746 => conv_std_logic_vector(137, 8),
44747 => conv_std_logic_vector(137, 8),
44748 => conv_std_logic_vector(138, 8),
44749 => conv_std_logic_vector(139, 8),
44750 => conv_std_logic_vector(140, 8),
44751 => conv_std_logic_vector(140, 8),
44752 => conv_std_logic_vector(141, 8),
44753 => conv_std_logic_vector(142, 8),
44754 => conv_std_logic_vector(142, 8),
44755 => conv_std_logic_vector(143, 8),
44756 => conv_std_logic_vector(144, 8),
44757 => conv_std_logic_vector(144, 8),
44758 => conv_std_logic_vector(145, 8),
44759 => conv_std_logic_vector(146, 8),
44760 => conv_std_logic_vector(146, 8),
44761 => conv_std_logic_vector(147, 8),
44762 => conv_std_logic_vector(148, 8),
44763 => conv_std_logic_vector(148, 8),
44764 => conv_std_logic_vector(149, 8),
44765 => conv_std_logic_vector(150, 8),
44766 => conv_std_logic_vector(150, 8),
44767 => conv_std_logic_vector(151, 8),
44768 => conv_std_logic_vector(152, 8),
44769 => conv_std_logic_vector(152, 8),
44770 => conv_std_logic_vector(153, 8),
44771 => conv_std_logic_vector(154, 8),
44772 => conv_std_logic_vector(154, 8),
44773 => conv_std_logic_vector(155, 8),
44774 => conv_std_logic_vector(156, 8),
44775 => conv_std_logic_vector(157, 8),
44776 => conv_std_logic_vector(157, 8),
44777 => conv_std_logic_vector(158, 8),
44778 => conv_std_logic_vector(159, 8),
44779 => conv_std_logic_vector(159, 8),
44780 => conv_std_logic_vector(160, 8),
44781 => conv_std_logic_vector(161, 8),
44782 => conv_std_logic_vector(161, 8),
44783 => conv_std_logic_vector(162, 8),
44784 => conv_std_logic_vector(163, 8),
44785 => conv_std_logic_vector(163, 8),
44786 => conv_std_logic_vector(164, 8),
44787 => conv_std_logic_vector(165, 8),
44788 => conv_std_logic_vector(165, 8),
44789 => conv_std_logic_vector(166, 8),
44790 => conv_std_logic_vector(167, 8),
44791 => conv_std_logic_vector(167, 8),
44792 => conv_std_logic_vector(168, 8),
44793 => conv_std_logic_vector(169, 8),
44794 => conv_std_logic_vector(169, 8),
44795 => conv_std_logic_vector(170, 8),
44796 => conv_std_logic_vector(171, 8),
44797 => conv_std_logic_vector(171, 8),
44798 => conv_std_logic_vector(172, 8),
44799 => conv_std_logic_vector(173, 8),
44800 => conv_std_logic_vector(0, 8),
44801 => conv_std_logic_vector(0, 8),
44802 => conv_std_logic_vector(1, 8),
44803 => conv_std_logic_vector(2, 8),
44804 => conv_std_logic_vector(2, 8),
44805 => conv_std_logic_vector(3, 8),
44806 => conv_std_logic_vector(4, 8),
44807 => conv_std_logic_vector(4, 8),
44808 => conv_std_logic_vector(5, 8),
44809 => conv_std_logic_vector(6, 8),
44810 => conv_std_logic_vector(6, 8),
44811 => conv_std_logic_vector(7, 8),
44812 => conv_std_logic_vector(8, 8),
44813 => conv_std_logic_vector(8, 8),
44814 => conv_std_logic_vector(9, 8),
44815 => conv_std_logic_vector(10, 8),
44816 => conv_std_logic_vector(10, 8),
44817 => conv_std_logic_vector(11, 8),
44818 => conv_std_logic_vector(12, 8),
44819 => conv_std_logic_vector(12, 8),
44820 => conv_std_logic_vector(13, 8),
44821 => conv_std_logic_vector(14, 8),
44822 => conv_std_logic_vector(15, 8),
44823 => conv_std_logic_vector(15, 8),
44824 => conv_std_logic_vector(16, 8),
44825 => conv_std_logic_vector(17, 8),
44826 => conv_std_logic_vector(17, 8),
44827 => conv_std_logic_vector(18, 8),
44828 => conv_std_logic_vector(19, 8),
44829 => conv_std_logic_vector(19, 8),
44830 => conv_std_logic_vector(20, 8),
44831 => conv_std_logic_vector(21, 8),
44832 => conv_std_logic_vector(21, 8),
44833 => conv_std_logic_vector(22, 8),
44834 => conv_std_logic_vector(23, 8),
44835 => conv_std_logic_vector(23, 8),
44836 => conv_std_logic_vector(24, 8),
44837 => conv_std_logic_vector(25, 8),
44838 => conv_std_logic_vector(25, 8),
44839 => conv_std_logic_vector(26, 8),
44840 => conv_std_logic_vector(27, 8),
44841 => conv_std_logic_vector(28, 8),
44842 => conv_std_logic_vector(28, 8),
44843 => conv_std_logic_vector(29, 8),
44844 => conv_std_logic_vector(30, 8),
44845 => conv_std_logic_vector(30, 8),
44846 => conv_std_logic_vector(31, 8),
44847 => conv_std_logic_vector(32, 8),
44848 => conv_std_logic_vector(32, 8),
44849 => conv_std_logic_vector(33, 8),
44850 => conv_std_logic_vector(34, 8),
44851 => conv_std_logic_vector(34, 8),
44852 => conv_std_logic_vector(35, 8),
44853 => conv_std_logic_vector(36, 8),
44854 => conv_std_logic_vector(36, 8),
44855 => conv_std_logic_vector(37, 8),
44856 => conv_std_logic_vector(38, 8),
44857 => conv_std_logic_vector(38, 8),
44858 => conv_std_logic_vector(39, 8),
44859 => conv_std_logic_vector(40, 8),
44860 => conv_std_logic_vector(41, 8),
44861 => conv_std_logic_vector(41, 8),
44862 => conv_std_logic_vector(42, 8),
44863 => conv_std_logic_vector(43, 8),
44864 => conv_std_logic_vector(43, 8),
44865 => conv_std_logic_vector(44, 8),
44866 => conv_std_logic_vector(45, 8),
44867 => conv_std_logic_vector(45, 8),
44868 => conv_std_logic_vector(46, 8),
44869 => conv_std_logic_vector(47, 8),
44870 => conv_std_logic_vector(47, 8),
44871 => conv_std_logic_vector(48, 8),
44872 => conv_std_logic_vector(49, 8),
44873 => conv_std_logic_vector(49, 8),
44874 => conv_std_logic_vector(50, 8),
44875 => conv_std_logic_vector(51, 8),
44876 => conv_std_logic_vector(51, 8),
44877 => conv_std_logic_vector(52, 8),
44878 => conv_std_logic_vector(53, 8),
44879 => conv_std_logic_vector(54, 8),
44880 => conv_std_logic_vector(54, 8),
44881 => conv_std_logic_vector(55, 8),
44882 => conv_std_logic_vector(56, 8),
44883 => conv_std_logic_vector(56, 8),
44884 => conv_std_logic_vector(57, 8),
44885 => conv_std_logic_vector(58, 8),
44886 => conv_std_logic_vector(58, 8),
44887 => conv_std_logic_vector(59, 8),
44888 => conv_std_logic_vector(60, 8),
44889 => conv_std_logic_vector(60, 8),
44890 => conv_std_logic_vector(61, 8),
44891 => conv_std_logic_vector(62, 8),
44892 => conv_std_logic_vector(62, 8),
44893 => conv_std_logic_vector(63, 8),
44894 => conv_std_logic_vector(64, 8),
44895 => conv_std_logic_vector(64, 8),
44896 => conv_std_logic_vector(65, 8),
44897 => conv_std_logic_vector(66, 8),
44898 => conv_std_logic_vector(66, 8),
44899 => conv_std_logic_vector(67, 8),
44900 => conv_std_logic_vector(68, 8),
44901 => conv_std_logic_vector(69, 8),
44902 => conv_std_logic_vector(69, 8),
44903 => conv_std_logic_vector(70, 8),
44904 => conv_std_logic_vector(71, 8),
44905 => conv_std_logic_vector(71, 8),
44906 => conv_std_logic_vector(72, 8),
44907 => conv_std_logic_vector(73, 8),
44908 => conv_std_logic_vector(73, 8),
44909 => conv_std_logic_vector(74, 8),
44910 => conv_std_logic_vector(75, 8),
44911 => conv_std_logic_vector(75, 8),
44912 => conv_std_logic_vector(76, 8),
44913 => conv_std_logic_vector(77, 8),
44914 => conv_std_logic_vector(77, 8),
44915 => conv_std_logic_vector(78, 8),
44916 => conv_std_logic_vector(79, 8),
44917 => conv_std_logic_vector(79, 8),
44918 => conv_std_logic_vector(80, 8),
44919 => conv_std_logic_vector(81, 8),
44920 => conv_std_logic_vector(82, 8),
44921 => conv_std_logic_vector(82, 8),
44922 => conv_std_logic_vector(83, 8),
44923 => conv_std_logic_vector(84, 8),
44924 => conv_std_logic_vector(84, 8),
44925 => conv_std_logic_vector(85, 8),
44926 => conv_std_logic_vector(86, 8),
44927 => conv_std_logic_vector(86, 8),
44928 => conv_std_logic_vector(87, 8),
44929 => conv_std_logic_vector(88, 8),
44930 => conv_std_logic_vector(88, 8),
44931 => conv_std_logic_vector(89, 8),
44932 => conv_std_logic_vector(90, 8),
44933 => conv_std_logic_vector(90, 8),
44934 => conv_std_logic_vector(91, 8),
44935 => conv_std_logic_vector(92, 8),
44936 => conv_std_logic_vector(92, 8),
44937 => conv_std_logic_vector(93, 8),
44938 => conv_std_logic_vector(94, 8),
44939 => conv_std_logic_vector(95, 8),
44940 => conv_std_logic_vector(95, 8),
44941 => conv_std_logic_vector(96, 8),
44942 => conv_std_logic_vector(97, 8),
44943 => conv_std_logic_vector(97, 8),
44944 => conv_std_logic_vector(98, 8),
44945 => conv_std_logic_vector(99, 8),
44946 => conv_std_logic_vector(99, 8),
44947 => conv_std_logic_vector(100, 8),
44948 => conv_std_logic_vector(101, 8),
44949 => conv_std_logic_vector(101, 8),
44950 => conv_std_logic_vector(102, 8),
44951 => conv_std_logic_vector(103, 8),
44952 => conv_std_logic_vector(103, 8),
44953 => conv_std_logic_vector(104, 8),
44954 => conv_std_logic_vector(105, 8),
44955 => conv_std_logic_vector(105, 8),
44956 => conv_std_logic_vector(106, 8),
44957 => conv_std_logic_vector(107, 8),
44958 => conv_std_logic_vector(108, 8),
44959 => conv_std_logic_vector(108, 8),
44960 => conv_std_logic_vector(109, 8),
44961 => conv_std_logic_vector(110, 8),
44962 => conv_std_logic_vector(110, 8),
44963 => conv_std_logic_vector(111, 8),
44964 => conv_std_logic_vector(112, 8),
44965 => conv_std_logic_vector(112, 8),
44966 => conv_std_logic_vector(113, 8),
44967 => conv_std_logic_vector(114, 8),
44968 => conv_std_logic_vector(114, 8),
44969 => conv_std_logic_vector(115, 8),
44970 => conv_std_logic_vector(116, 8),
44971 => conv_std_logic_vector(116, 8),
44972 => conv_std_logic_vector(117, 8),
44973 => conv_std_logic_vector(118, 8),
44974 => conv_std_logic_vector(118, 8),
44975 => conv_std_logic_vector(119, 8),
44976 => conv_std_logic_vector(120, 8),
44977 => conv_std_logic_vector(120, 8),
44978 => conv_std_logic_vector(121, 8),
44979 => conv_std_logic_vector(122, 8),
44980 => conv_std_logic_vector(123, 8),
44981 => conv_std_logic_vector(123, 8),
44982 => conv_std_logic_vector(124, 8),
44983 => conv_std_logic_vector(125, 8),
44984 => conv_std_logic_vector(125, 8),
44985 => conv_std_logic_vector(126, 8),
44986 => conv_std_logic_vector(127, 8),
44987 => conv_std_logic_vector(127, 8),
44988 => conv_std_logic_vector(128, 8),
44989 => conv_std_logic_vector(129, 8),
44990 => conv_std_logic_vector(129, 8),
44991 => conv_std_logic_vector(130, 8),
44992 => conv_std_logic_vector(131, 8),
44993 => conv_std_logic_vector(131, 8),
44994 => conv_std_logic_vector(132, 8),
44995 => conv_std_logic_vector(133, 8),
44996 => conv_std_logic_vector(133, 8),
44997 => conv_std_logic_vector(134, 8),
44998 => conv_std_logic_vector(135, 8),
44999 => conv_std_logic_vector(136, 8),
45000 => conv_std_logic_vector(136, 8),
45001 => conv_std_logic_vector(137, 8),
45002 => conv_std_logic_vector(138, 8),
45003 => conv_std_logic_vector(138, 8),
45004 => conv_std_logic_vector(139, 8),
45005 => conv_std_logic_vector(140, 8),
45006 => conv_std_logic_vector(140, 8),
45007 => conv_std_logic_vector(141, 8),
45008 => conv_std_logic_vector(142, 8),
45009 => conv_std_logic_vector(142, 8),
45010 => conv_std_logic_vector(143, 8),
45011 => conv_std_logic_vector(144, 8),
45012 => conv_std_logic_vector(144, 8),
45013 => conv_std_logic_vector(145, 8),
45014 => conv_std_logic_vector(146, 8),
45015 => conv_std_logic_vector(146, 8),
45016 => conv_std_logic_vector(147, 8),
45017 => conv_std_logic_vector(148, 8),
45018 => conv_std_logic_vector(149, 8),
45019 => conv_std_logic_vector(149, 8),
45020 => conv_std_logic_vector(150, 8),
45021 => conv_std_logic_vector(151, 8),
45022 => conv_std_logic_vector(151, 8),
45023 => conv_std_logic_vector(152, 8),
45024 => conv_std_logic_vector(153, 8),
45025 => conv_std_logic_vector(153, 8),
45026 => conv_std_logic_vector(154, 8),
45027 => conv_std_logic_vector(155, 8),
45028 => conv_std_logic_vector(155, 8),
45029 => conv_std_logic_vector(156, 8),
45030 => conv_std_logic_vector(157, 8),
45031 => conv_std_logic_vector(157, 8),
45032 => conv_std_logic_vector(158, 8),
45033 => conv_std_logic_vector(159, 8),
45034 => conv_std_logic_vector(159, 8),
45035 => conv_std_logic_vector(160, 8),
45036 => conv_std_logic_vector(161, 8),
45037 => conv_std_logic_vector(162, 8),
45038 => conv_std_logic_vector(162, 8),
45039 => conv_std_logic_vector(163, 8),
45040 => conv_std_logic_vector(164, 8),
45041 => conv_std_logic_vector(164, 8),
45042 => conv_std_logic_vector(165, 8),
45043 => conv_std_logic_vector(166, 8),
45044 => conv_std_logic_vector(166, 8),
45045 => conv_std_logic_vector(167, 8),
45046 => conv_std_logic_vector(168, 8),
45047 => conv_std_logic_vector(168, 8),
45048 => conv_std_logic_vector(169, 8),
45049 => conv_std_logic_vector(170, 8),
45050 => conv_std_logic_vector(170, 8),
45051 => conv_std_logic_vector(171, 8),
45052 => conv_std_logic_vector(172, 8),
45053 => conv_std_logic_vector(172, 8),
45054 => conv_std_logic_vector(173, 8),
45055 => conv_std_logic_vector(174, 8),
45056 => conv_std_logic_vector(0, 8),
45057 => conv_std_logic_vector(0, 8),
45058 => conv_std_logic_vector(1, 8),
45059 => conv_std_logic_vector(2, 8),
45060 => conv_std_logic_vector(2, 8),
45061 => conv_std_logic_vector(3, 8),
45062 => conv_std_logic_vector(4, 8),
45063 => conv_std_logic_vector(4, 8),
45064 => conv_std_logic_vector(5, 8),
45065 => conv_std_logic_vector(6, 8),
45066 => conv_std_logic_vector(6, 8),
45067 => conv_std_logic_vector(7, 8),
45068 => conv_std_logic_vector(8, 8),
45069 => conv_std_logic_vector(8, 8),
45070 => conv_std_logic_vector(9, 8),
45071 => conv_std_logic_vector(10, 8),
45072 => conv_std_logic_vector(11, 8),
45073 => conv_std_logic_vector(11, 8),
45074 => conv_std_logic_vector(12, 8),
45075 => conv_std_logic_vector(13, 8),
45076 => conv_std_logic_vector(13, 8),
45077 => conv_std_logic_vector(14, 8),
45078 => conv_std_logic_vector(15, 8),
45079 => conv_std_logic_vector(15, 8),
45080 => conv_std_logic_vector(16, 8),
45081 => conv_std_logic_vector(17, 8),
45082 => conv_std_logic_vector(17, 8),
45083 => conv_std_logic_vector(18, 8),
45084 => conv_std_logic_vector(19, 8),
45085 => conv_std_logic_vector(19, 8),
45086 => conv_std_logic_vector(20, 8),
45087 => conv_std_logic_vector(21, 8),
45088 => conv_std_logic_vector(22, 8),
45089 => conv_std_logic_vector(22, 8),
45090 => conv_std_logic_vector(23, 8),
45091 => conv_std_logic_vector(24, 8),
45092 => conv_std_logic_vector(24, 8),
45093 => conv_std_logic_vector(25, 8),
45094 => conv_std_logic_vector(26, 8),
45095 => conv_std_logic_vector(26, 8),
45096 => conv_std_logic_vector(27, 8),
45097 => conv_std_logic_vector(28, 8),
45098 => conv_std_logic_vector(28, 8),
45099 => conv_std_logic_vector(29, 8),
45100 => conv_std_logic_vector(30, 8),
45101 => conv_std_logic_vector(30, 8),
45102 => conv_std_logic_vector(31, 8),
45103 => conv_std_logic_vector(32, 8),
45104 => conv_std_logic_vector(33, 8),
45105 => conv_std_logic_vector(33, 8),
45106 => conv_std_logic_vector(34, 8),
45107 => conv_std_logic_vector(35, 8),
45108 => conv_std_logic_vector(35, 8),
45109 => conv_std_logic_vector(36, 8),
45110 => conv_std_logic_vector(37, 8),
45111 => conv_std_logic_vector(37, 8),
45112 => conv_std_logic_vector(38, 8),
45113 => conv_std_logic_vector(39, 8),
45114 => conv_std_logic_vector(39, 8),
45115 => conv_std_logic_vector(40, 8),
45116 => conv_std_logic_vector(41, 8),
45117 => conv_std_logic_vector(41, 8),
45118 => conv_std_logic_vector(42, 8),
45119 => conv_std_logic_vector(43, 8),
45120 => conv_std_logic_vector(44, 8),
45121 => conv_std_logic_vector(44, 8),
45122 => conv_std_logic_vector(45, 8),
45123 => conv_std_logic_vector(46, 8),
45124 => conv_std_logic_vector(46, 8),
45125 => conv_std_logic_vector(47, 8),
45126 => conv_std_logic_vector(48, 8),
45127 => conv_std_logic_vector(48, 8),
45128 => conv_std_logic_vector(49, 8),
45129 => conv_std_logic_vector(50, 8),
45130 => conv_std_logic_vector(50, 8),
45131 => conv_std_logic_vector(51, 8),
45132 => conv_std_logic_vector(52, 8),
45133 => conv_std_logic_vector(52, 8),
45134 => conv_std_logic_vector(53, 8),
45135 => conv_std_logic_vector(54, 8),
45136 => conv_std_logic_vector(55, 8),
45137 => conv_std_logic_vector(55, 8),
45138 => conv_std_logic_vector(56, 8),
45139 => conv_std_logic_vector(57, 8),
45140 => conv_std_logic_vector(57, 8),
45141 => conv_std_logic_vector(58, 8),
45142 => conv_std_logic_vector(59, 8),
45143 => conv_std_logic_vector(59, 8),
45144 => conv_std_logic_vector(60, 8),
45145 => conv_std_logic_vector(61, 8),
45146 => conv_std_logic_vector(61, 8),
45147 => conv_std_logic_vector(62, 8),
45148 => conv_std_logic_vector(63, 8),
45149 => conv_std_logic_vector(63, 8),
45150 => conv_std_logic_vector(64, 8),
45151 => conv_std_logic_vector(65, 8),
45152 => conv_std_logic_vector(66, 8),
45153 => conv_std_logic_vector(66, 8),
45154 => conv_std_logic_vector(67, 8),
45155 => conv_std_logic_vector(68, 8),
45156 => conv_std_logic_vector(68, 8),
45157 => conv_std_logic_vector(69, 8),
45158 => conv_std_logic_vector(70, 8),
45159 => conv_std_logic_vector(70, 8),
45160 => conv_std_logic_vector(71, 8),
45161 => conv_std_logic_vector(72, 8),
45162 => conv_std_logic_vector(72, 8),
45163 => conv_std_logic_vector(73, 8),
45164 => conv_std_logic_vector(74, 8),
45165 => conv_std_logic_vector(74, 8),
45166 => conv_std_logic_vector(75, 8),
45167 => conv_std_logic_vector(76, 8),
45168 => conv_std_logic_vector(77, 8),
45169 => conv_std_logic_vector(77, 8),
45170 => conv_std_logic_vector(78, 8),
45171 => conv_std_logic_vector(79, 8),
45172 => conv_std_logic_vector(79, 8),
45173 => conv_std_logic_vector(80, 8),
45174 => conv_std_logic_vector(81, 8),
45175 => conv_std_logic_vector(81, 8),
45176 => conv_std_logic_vector(82, 8),
45177 => conv_std_logic_vector(83, 8),
45178 => conv_std_logic_vector(83, 8),
45179 => conv_std_logic_vector(84, 8),
45180 => conv_std_logic_vector(85, 8),
45181 => conv_std_logic_vector(85, 8),
45182 => conv_std_logic_vector(86, 8),
45183 => conv_std_logic_vector(87, 8),
45184 => conv_std_logic_vector(88, 8),
45185 => conv_std_logic_vector(88, 8),
45186 => conv_std_logic_vector(89, 8),
45187 => conv_std_logic_vector(90, 8),
45188 => conv_std_logic_vector(90, 8),
45189 => conv_std_logic_vector(91, 8),
45190 => conv_std_logic_vector(92, 8),
45191 => conv_std_logic_vector(92, 8),
45192 => conv_std_logic_vector(93, 8),
45193 => conv_std_logic_vector(94, 8),
45194 => conv_std_logic_vector(94, 8),
45195 => conv_std_logic_vector(95, 8),
45196 => conv_std_logic_vector(96, 8),
45197 => conv_std_logic_vector(96, 8),
45198 => conv_std_logic_vector(97, 8),
45199 => conv_std_logic_vector(98, 8),
45200 => conv_std_logic_vector(99, 8),
45201 => conv_std_logic_vector(99, 8),
45202 => conv_std_logic_vector(100, 8),
45203 => conv_std_logic_vector(101, 8),
45204 => conv_std_logic_vector(101, 8),
45205 => conv_std_logic_vector(102, 8),
45206 => conv_std_logic_vector(103, 8),
45207 => conv_std_logic_vector(103, 8),
45208 => conv_std_logic_vector(104, 8),
45209 => conv_std_logic_vector(105, 8),
45210 => conv_std_logic_vector(105, 8),
45211 => conv_std_logic_vector(106, 8),
45212 => conv_std_logic_vector(107, 8),
45213 => conv_std_logic_vector(107, 8),
45214 => conv_std_logic_vector(108, 8),
45215 => conv_std_logic_vector(109, 8),
45216 => conv_std_logic_vector(110, 8),
45217 => conv_std_logic_vector(110, 8),
45218 => conv_std_logic_vector(111, 8),
45219 => conv_std_logic_vector(112, 8),
45220 => conv_std_logic_vector(112, 8),
45221 => conv_std_logic_vector(113, 8),
45222 => conv_std_logic_vector(114, 8),
45223 => conv_std_logic_vector(114, 8),
45224 => conv_std_logic_vector(115, 8),
45225 => conv_std_logic_vector(116, 8),
45226 => conv_std_logic_vector(116, 8),
45227 => conv_std_logic_vector(117, 8),
45228 => conv_std_logic_vector(118, 8),
45229 => conv_std_logic_vector(118, 8),
45230 => conv_std_logic_vector(119, 8),
45231 => conv_std_logic_vector(120, 8),
45232 => conv_std_logic_vector(121, 8),
45233 => conv_std_logic_vector(121, 8),
45234 => conv_std_logic_vector(122, 8),
45235 => conv_std_logic_vector(123, 8),
45236 => conv_std_logic_vector(123, 8),
45237 => conv_std_logic_vector(124, 8),
45238 => conv_std_logic_vector(125, 8),
45239 => conv_std_logic_vector(125, 8),
45240 => conv_std_logic_vector(126, 8),
45241 => conv_std_logic_vector(127, 8),
45242 => conv_std_logic_vector(127, 8),
45243 => conv_std_logic_vector(128, 8),
45244 => conv_std_logic_vector(129, 8),
45245 => conv_std_logic_vector(129, 8),
45246 => conv_std_logic_vector(130, 8),
45247 => conv_std_logic_vector(131, 8),
45248 => conv_std_logic_vector(132, 8),
45249 => conv_std_logic_vector(132, 8),
45250 => conv_std_logic_vector(133, 8),
45251 => conv_std_logic_vector(134, 8),
45252 => conv_std_logic_vector(134, 8),
45253 => conv_std_logic_vector(135, 8),
45254 => conv_std_logic_vector(136, 8),
45255 => conv_std_logic_vector(136, 8),
45256 => conv_std_logic_vector(137, 8),
45257 => conv_std_logic_vector(138, 8),
45258 => conv_std_logic_vector(138, 8),
45259 => conv_std_logic_vector(139, 8),
45260 => conv_std_logic_vector(140, 8),
45261 => conv_std_logic_vector(140, 8),
45262 => conv_std_logic_vector(141, 8),
45263 => conv_std_logic_vector(142, 8),
45264 => conv_std_logic_vector(143, 8),
45265 => conv_std_logic_vector(143, 8),
45266 => conv_std_logic_vector(144, 8),
45267 => conv_std_logic_vector(145, 8),
45268 => conv_std_logic_vector(145, 8),
45269 => conv_std_logic_vector(146, 8),
45270 => conv_std_logic_vector(147, 8),
45271 => conv_std_logic_vector(147, 8),
45272 => conv_std_logic_vector(148, 8),
45273 => conv_std_logic_vector(149, 8),
45274 => conv_std_logic_vector(149, 8),
45275 => conv_std_logic_vector(150, 8),
45276 => conv_std_logic_vector(151, 8),
45277 => conv_std_logic_vector(151, 8),
45278 => conv_std_logic_vector(152, 8),
45279 => conv_std_logic_vector(153, 8),
45280 => conv_std_logic_vector(154, 8),
45281 => conv_std_logic_vector(154, 8),
45282 => conv_std_logic_vector(155, 8),
45283 => conv_std_logic_vector(156, 8),
45284 => conv_std_logic_vector(156, 8),
45285 => conv_std_logic_vector(157, 8),
45286 => conv_std_logic_vector(158, 8),
45287 => conv_std_logic_vector(158, 8),
45288 => conv_std_logic_vector(159, 8),
45289 => conv_std_logic_vector(160, 8),
45290 => conv_std_logic_vector(160, 8),
45291 => conv_std_logic_vector(161, 8),
45292 => conv_std_logic_vector(162, 8),
45293 => conv_std_logic_vector(162, 8),
45294 => conv_std_logic_vector(163, 8),
45295 => conv_std_logic_vector(164, 8),
45296 => conv_std_logic_vector(165, 8),
45297 => conv_std_logic_vector(165, 8),
45298 => conv_std_logic_vector(166, 8),
45299 => conv_std_logic_vector(167, 8),
45300 => conv_std_logic_vector(167, 8),
45301 => conv_std_logic_vector(168, 8),
45302 => conv_std_logic_vector(169, 8),
45303 => conv_std_logic_vector(169, 8),
45304 => conv_std_logic_vector(170, 8),
45305 => conv_std_logic_vector(171, 8),
45306 => conv_std_logic_vector(171, 8),
45307 => conv_std_logic_vector(172, 8),
45308 => conv_std_logic_vector(173, 8),
45309 => conv_std_logic_vector(173, 8),
45310 => conv_std_logic_vector(174, 8),
45311 => conv_std_logic_vector(175, 8),
45312 => conv_std_logic_vector(0, 8),
45313 => conv_std_logic_vector(0, 8),
45314 => conv_std_logic_vector(1, 8),
45315 => conv_std_logic_vector(2, 8),
45316 => conv_std_logic_vector(2, 8),
45317 => conv_std_logic_vector(3, 8),
45318 => conv_std_logic_vector(4, 8),
45319 => conv_std_logic_vector(4, 8),
45320 => conv_std_logic_vector(5, 8),
45321 => conv_std_logic_vector(6, 8),
45322 => conv_std_logic_vector(6, 8),
45323 => conv_std_logic_vector(7, 8),
45324 => conv_std_logic_vector(8, 8),
45325 => conv_std_logic_vector(8, 8),
45326 => conv_std_logic_vector(9, 8),
45327 => conv_std_logic_vector(10, 8),
45328 => conv_std_logic_vector(11, 8),
45329 => conv_std_logic_vector(11, 8),
45330 => conv_std_logic_vector(12, 8),
45331 => conv_std_logic_vector(13, 8),
45332 => conv_std_logic_vector(13, 8),
45333 => conv_std_logic_vector(14, 8),
45334 => conv_std_logic_vector(15, 8),
45335 => conv_std_logic_vector(15, 8),
45336 => conv_std_logic_vector(16, 8),
45337 => conv_std_logic_vector(17, 8),
45338 => conv_std_logic_vector(17, 8),
45339 => conv_std_logic_vector(18, 8),
45340 => conv_std_logic_vector(19, 8),
45341 => conv_std_logic_vector(20, 8),
45342 => conv_std_logic_vector(20, 8),
45343 => conv_std_logic_vector(21, 8),
45344 => conv_std_logic_vector(22, 8),
45345 => conv_std_logic_vector(22, 8),
45346 => conv_std_logic_vector(23, 8),
45347 => conv_std_logic_vector(24, 8),
45348 => conv_std_logic_vector(24, 8),
45349 => conv_std_logic_vector(25, 8),
45350 => conv_std_logic_vector(26, 8),
45351 => conv_std_logic_vector(26, 8),
45352 => conv_std_logic_vector(27, 8),
45353 => conv_std_logic_vector(28, 8),
45354 => conv_std_logic_vector(29, 8),
45355 => conv_std_logic_vector(29, 8),
45356 => conv_std_logic_vector(30, 8),
45357 => conv_std_logic_vector(31, 8),
45358 => conv_std_logic_vector(31, 8),
45359 => conv_std_logic_vector(32, 8),
45360 => conv_std_logic_vector(33, 8),
45361 => conv_std_logic_vector(33, 8),
45362 => conv_std_logic_vector(34, 8),
45363 => conv_std_logic_vector(35, 8),
45364 => conv_std_logic_vector(35, 8),
45365 => conv_std_logic_vector(36, 8),
45366 => conv_std_logic_vector(37, 8),
45367 => conv_std_logic_vector(38, 8),
45368 => conv_std_logic_vector(38, 8),
45369 => conv_std_logic_vector(39, 8),
45370 => conv_std_logic_vector(40, 8),
45371 => conv_std_logic_vector(40, 8),
45372 => conv_std_logic_vector(41, 8),
45373 => conv_std_logic_vector(42, 8),
45374 => conv_std_logic_vector(42, 8),
45375 => conv_std_logic_vector(43, 8),
45376 => conv_std_logic_vector(44, 8),
45377 => conv_std_logic_vector(44, 8),
45378 => conv_std_logic_vector(45, 8),
45379 => conv_std_logic_vector(46, 8),
45380 => conv_std_logic_vector(47, 8),
45381 => conv_std_logic_vector(47, 8),
45382 => conv_std_logic_vector(48, 8),
45383 => conv_std_logic_vector(49, 8),
45384 => conv_std_logic_vector(49, 8),
45385 => conv_std_logic_vector(50, 8),
45386 => conv_std_logic_vector(51, 8),
45387 => conv_std_logic_vector(51, 8),
45388 => conv_std_logic_vector(52, 8),
45389 => conv_std_logic_vector(53, 8),
45390 => conv_std_logic_vector(53, 8),
45391 => conv_std_logic_vector(54, 8),
45392 => conv_std_logic_vector(55, 8),
45393 => conv_std_logic_vector(56, 8),
45394 => conv_std_logic_vector(56, 8),
45395 => conv_std_logic_vector(57, 8),
45396 => conv_std_logic_vector(58, 8),
45397 => conv_std_logic_vector(58, 8),
45398 => conv_std_logic_vector(59, 8),
45399 => conv_std_logic_vector(60, 8),
45400 => conv_std_logic_vector(60, 8),
45401 => conv_std_logic_vector(61, 8),
45402 => conv_std_logic_vector(62, 8),
45403 => conv_std_logic_vector(62, 8),
45404 => conv_std_logic_vector(63, 8),
45405 => conv_std_logic_vector(64, 8),
45406 => conv_std_logic_vector(64, 8),
45407 => conv_std_logic_vector(65, 8),
45408 => conv_std_logic_vector(66, 8),
45409 => conv_std_logic_vector(67, 8),
45410 => conv_std_logic_vector(67, 8),
45411 => conv_std_logic_vector(68, 8),
45412 => conv_std_logic_vector(69, 8),
45413 => conv_std_logic_vector(69, 8),
45414 => conv_std_logic_vector(70, 8),
45415 => conv_std_logic_vector(71, 8),
45416 => conv_std_logic_vector(71, 8),
45417 => conv_std_logic_vector(72, 8),
45418 => conv_std_logic_vector(73, 8),
45419 => conv_std_logic_vector(73, 8),
45420 => conv_std_logic_vector(74, 8),
45421 => conv_std_logic_vector(75, 8),
45422 => conv_std_logic_vector(76, 8),
45423 => conv_std_logic_vector(76, 8),
45424 => conv_std_logic_vector(77, 8),
45425 => conv_std_logic_vector(78, 8),
45426 => conv_std_logic_vector(78, 8),
45427 => conv_std_logic_vector(79, 8),
45428 => conv_std_logic_vector(80, 8),
45429 => conv_std_logic_vector(80, 8),
45430 => conv_std_logic_vector(81, 8),
45431 => conv_std_logic_vector(82, 8),
45432 => conv_std_logic_vector(82, 8),
45433 => conv_std_logic_vector(83, 8),
45434 => conv_std_logic_vector(84, 8),
45435 => conv_std_logic_vector(85, 8),
45436 => conv_std_logic_vector(85, 8),
45437 => conv_std_logic_vector(86, 8),
45438 => conv_std_logic_vector(87, 8),
45439 => conv_std_logic_vector(87, 8),
45440 => conv_std_logic_vector(88, 8),
45441 => conv_std_logic_vector(89, 8),
45442 => conv_std_logic_vector(89, 8),
45443 => conv_std_logic_vector(90, 8),
45444 => conv_std_logic_vector(91, 8),
45445 => conv_std_logic_vector(91, 8),
45446 => conv_std_logic_vector(92, 8),
45447 => conv_std_logic_vector(93, 8),
45448 => conv_std_logic_vector(94, 8),
45449 => conv_std_logic_vector(94, 8),
45450 => conv_std_logic_vector(95, 8),
45451 => conv_std_logic_vector(96, 8),
45452 => conv_std_logic_vector(96, 8),
45453 => conv_std_logic_vector(97, 8),
45454 => conv_std_logic_vector(98, 8),
45455 => conv_std_logic_vector(98, 8),
45456 => conv_std_logic_vector(99, 8),
45457 => conv_std_logic_vector(100, 8),
45458 => conv_std_logic_vector(100, 8),
45459 => conv_std_logic_vector(101, 8),
45460 => conv_std_logic_vector(102, 8),
45461 => conv_std_logic_vector(103, 8),
45462 => conv_std_logic_vector(103, 8),
45463 => conv_std_logic_vector(104, 8),
45464 => conv_std_logic_vector(105, 8),
45465 => conv_std_logic_vector(105, 8),
45466 => conv_std_logic_vector(106, 8),
45467 => conv_std_logic_vector(107, 8),
45468 => conv_std_logic_vector(107, 8),
45469 => conv_std_logic_vector(108, 8),
45470 => conv_std_logic_vector(109, 8),
45471 => conv_std_logic_vector(109, 8),
45472 => conv_std_logic_vector(110, 8),
45473 => conv_std_logic_vector(111, 8),
45474 => conv_std_logic_vector(112, 8),
45475 => conv_std_logic_vector(112, 8),
45476 => conv_std_logic_vector(113, 8),
45477 => conv_std_logic_vector(114, 8),
45478 => conv_std_logic_vector(114, 8),
45479 => conv_std_logic_vector(115, 8),
45480 => conv_std_logic_vector(116, 8),
45481 => conv_std_logic_vector(116, 8),
45482 => conv_std_logic_vector(117, 8),
45483 => conv_std_logic_vector(118, 8),
45484 => conv_std_logic_vector(118, 8),
45485 => conv_std_logic_vector(119, 8),
45486 => conv_std_logic_vector(120, 8),
45487 => conv_std_logic_vector(120, 8),
45488 => conv_std_logic_vector(121, 8),
45489 => conv_std_logic_vector(122, 8),
45490 => conv_std_logic_vector(123, 8),
45491 => conv_std_logic_vector(123, 8),
45492 => conv_std_logic_vector(124, 8),
45493 => conv_std_logic_vector(125, 8),
45494 => conv_std_logic_vector(125, 8),
45495 => conv_std_logic_vector(126, 8),
45496 => conv_std_logic_vector(127, 8),
45497 => conv_std_logic_vector(127, 8),
45498 => conv_std_logic_vector(128, 8),
45499 => conv_std_logic_vector(129, 8),
45500 => conv_std_logic_vector(129, 8),
45501 => conv_std_logic_vector(130, 8),
45502 => conv_std_logic_vector(131, 8),
45503 => conv_std_logic_vector(132, 8),
45504 => conv_std_logic_vector(132, 8),
45505 => conv_std_logic_vector(133, 8),
45506 => conv_std_logic_vector(134, 8),
45507 => conv_std_logic_vector(134, 8),
45508 => conv_std_logic_vector(135, 8),
45509 => conv_std_logic_vector(136, 8),
45510 => conv_std_logic_vector(136, 8),
45511 => conv_std_logic_vector(137, 8),
45512 => conv_std_logic_vector(138, 8),
45513 => conv_std_logic_vector(138, 8),
45514 => conv_std_logic_vector(139, 8),
45515 => conv_std_logic_vector(140, 8),
45516 => conv_std_logic_vector(141, 8),
45517 => conv_std_logic_vector(141, 8),
45518 => conv_std_logic_vector(142, 8),
45519 => conv_std_logic_vector(143, 8),
45520 => conv_std_logic_vector(143, 8),
45521 => conv_std_logic_vector(144, 8),
45522 => conv_std_logic_vector(145, 8),
45523 => conv_std_logic_vector(145, 8),
45524 => conv_std_logic_vector(146, 8),
45525 => conv_std_logic_vector(147, 8),
45526 => conv_std_logic_vector(147, 8),
45527 => conv_std_logic_vector(148, 8),
45528 => conv_std_logic_vector(149, 8),
45529 => conv_std_logic_vector(150, 8),
45530 => conv_std_logic_vector(150, 8),
45531 => conv_std_logic_vector(151, 8),
45532 => conv_std_logic_vector(152, 8),
45533 => conv_std_logic_vector(152, 8),
45534 => conv_std_logic_vector(153, 8),
45535 => conv_std_logic_vector(154, 8),
45536 => conv_std_logic_vector(154, 8),
45537 => conv_std_logic_vector(155, 8),
45538 => conv_std_logic_vector(156, 8),
45539 => conv_std_logic_vector(156, 8),
45540 => conv_std_logic_vector(157, 8),
45541 => conv_std_logic_vector(158, 8),
45542 => conv_std_logic_vector(159, 8),
45543 => conv_std_logic_vector(159, 8),
45544 => conv_std_logic_vector(160, 8),
45545 => conv_std_logic_vector(161, 8),
45546 => conv_std_logic_vector(161, 8),
45547 => conv_std_logic_vector(162, 8),
45548 => conv_std_logic_vector(163, 8),
45549 => conv_std_logic_vector(163, 8),
45550 => conv_std_logic_vector(164, 8),
45551 => conv_std_logic_vector(165, 8),
45552 => conv_std_logic_vector(165, 8),
45553 => conv_std_logic_vector(166, 8),
45554 => conv_std_logic_vector(167, 8),
45555 => conv_std_logic_vector(168, 8),
45556 => conv_std_logic_vector(168, 8),
45557 => conv_std_logic_vector(169, 8),
45558 => conv_std_logic_vector(170, 8),
45559 => conv_std_logic_vector(170, 8),
45560 => conv_std_logic_vector(171, 8),
45561 => conv_std_logic_vector(172, 8),
45562 => conv_std_logic_vector(172, 8),
45563 => conv_std_logic_vector(173, 8),
45564 => conv_std_logic_vector(174, 8),
45565 => conv_std_logic_vector(174, 8),
45566 => conv_std_logic_vector(175, 8),
45567 => conv_std_logic_vector(176, 8),
45568 => conv_std_logic_vector(0, 8),
45569 => conv_std_logic_vector(0, 8),
45570 => conv_std_logic_vector(1, 8),
45571 => conv_std_logic_vector(2, 8),
45572 => conv_std_logic_vector(2, 8),
45573 => conv_std_logic_vector(3, 8),
45574 => conv_std_logic_vector(4, 8),
45575 => conv_std_logic_vector(4, 8),
45576 => conv_std_logic_vector(5, 8),
45577 => conv_std_logic_vector(6, 8),
45578 => conv_std_logic_vector(6, 8),
45579 => conv_std_logic_vector(7, 8),
45580 => conv_std_logic_vector(8, 8),
45581 => conv_std_logic_vector(9, 8),
45582 => conv_std_logic_vector(9, 8),
45583 => conv_std_logic_vector(10, 8),
45584 => conv_std_logic_vector(11, 8),
45585 => conv_std_logic_vector(11, 8),
45586 => conv_std_logic_vector(12, 8),
45587 => conv_std_logic_vector(13, 8),
45588 => conv_std_logic_vector(13, 8),
45589 => conv_std_logic_vector(14, 8),
45590 => conv_std_logic_vector(15, 8),
45591 => conv_std_logic_vector(15, 8),
45592 => conv_std_logic_vector(16, 8),
45593 => conv_std_logic_vector(17, 8),
45594 => conv_std_logic_vector(18, 8),
45595 => conv_std_logic_vector(18, 8),
45596 => conv_std_logic_vector(19, 8),
45597 => conv_std_logic_vector(20, 8),
45598 => conv_std_logic_vector(20, 8),
45599 => conv_std_logic_vector(21, 8),
45600 => conv_std_logic_vector(22, 8),
45601 => conv_std_logic_vector(22, 8),
45602 => conv_std_logic_vector(23, 8),
45603 => conv_std_logic_vector(24, 8),
45604 => conv_std_logic_vector(25, 8),
45605 => conv_std_logic_vector(25, 8),
45606 => conv_std_logic_vector(26, 8),
45607 => conv_std_logic_vector(27, 8),
45608 => conv_std_logic_vector(27, 8),
45609 => conv_std_logic_vector(28, 8),
45610 => conv_std_logic_vector(29, 8),
45611 => conv_std_logic_vector(29, 8),
45612 => conv_std_logic_vector(30, 8),
45613 => conv_std_logic_vector(31, 8),
45614 => conv_std_logic_vector(31, 8),
45615 => conv_std_logic_vector(32, 8),
45616 => conv_std_logic_vector(33, 8),
45617 => conv_std_logic_vector(34, 8),
45618 => conv_std_logic_vector(34, 8),
45619 => conv_std_logic_vector(35, 8),
45620 => conv_std_logic_vector(36, 8),
45621 => conv_std_logic_vector(36, 8),
45622 => conv_std_logic_vector(37, 8),
45623 => conv_std_logic_vector(38, 8),
45624 => conv_std_logic_vector(38, 8),
45625 => conv_std_logic_vector(39, 8),
45626 => conv_std_logic_vector(40, 8),
45627 => conv_std_logic_vector(41, 8),
45628 => conv_std_logic_vector(41, 8),
45629 => conv_std_logic_vector(42, 8),
45630 => conv_std_logic_vector(43, 8),
45631 => conv_std_logic_vector(43, 8),
45632 => conv_std_logic_vector(44, 8),
45633 => conv_std_logic_vector(45, 8),
45634 => conv_std_logic_vector(45, 8),
45635 => conv_std_logic_vector(46, 8),
45636 => conv_std_logic_vector(47, 8),
45637 => conv_std_logic_vector(47, 8),
45638 => conv_std_logic_vector(48, 8),
45639 => conv_std_logic_vector(49, 8),
45640 => conv_std_logic_vector(50, 8),
45641 => conv_std_logic_vector(50, 8),
45642 => conv_std_logic_vector(51, 8),
45643 => conv_std_logic_vector(52, 8),
45644 => conv_std_logic_vector(52, 8),
45645 => conv_std_logic_vector(53, 8),
45646 => conv_std_logic_vector(54, 8),
45647 => conv_std_logic_vector(54, 8),
45648 => conv_std_logic_vector(55, 8),
45649 => conv_std_logic_vector(56, 8),
45650 => conv_std_logic_vector(57, 8),
45651 => conv_std_logic_vector(57, 8),
45652 => conv_std_logic_vector(58, 8),
45653 => conv_std_logic_vector(59, 8),
45654 => conv_std_logic_vector(59, 8),
45655 => conv_std_logic_vector(60, 8),
45656 => conv_std_logic_vector(61, 8),
45657 => conv_std_logic_vector(61, 8),
45658 => conv_std_logic_vector(62, 8),
45659 => conv_std_logic_vector(63, 8),
45660 => conv_std_logic_vector(63, 8),
45661 => conv_std_logic_vector(64, 8),
45662 => conv_std_logic_vector(65, 8),
45663 => conv_std_logic_vector(66, 8),
45664 => conv_std_logic_vector(66, 8),
45665 => conv_std_logic_vector(67, 8),
45666 => conv_std_logic_vector(68, 8),
45667 => conv_std_logic_vector(68, 8),
45668 => conv_std_logic_vector(69, 8),
45669 => conv_std_logic_vector(70, 8),
45670 => conv_std_logic_vector(70, 8),
45671 => conv_std_logic_vector(71, 8),
45672 => conv_std_logic_vector(72, 8),
45673 => conv_std_logic_vector(73, 8),
45674 => conv_std_logic_vector(73, 8),
45675 => conv_std_logic_vector(74, 8),
45676 => conv_std_logic_vector(75, 8),
45677 => conv_std_logic_vector(75, 8),
45678 => conv_std_logic_vector(76, 8),
45679 => conv_std_logic_vector(77, 8),
45680 => conv_std_logic_vector(77, 8),
45681 => conv_std_logic_vector(78, 8),
45682 => conv_std_logic_vector(79, 8),
45683 => conv_std_logic_vector(79, 8),
45684 => conv_std_logic_vector(80, 8),
45685 => conv_std_logic_vector(81, 8),
45686 => conv_std_logic_vector(82, 8),
45687 => conv_std_logic_vector(82, 8),
45688 => conv_std_logic_vector(83, 8),
45689 => conv_std_logic_vector(84, 8),
45690 => conv_std_logic_vector(84, 8),
45691 => conv_std_logic_vector(85, 8),
45692 => conv_std_logic_vector(86, 8),
45693 => conv_std_logic_vector(86, 8),
45694 => conv_std_logic_vector(87, 8),
45695 => conv_std_logic_vector(88, 8),
45696 => conv_std_logic_vector(89, 8),
45697 => conv_std_logic_vector(89, 8),
45698 => conv_std_logic_vector(90, 8),
45699 => conv_std_logic_vector(91, 8),
45700 => conv_std_logic_vector(91, 8),
45701 => conv_std_logic_vector(92, 8),
45702 => conv_std_logic_vector(93, 8),
45703 => conv_std_logic_vector(93, 8),
45704 => conv_std_logic_vector(94, 8),
45705 => conv_std_logic_vector(95, 8),
45706 => conv_std_logic_vector(95, 8),
45707 => conv_std_logic_vector(96, 8),
45708 => conv_std_logic_vector(97, 8),
45709 => conv_std_logic_vector(98, 8),
45710 => conv_std_logic_vector(98, 8),
45711 => conv_std_logic_vector(99, 8),
45712 => conv_std_logic_vector(100, 8),
45713 => conv_std_logic_vector(100, 8),
45714 => conv_std_logic_vector(101, 8),
45715 => conv_std_logic_vector(102, 8),
45716 => conv_std_logic_vector(102, 8),
45717 => conv_std_logic_vector(103, 8),
45718 => conv_std_logic_vector(104, 8),
45719 => conv_std_logic_vector(104, 8),
45720 => conv_std_logic_vector(105, 8),
45721 => conv_std_logic_vector(106, 8),
45722 => conv_std_logic_vector(107, 8),
45723 => conv_std_logic_vector(107, 8),
45724 => conv_std_logic_vector(108, 8),
45725 => conv_std_logic_vector(109, 8),
45726 => conv_std_logic_vector(109, 8),
45727 => conv_std_logic_vector(110, 8),
45728 => conv_std_logic_vector(111, 8),
45729 => conv_std_logic_vector(111, 8),
45730 => conv_std_logic_vector(112, 8),
45731 => conv_std_logic_vector(113, 8),
45732 => conv_std_logic_vector(114, 8),
45733 => conv_std_logic_vector(114, 8),
45734 => conv_std_logic_vector(115, 8),
45735 => conv_std_logic_vector(116, 8),
45736 => conv_std_logic_vector(116, 8),
45737 => conv_std_logic_vector(117, 8),
45738 => conv_std_logic_vector(118, 8),
45739 => conv_std_logic_vector(118, 8),
45740 => conv_std_logic_vector(119, 8),
45741 => conv_std_logic_vector(120, 8),
45742 => conv_std_logic_vector(120, 8),
45743 => conv_std_logic_vector(121, 8),
45744 => conv_std_logic_vector(122, 8),
45745 => conv_std_logic_vector(123, 8),
45746 => conv_std_logic_vector(123, 8),
45747 => conv_std_logic_vector(124, 8),
45748 => conv_std_logic_vector(125, 8),
45749 => conv_std_logic_vector(125, 8),
45750 => conv_std_logic_vector(126, 8),
45751 => conv_std_logic_vector(127, 8),
45752 => conv_std_logic_vector(127, 8),
45753 => conv_std_logic_vector(128, 8),
45754 => conv_std_logic_vector(129, 8),
45755 => conv_std_logic_vector(130, 8),
45756 => conv_std_logic_vector(130, 8),
45757 => conv_std_logic_vector(131, 8),
45758 => conv_std_logic_vector(132, 8),
45759 => conv_std_logic_vector(132, 8),
45760 => conv_std_logic_vector(133, 8),
45761 => conv_std_logic_vector(134, 8),
45762 => conv_std_logic_vector(134, 8),
45763 => conv_std_logic_vector(135, 8),
45764 => conv_std_logic_vector(136, 8),
45765 => conv_std_logic_vector(136, 8),
45766 => conv_std_logic_vector(137, 8),
45767 => conv_std_logic_vector(138, 8),
45768 => conv_std_logic_vector(139, 8),
45769 => conv_std_logic_vector(139, 8),
45770 => conv_std_logic_vector(140, 8),
45771 => conv_std_logic_vector(141, 8),
45772 => conv_std_logic_vector(141, 8),
45773 => conv_std_logic_vector(142, 8),
45774 => conv_std_logic_vector(143, 8),
45775 => conv_std_logic_vector(143, 8),
45776 => conv_std_logic_vector(144, 8),
45777 => conv_std_logic_vector(145, 8),
45778 => conv_std_logic_vector(146, 8),
45779 => conv_std_logic_vector(146, 8),
45780 => conv_std_logic_vector(147, 8),
45781 => conv_std_logic_vector(148, 8),
45782 => conv_std_logic_vector(148, 8),
45783 => conv_std_logic_vector(149, 8),
45784 => conv_std_logic_vector(150, 8),
45785 => conv_std_logic_vector(150, 8),
45786 => conv_std_logic_vector(151, 8),
45787 => conv_std_logic_vector(152, 8),
45788 => conv_std_logic_vector(152, 8),
45789 => conv_std_logic_vector(153, 8),
45790 => conv_std_logic_vector(154, 8),
45791 => conv_std_logic_vector(155, 8),
45792 => conv_std_logic_vector(155, 8),
45793 => conv_std_logic_vector(156, 8),
45794 => conv_std_logic_vector(157, 8),
45795 => conv_std_logic_vector(157, 8),
45796 => conv_std_logic_vector(158, 8),
45797 => conv_std_logic_vector(159, 8),
45798 => conv_std_logic_vector(159, 8),
45799 => conv_std_logic_vector(160, 8),
45800 => conv_std_logic_vector(161, 8),
45801 => conv_std_logic_vector(162, 8),
45802 => conv_std_logic_vector(162, 8),
45803 => conv_std_logic_vector(163, 8),
45804 => conv_std_logic_vector(164, 8),
45805 => conv_std_logic_vector(164, 8),
45806 => conv_std_logic_vector(165, 8),
45807 => conv_std_logic_vector(166, 8),
45808 => conv_std_logic_vector(166, 8),
45809 => conv_std_logic_vector(167, 8),
45810 => conv_std_logic_vector(168, 8),
45811 => conv_std_logic_vector(168, 8),
45812 => conv_std_logic_vector(169, 8),
45813 => conv_std_logic_vector(170, 8),
45814 => conv_std_logic_vector(171, 8),
45815 => conv_std_logic_vector(171, 8),
45816 => conv_std_logic_vector(172, 8),
45817 => conv_std_logic_vector(173, 8),
45818 => conv_std_logic_vector(173, 8),
45819 => conv_std_logic_vector(174, 8),
45820 => conv_std_logic_vector(175, 8),
45821 => conv_std_logic_vector(175, 8),
45822 => conv_std_logic_vector(176, 8),
45823 => conv_std_logic_vector(177, 8),
45824 => conv_std_logic_vector(0, 8),
45825 => conv_std_logic_vector(0, 8),
45826 => conv_std_logic_vector(1, 8),
45827 => conv_std_logic_vector(2, 8),
45828 => conv_std_logic_vector(2, 8),
45829 => conv_std_logic_vector(3, 8),
45830 => conv_std_logic_vector(4, 8),
45831 => conv_std_logic_vector(4, 8),
45832 => conv_std_logic_vector(5, 8),
45833 => conv_std_logic_vector(6, 8),
45834 => conv_std_logic_vector(6, 8),
45835 => conv_std_logic_vector(7, 8),
45836 => conv_std_logic_vector(8, 8),
45837 => conv_std_logic_vector(9, 8),
45838 => conv_std_logic_vector(9, 8),
45839 => conv_std_logic_vector(10, 8),
45840 => conv_std_logic_vector(11, 8),
45841 => conv_std_logic_vector(11, 8),
45842 => conv_std_logic_vector(12, 8),
45843 => conv_std_logic_vector(13, 8),
45844 => conv_std_logic_vector(13, 8),
45845 => conv_std_logic_vector(14, 8),
45846 => conv_std_logic_vector(15, 8),
45847 => conv_std_logic_vector(16, 8),
45848 => conv_std_logic_vector(16, 8),
45849 => conv_std_logic_vector(17, 8),
45850 => conv_std_logic_vector(18, 8),
45851 => conv_std_logic_vector(18, 8),
45852 => conv_std_logic_vector(19, 8),
45853 => conv_std_logic_vector(20, 8),
45854 => conv_std_logic_vector(20, 8),
45855 => conv_std_logic_vector(21, 8),
45856 => conv_std_logic_vector(22, 8),
45857 => conv_std_logic_vector(23, 8),
45858 => conv_std_logic_vector(23, 8),
45859 => conv_std_logic_vector(24, 8),
45860 => conv_std_logic_vector(25, 8),
45861 => conv_std_logic_vector(25, 8),
45862 => conv_std_logic_vector(26, 8),
45863 => conv_std_logic_vector(27, 8),
45864 => conv_std_logic_vector(27, 8),
45865 => conv_std_logic_vector(28, 8),
45866 => conv_std_logic_vector(29, 8),
45867 => conv_std_logic_vector(30, 8),
45868 => conv_std_logic_vector(30, 8),
45869 => conv_std_logic_vector(31, 8),
45870 => conv_std_logic_vector(32, 8),
45871 => conv_std_logic_vector(32, 8),
45872 => conv_std_logic_vector(33, 8),
45873 => conv_std_logic_vector(34, 8),
45874 => conv_std_logic_vector(34, 8),
45875 => conv_std_logic_vector(35, 8),
45876 => conv_std_logic_vector(36, 8),
45877 => conv_std_logic_vector(37, 8),
45878 => conv_std_logic_vector(37, 8),
45879 => conv_std_logic_vector(38, 8),
45880 => conv_std_logic_vector(39, 8),
45881 => conv_std_logic_vector(39, 8),
45882 => conv_std_logic_vector(40, 8),
45883 => conv_std_logic_vector(41, 8),
45884 => conv_std_logic_vector(41, 8),
45885 => conv_std_logic_vector(42, 8),
45886 => conv_std_logic_vector(43, 8),
45887 => conv_std_logic_vector(44, 8),
45888 => conv_std_logic_vector(44, 8),
45889 => conv_std_logic_vector(45, 8),
45890 => conv_std_logic_vector(46, 8),
45891 => conv_std_logic_vector(46, 8),
45892 => conv_std_logic_vector(47, 8),
45893 => conv_std_logic_vector(48, 8),
45894 => conv_std_logic_vector(48, 8),
45895 => conv_std_logic_vector(49, 8),
45896 => conv_std_logic_vector(50, 8),
45897 => conv_std_logic_vector(51, 8),
45898 => conv_std_logic_vector(51, 8),
45899 => conv_std_logic_vector(52, 8),
45900 => conv_std_logic_vector(53, 8),
45901 => conv_std_logic_vector(53, 8),
45902 => conv_std_logic_vector(54, 8),
45903 => conv_std_logic_vector(55, 8),
45904 => conv_std_logic_vector(55, 8),
45905 => conv_std_logic_vector(56, 8),
45906 => conv_std_logic_vector(57, 8),
45907 => conv_std_logic_vector(58, 8),
45908 => conv_std_logic_vector(58, 8),
45909 => conv_std_logic_vector(59, 8),
45910 => conv_std_logic_vector(60, 8),
45911 => conv_std_logic_vector(60, 8),
45912 => conv_std_logic_vector(61, 8),
45913 => conv_std_logic_vector(62, 8),
45914 => conv_std_logic_vector(62, 8),
45915 => conv_std_logic_vector(63, 8),
45916 => conv_std_logic_vector(64, 8),
45917 => conv_std_logic_vector(65, 8),
45918 => conv_std_logic_vector(65, 8),
45919 => conv_std_logic_vector(66, 8),
45920 => conv_std_logic_vector(67, 8),
45921 => conv_std_logic_vector(67, 8),
45922 => conv_std_logic_vector(68, 8),
45923 => conv_std_logic_vector(69, 8),
45924 => conv_std_logic_vector(69, 8),
45925 => conv_std_logic_vector(70, 8),
45926 => conv_std_logic_vector(71, 8),
45927 => conv_std_logic_vector(72, 8),
45928 => conv_std_logic_vector(72, 8),
45929 => conv_std_logic_vector(73, 8),
45930 => conv_std_logic_vector(74, 8),
45931 => conv_std_logic_vector(74, 8),
45932 => conv_std_logic_vector(75, 8),
45933 => conv_std_logic_vector(76, 8),
45934 => conv_std_logic_vector(76, 8),
45935 => conv_std_logic_vector(77, 8),
45936 => conv_std_logic_vector(78, 8),
45937 => conv_std_logic_vector(79, 8),
45938 => conv_std_logic_vector(79, 8),
45939 => conv_std_logic_vector(80, 8),
45940 => conv_std_logic_vector(81, 8),
45941 => conv_std_logic_vector(81, 8),
45942 => conv_std_logic_vector(82, 8),
45943 => conv_std_logic_vector(83, 8),
45944 => conv_std_logic_vector(83, 8),
45945 => conv_std_logic_vector(84, 8),
45946 => conv_std_logic_vector(85, 8),
45947 => conv_std_logic_vector(86, 8),
45948 => conv_std_logic_vector(86, 8),
45949 => conv_std_logic_vector(87, 8),
45950 => conv_std_logic_vector(88, 8),
45951 => conv_std_logic_vector(88, 8),
45952 => conv_std_logic_vector(89, 8),
45953 => conv_std_logic_vector(90, 8),
45954 => conv_std_logic_vector(90, 8),
45955 => conv_std_logic_vector(91, 8),
45956 => conv_std_logic_vector(92, 8),
45957 => conv_std_logic_vector(92, 8),
45958 => conv_std_logic_vector(93, 8),
45959 => conv_std_logic_vector(94, 8),
45960 => conv_std_logic_vector(95, 8),
45961 => conv_std_logic_vector(95, 8),
45962 => conv_std_logic_vector(96, 8),
45963 => conv_std_logic_vector(97, 8),
45964 => conv_std_logic_vector(97, 8),
45965 => conv_std_logic_vector(98, 8),
45966 => conv_std_logic_vector(99, 8),
45967 => conv_std_logic_vector(99, 8),
45968 => conv_std_logic_vector(100, 8),
45969 => conv_std_logic_vector(101, 8),
45970 => conv_std_logic_vector(102, 8),
45971 => conv_std_logic_vector(102, 8),
45972 => conv_std_logic_vector(103, 8),
45973 => conv_std_logic_vector(104, 8),
45974 => conv_std_logic_vector(104, 8),
45975 => conv_std_logic_vector(105, 8),
45976 => conv_std_logic_vector(106, 8),
45977 => conv_std_logic_vector(106, 8),
45978 => conv_std_logic_vector(107, 8),
45979 => conv_std_logic_vector(108, 8),
45980 => conv_std_logic_vector(109, 8),
45981 => conv_std_logic_vector(109, 8),
45982 => conv_std_logic_vector(110, 8),
45983 => conv_std_logic_vector(111, 8),
45984 => conv_std_logic_vector(111, 8),
45985 => conv_std_logic_vector(112, 8),
45986 => conv_std_logic_vector(113, 8),
45987 => conv_std_logic_vector(113, 8),
45988 => conv_std_logic_vector(114, 8),
45989 => conv_std_logic_vector(115, 8),
45990 => conv_std_logic_vector(116, 8),
45991 => conv_std_logic_vector(116, 8),
45992 => conv_std_logic_vector(117, 8),
45993 => conv_std_logic_vector(118, 8),
45994 => conv_std_logic_vector(118, 8),
45995 => conv_std_logic_vector(119, 8),
45996 => conv_std_logic_vector(120, 8),
45997 => conv_std_logic_vector(120, 8),
45998 => conv_std_logic_vector(121, 8),
45999 => conv_std_logic_vector(122, 8),
46000 => conv_std_logic_vector(123, 8),
46001 => conv_std_logic_vector(123, 8),
46002 => conv_std_logic_vector(124, 8),
46003 => conv_std_logic_vector(125, 8),
46004 => conv_std_logic_vector(125, 8),
46005 => conv_std_logic_vector(126, 8),
46006 => conv_std_logic_vector(127, 8),
46007 => conv_std_logic_vector(127, 8),
46008 => conv_std_logic_vector(128, 8),
46009 => conv_std_logic_vector(129, 8),
46010 => conv_std_logic_vector(130, 8),
46011 => conv_std_logic_vector(130, 8),
46012 => conv_std_logic_vector(131, 8),
46013 => conv_std_logic_vector(132, 8),
46014 => conv_std_logic_vector(132, 8),
46015 => conv_std_logic_vector(133, 8),
46016 => conv_std_logic_vector(134, 8),
46017 => conv_std_logic_vector(134, 8),
46018 => conv_std_logic_vector(135, 8),
46019 => conv_std_logic_vector(136, 8),
46020 => conv_std_logic_vector(137, 8),
46021 => conv_std_logic_vector(137, 8),
46022 => conv_std_logic_vector(138, 8),
46023 => conv_std_logic_vector(139, 8),
46024 => conv_std_logic_vector(139, 8),
46025 => conv_std_logic_vector(140, 8),
46026 => conv_std_logic_vector(141, 8),
46027 => conv_std_logic_vector(141, 8),
46028 => conv_std_logic_vector(142, 8),
46029 => conv_std_logic_vector(143, 8),
46030 => conv_std_logic_vector(144, 8),
46031 => conv_std_logic_vector(144, 8),
46032 => conv_std_logic_vector(145, 8),
46033 => conv_std_logic_vector(146, 8),
46034 => conv_std_logic_vector(146, 8),
46035 => conv_std_logic_vector(147, 8),
46036 => conv_std_logic_vector(148, 8),
46037 => conv_std_logic_vector(148, 8),
46038 => conv_std_logic_vector(149, 8),
46039 => conv_std_logic_vector(150, 8),
46040 => conv_std_logic_vector(151, 8),
46041 => conv_std_logic_vector(151, 8),
46042 => conv_std_logic_vector(152, 8),
46043 => conv_std_logic_vector(153, 8),
46044 => conv_std_logic_vector(153, 8),
46045 => conv_std_logic_vector(154, 8),
46046 => conv_std_logic_vector(155, 8),
46047 => conv_std_logic_vector(155, 8),
46048 => conv_std_logic_vector(156, 8),
46049 => conv_std_logic_vector(157, 8),
46050 => conv_std_logic_vector(158, 8),
46051 => conv_std_logic_vector(158, 8),
46052 => conv_std_logic_vector(159, 8),
46053 => conv_std_logic_vector(160, 8),
46054 => conv_std_logic_vector(160, 8),
46055 => conv_std_logic_vector(161, 8),
46056 => conv_std_logic_vector(162, 8),
46057 => conv_std_logic_vector(162, 8),
46058 => conv_std_logic_vector(163, 8),
46059 => conv_std_logic_vector(164, 8),
46060 => conv_std_logic_vector(165, 8),
46061 => conv_std_logic_vector(165, 8),
46062 => conv_std_logic_vector(166, 8),
46063 => conv_std_logic_vector(167, 8),
46064 => conv_std_logic_vector(167, 8),
46065 => conv_std_logic_vector(168, 8),
46066 => conv_std_logic_vector(169, 8),
46067 => conv_std_logic_vector(169, 8),
46068 => conv_std_logic_vector(170, 8),
46069 => conv_std_logic_vector(171, 8),
46070 => conv_std_logic_vector(172, 8),
46071 => conv_std_logic_vector(172, 8),
46072 => conv_std_logic_vector(173, 8),
46073 => conv_std_logic_vector(174, 8),
46074 => conv_std_logic_vector(174, 8),
46075 => conv_std_logic_vector(175, 8),
46076 => conv_std_logic_vector(176, 8),
46077 => conv_std_logic_vector(176, 8),
46078 => conv_std_logic_vector(177, 8),
46079 => conv_std_logic_vector(178, 8),
46080 => conv_std_logic_vector(0, 8),
46081 => conv_std_logic_vector(0, 8),
46082 => conv_std_logic_vector(1, 8),
46083 => conv_std_logic_vector(2, 8),
46084 => conv_std_logic_vector(2, 8),
46085 => conv_std_logic_vector(3, 8),
46086 => conv_std_logic_vector(4, 8),
46087 => conv_std_logic_vector(4, 8),
46088 => conv_std_logic_vector(5, 8),
46089 => conv_std_logic_vector(6, 8),
46090 => conv_std_logic_vector(7, 8),
46091 => conv_std_logic_vector(7, 8),
46092 => conv_std_logic_vector(8, 8),
46093 => conv_std_logic_vector(9, 8),
46094 => conv_std_logic_vector(9, 8),
46095 => conv_std_logic_vector(10, 8),
46096 => conv_std_logic_vector(11, 8),
46097 => conv_std_logic_vector(11, 8),
46098 => conv_std_logic_vector(12, 8),
46099 => conv_std_logic_vector(13, 8),
46100 => conv_std_logic_vector(14, 8),
46101 => conv_std_logic_vector(14, 8),
46102 => conv_std_logic_vector(15, 8),
46103 => conv_std_logic_vector(16, 8),
46104 => conv_std_logic_vector(16, 8),
46105 => conv_std_logic_vector(17, 8),
46106 => conv_std_logic_vector(18, 8),
46107 => conv_std_logic_vector(18, 8),
46108 => conv_std_logic_vector(19, 8),
46109 => conv_std_logic_vector(20, 8),
46110 => conv_std_logic_vector(21, 8),
46111 => conv_std_logic_vector(21, 8),
46112 => conv_std_logic_vector(22, 8),
46113 => conv_std_logic_vector(23, 8),
46114 => conv_std_logic_vector(23, 8),
46115 => conv_std_logic_vector(24, 8),
46116 => conv_std_logic_vector(25, 8),
46117 => conv_std_logic_vector(26, 8),
46118 => conv_std_logic_vector(26, 8),
46119 => conv_std_logic_vector(27, 8),
46120 => conv_std_logic_vector(28, 8),
46121 => conv_std_logic_vector(28, 8),
46122 => conv_std_logic_vector(29, 8),
46123 => conv_std_logic_vector(30, 8),
46124 => conv_std_logic_vector(30, 8),
46125 => conv_std_logic_vector(31, 8),
46126 => conv_std_logic_vector(32, 8),
46127 => conv_std_logic_vector(33, 8),
46128 => conv_std_logic_vector(33, 8),
46129 => conv_std_logic_vector(34, 8),
46130 => conv_std_logic_vector(35, 8),
46131 => conv_std_logic_vector(35, 8),
46132 => conv_std_logic_vector(36, 8),
46133 => conv_std_logic_vector(37, 8),
46134 => conv_std_logic_vector(37, 8),
46135 => conv_std_logic_vector(38, 8),
46136 => conv_std_logic_vector(39, 8),
46137 => conv_std_logic_vector(40, 8),
46138 => conv_std_logic_vector(40, 8),
46139 => conv_std_logic_vector(41, 8),
46140 => conv_std_logic_vector(42, 8),
46141 => conv_std_logic_vector(42, 8),
46142 => conv_std_logic_vector(43, 8),
46143 => conv_std_logic_vector(44, 8),
46144 => conv_std_logic_vector(45, 8),
46145 => conv_std_logic_vector(45, 8),
46146 => conv_std_logic_vector(46, 8),
46147 => conv_std_logic_vector(47, 8),
46148 => conv_std_logic_vector(47, 8),
46149 => conv_std_logic_vector(48, 8),
46150 => conv_std_logic_vector(49, 8),
46151 => conv_std_logic_vector(49, 8),
46152 => conv_std_logic_vector(50, 8),
46153 => conv_std_logic_vector(51, 8),
46154 => conv_std_logic_vector(52, 8),
46155 => conv_std_logic_vector(52, 8),
46156 => conv_std_logic_vector(53, 8),
46157 => conv_std_logic_vector(54, 8),
46158 => conv_std_logic_vector(54, 8),
46159 => conv_std_logic_vector(55, 8),
46160 => conv_std_logic_vector(56, 8),
46161 => conv_std_logic_vector(56, 8),
46162 => conv_std_logic_vector(57, 8),
46163 => conv_std_logic_vector(58, 8),
46164 => conv_std_logic_vector(59, 8),
46165 => conv_std_logic_vector(59, 8),
46166 => conv_std_logic_vector(60, 8),
46167 => conv_std_logic_vector(61, 8),
46168 => conv_std_logic_vector(61, 8),
46169 => conv_std_logic_vector(62, 8),
46170 => conv_std_logic_vector(63, 8),
46171 => conv_std_logic_vector(63, 8),
46172 => conv_std_logic_vector(64, 8),
46173 => conv_std_logic_vector(65, 8),
46174 => conv_std_logic_vector(66, 8),
46175 => conv_std_logic_vector(66, 8),
46176 => conv_std_logic_vector(67, 8),
46177 => conv_std_logic_vector(68, 8),
46178 => conv_std_logic_vector(68, 8),
46179 => conv_std_logic_vector(69, 8),
46180 => conv_std_logic_vector(70, 8),
46181 => conv_std_logic_vector(71, 8),
46182 => conv_std_logic_vector(71, 8),
46183 => conv_std_logic_vector(72, 8),
46184 => conv_std_logic_vector(73, 8),
46185 => conv_std_logic_vector(73, 8),
46186 => conv_std_logic_vector(74, 8),
46187 => conv_std_logic_vector(75, 8),
46188 => conv_std_logic_vector(75, 8),
46189 => conv_std_logic_vector(76, 8),
46190 => conv_std_logic_vector(77, 8),
46191 => conv_std_logic_vector(78, 8),
46192 => conv_std_logic_vector(78, 8),
46193 => conv_std_logic_vector(79, 8),
46194 => conv_std_logic_vector(80, 8),
46195 => conv_std_logic_vector(80, 8),
46196 => conv_std_logic_vector(81, 8),
46197 => conv_std_logic_vector(82, 8),
46198 => conv_std_logic_vector(82, 8),
46199 => conv_std_logic_vector(83, 8),
46200 => conv_std_logic_vector(84, 8),
46201 => conv_std_logic_vector(85, 8),
46202 => conv_std_logic_vector(85, 8),
46203 => conv_std_logic_vector(86, 8),
46204 => conv_std_logic_vector(87, 8),
46205 => conv_std_logic_vector(87, 8),
46206 => conv_std_logic_vector(88, 8),
46207 => conv_std_logic_vector(89, 8),
46208 => conv_std_logic_vector(90, 8),
46209 => conv_std_logic_vector(90, 8),
46210 => conv_std_logic_vector(91, 8),
46211 => conv_std_logic_vector(92, 8),
46212 => conv_std_logic_vector(92, 8),
46213 => conv_std_logic_vector(93, 8),
46214 => conv_std_logic_vector(94, 8),
46215 => conv_std_logic_vector(94, 8),
46216 => conv_std_logic_vector(95, 8),
46217 => conv_std_logic_vector(96, 8),
46218 => conv_std_logic_vector(97, 8),
46219 => conv_std_logic_vector(97, 8),
46220 => conv_std_logic_vector(98, 8),
46221 => conv_std_logic_vector(99, 8),
46222 => conv_std_logic_vector(99, 8),
46223 => conv_std_logic_vector(100, 8),
46224 => conv_std_logic_vector(101, 8),
46225 => conv_std_logic_vector(101, 8),
46226 => conv_std_logic_vector(102, 8),
46227 => conv_std_logic_vector(103, 8),
46228 => conv_std_logic_vector(104, 8),
46229 => conv_std_logic_vector(104, 8),
46230 => conv_std_logic_vector(105, 8),
46231 => conv_std_logic_vector(106, 8),
46232 => conv_std_logic_vector(106, 8),
46233 => conv_std_logic_vector(107, 8),
46234 => conv_std_logic_vector(108, 8),
46235 => conv_std_logic_vector(108, 8),
46236 => conv_std_logic_vector(109, 8),
46237 => conv_std_logic_vector(110, 8),
46238 => conv_std_logic_vector(111, 8),
46239 => conv_std_logic_vector(111, 8),
46240 => conv_std_logic_vector(112, 8),
46241 => conv_std_logic_vector(113, 8),
46242 => conv_std_logic_vector(113, 8),
46243 => conv_std_logic_vector(114, 8),
46244 => conv_std_logic_vector(115, 8),
46245 => conv_std_logic_vector(116, 8),
46246 => conv_std_logic_vector(116, 8),
46247 => conv_std_logic_vector(117, 8),
46248 => conv_std_logic_vector(118, 8),
46249 => conv_std_logic_vector(118, 8),
46250 => conv_std_logic_vector(119, 8),
46251 => conv_std_logic_vector(120, 8),
46252 => conv_std_logic_vector(120, 8),
46253 => conv_std_logic_vector(121, 8),
46254 => conv_std_logic_vector(122, 8),
46255 => conv_std_logic_vector(123, 8),
46256 => conv_std_logic_vector(123, 8),
46257 => conv_std_logic_vector(124, 8),
46258 => conv_std_logic_vector(125, 8),
46259 => conv_std_logic_vector(125, 8),
46260 => conv_std_logic_vector(126, 8),
46261 => conv_std_logic_vector(127, 8),
46262 => conv_std_logic_vector(127, 8),
46263 => conv_std_logic_vector(128, 8),
46264 => conv_std_logic_vector(129, 8),
46265 => conv_std_logic_vector(130, 8),
46266 => conv_std_logic_vector(130, 8),
46267 => conv_std_logic_vector(131, 8),
46268 => conv_std_logic_vector(132, 8),
46269 => conv_std_logic_vector(132, 8),
46270 => conv_std_logic_vector(133, 8),
46271 => conv_std_logic_vector(134, 8),
46272 => conv_std_logic_vector(135, 8),
46273 => conv_std_logic_vector(135, 8),
46274 => conv_std_logic_vector(136, 8),
46275 => conv_std_logic_vector(137, 8),
46276 => conv_std_logic_vector(137, 8),
46277 => conv_std_logic_vector(138, 8),
46278 => conv_std_logic_vector(139, 8),
46279 => conv_std_logic_vector(139, 8),
46280 => conv_std_logic_vector(140, 8),
46281 => conv_std_logic_vector(141, 8),
46282 => conv_std_logic_vector(142, 8),
46283 => conv_std_logic_vector(142, 8),
46284 => conv_std_logic_vector(143, 8),
46285 => conv_std_logic_vector(144, 8),
46286 => conv_std_logic_vector(144, 8),
46287 => conv_std_logic_vector(145, 8),
46288 => conv_std_logic_vector(146, 8),
46289 => conv_std_logic_vector(146, 8),
46290 => conv_std_logic_vector(147, 8),
46291 => conv_std_logic_vector(148, 8),
46292 => conv_std_logic_vector(149, 8),
46293 => conv_std_logic_vector(149, 8),
46294 => conv_std_logic_vector(150, 8),
46295 => conv_std_logic_vector(151, 8),
46296 => conv_std_logic_vector(151, 8),
46297 => conv_std_logic_vector(152, 8),
46298 => conv_std_logic_vector(153, 8),
46299 => conv_std_logic_vector(153, 8),
46300 => conv_std_logic_vector(154, 8),
46301 => conv_std_logic_vector(155, 8),
46302 => conv_std_logic_vector(156, 8),
46303 => conv_std_logic_vector(156, 8),
46304 => conv_std_logic_vector(157, 8),
46305 => conv_std_logic_vector(158, 8),
46306 => conv_std_logic_vector(158, 8),
46307 => conv_std_logic_vector(159, 8),
46308 => conv_std_logic_vector(160, 8),
46309 => conv_std_logic_vector(161, 8),
46310 => conv_std_logic_vector(161, 8),
46311 => conv_std_logic_vector(162, 8),
46312 => conv_std_logic_vector(163, 8),
46313 => conv_std_logic_vector(163, 8),
46314 => conv_std_logic_vector(164, 8),
46315 => conv_std_logic_vector(165, 8),
46316 => conv_std_logic_vector(165, 8),
46317 => conv_std_logic_vector(166, 8),
46318 => conv_std_logic_vector(167, 8),
46319 => conv_std_logic_vector(168, 8),
46320 => conv_std_logic_vector(168, 8),
46321 => conv_std_logic_vector(169, 8),
46322 => conv_std_logic_vector(170, 8),
46323 => conv_std_logic_vector(170, 8),
46324 => conv_std_logic_vector(171, 8),
46325 => conv_std_logic_vector(172, 8),
46326 => conv_std_logic_vector(172, 8),
46327 => conv_std_logic_vector(173, 8),
46328 => conv_std_logic_vector(174, 8),
46329 => conv_std_logic_vector(175, 8),
46330 => conv_std_logic_vector(175, 8),
46331 => conv_std_logic_vector(176, 8),
46332 => conv_std_logic_vector(177, 8),
46333 => conv_std_logic_vector(177, 8),
46334 => conv_std_logic_vector(178, 8),
46335 => conv_std_logic_vector(179, 8),
46336 => conv_std_logic_vector(0, 8),
46337 => conv_std_logic_vector(0, 8),
46338 => conv_std_logic_vector(1, 8),
46339 => conv_std_logic_vector(2, 8),
46340 => conv_std_logic_vector(2, 8),
46341 => conv_std_logic_vector(3, 8),
46342 => conv_std_logic_vector(4, 8),
46343 => conv_std_logic_vector(4, 8),
46344 => conv_std_logic_vector(5, 8),
46345 => conv_std_logic_vector(6, 8),
46346 => conv_std_logic_vector(7, 8),
46347 => conv_std_logic_vector(7, 8),
46348 => conv_std_logic_vector(8, 8),
46349 => conv_std_logic_vector(9, 8),
46350 => conv_std_logic_vector(9, 8),
46351 => conv_std_logic_vector(10, 8),
46352 => conv_std_logic_vector(11, 8),
46353 => conv_std_logic_vector(12, 8),
46354 => conv_std_logic_vector(12, 8),
46355 => conv_std_logic_vector(13, 8),
46356 => conv_std_logic_vector(14, 8),
46357 => conv_std_logic_vector(14, 8),
46358 => conv_std_logic_vector(15, 8),
46359 => conv_std_logic_vector(16, 8),
46360 => conv_std_logic_vector(16, 8),
46361 => conv_std_logic_vector(17, 8),
46362 => conv_std_logic_vector(18, 8),
46363 => conv_std_logic_vector(19, 8),
46364 => conv_std_logic_vector(19, 8),
46365 => conv_std_logic_vector(20, 8),
46366 => conv_std_logic_vector(21, 8),
46367 => conv_std_logic_vector(21, 8),
46368 => conv_std_logic_vector(22, 8),
46369 => conv_std_logic_vector(23, 8),
46370 => conv_std_logic_vector(24, 8),
46371 => conv_std_logic_vector(24, 8),
46372 => conv_std_logic_vector(25, 8),
46373 => conv_std_logic_vector(26, 8),
46374 => conv_std_logic_vector(26, 8),
46375 => conv_std_logic_vector(27, 8),
46376 => conv_std_logic_vector(28, 8),
46377 => conv_std_logic_vector(28, 8),
46378 => conv_std_logic_vector(29, 8),
46379 => conv_std_logic_vector(30, 8),
46380 => conv_std_logic_vector(31, 8),
46381 => conv_std_logic_vector(31, 8),
46382 => conv_std_logic_vector(32, 8),
46383 => conv_std_logic_vector(33, 8),
46384 => conv_std_logic_vector(33, 8),
46385 => conv_std_logic_vector(34, 8),
46386 => conv_std_logic_vector(35, 8),
46387 => conv_std_logic_vector(36, 8),
46388 => conv_std_logic_vector(36, 8),
46389 => conv_std_logic_vector(37, 8),
46390 => conv_std_logic_vector(38, 8),
46391 => conv_std_logic_vector(38, 8),
46392 => conv_std_logic_vector(39, 8),
46393 => conv_std_logic_vector(40, 8),
46394 => conv_std_logic_vector(41, 8),
46395 => conv_std_logic_vector(41, 8),
46396 => conv_std_logic_vector(42, 8),
46397 => conv_std_logic_vector(43, 8),
46398 => conv_std_logic_vector(43, 8),
46399 => conv_std_logic_vector(44, 8),
46400 => conv_std_logic_vector(45, 8),
46401 => conv_std_logic_vector(45, 8),
46402 => conv_std_logic_vector(46, 8),
46403 => conv_std_logic_vector(47, 8),
46404 => conv_std_logic_vector(48, 8),
46405 => conv_std_logic_vector(48, 8),
46406 => conv_std_logic_vector(49, 8),
46407 => conv_std_logic_vector(50, 8),
46408 => conv_std_logic_vector(50, 8),
46409 => conv_std_logic_vector(51, 8),
46410 => conv_std_logic_vector(52, 8),
46411 => conv_std_logic_vector(53, 8),
46412 => conv_std_logic_vector(53, 8),
46413 => conv_std_logic_vector(54, 8),
46414 => conv_std_logic_vector(55, 8),
46415 => conv_std_logic_vector(55, 8),
46416 => conv_std_logic_vector(56, 8),
46417 => conv_std_logic_vector(57, 8),
46418 => conv_std_logic_vector(57, 8),
46419 => conv_std_logic_vector(58, 8),
46420 => conv_std_logic_vector(59, 8),
46421 => conv_std_logic_vector(60, 8),
46422 => conv_std_logic_vector(60, 8),
46423 => conv_std_logic_vector(61, 8),
46424 => conv_std_logic_vector(62, 8),
46425 => conv_std_logic_vector(62, 8),
46426 => conv_std_logic_vector(63, 8),
46427 => conv_std_logic_vector(64, 8),
46428 => conv_std_logic_vector(65, 8),
46429 => conv_std_logic_vector(65, 8),
46430 => conv_std_logic_vector(66, 8),
46431 => conv_std_logic_vector(67, 8),
46432 => conv_std_logic_vector(67, 8),
46433 => conv_std_logic_vector(68, 8),
46434 => conv_std_logic_vector(69, 8),
46435 => conv_std_logic_vector(69, 8),
46436 => conv_std_logic_vector(70, 8),
46437 => conv_std_logic_vector(71, 8),
46438 => conv_std_logic_vector(72, 8),
46439 => conv_std_logic_vector(72, 8),
46440 => conv_std_logic_vector(73, 8),
46441 => conv_std_logic_vector(74, 8),
46442 => conv_std_logic_vector(74, 8),
46443 => conv_std_logic_vector(75, 8),
46444 => conv_std_logic_vector(76, 8),
46445 => conv_std_logic_vector(77, 8),
46446 => conv_std_logic_vector(77, 8),
46447 => conv_std_logic_vector(78, 8),
46448 => conv_std_logic_vector(79, 8),
46449 => conv_std_logic_vector(79, 8),
46450 => conv_std_logic_vector(80, 8),
46451 => conv_std_logic_vector(81, 8),
46452 => conv_std_logic_vector(82, 8),
46453 => conv_std_logic_vector(82, 8),
46454 => conv_std_logic_vector(83, 8),
46455 => conv_std_logic_vector(84, 8),
46456 => conv_std_logic_vector(84, 8),
46457 => conv_std_logic_vector(85, 8),
46458 => conv_std_logic_vector(86, 8),
46459 => conv_std_logic_vector(86, 8),
46460 => conv_std_logic_vector(87, 8),
46461 => conv_std_logic_vector(88, 8),
46462 => conv_std_logic_vector(89, 8),
46463 => conv_std_logic_vector(89, 8),
46464 => conv_std_logic_vector(90, 8),
46465 => conv_std_logic_vector(91, 8),
46466 => conv_std_logic_vector(91, 8),
46467 => conv_std_logic_vector(92, 8),
46468 => conv_std_logic_vector(93, 8),
46469 => conv_std_logic_vector(94, 8),
46470 => conv_std_logic_vector(94, 8),
46471 => conv_std_logic_vector(95, 8),
46472 => conv_std_logic_vector(96, 8),
46473 => conv_std_logic_vector(96, 8),
46474 => conv_std_logic_vector(97, 8),
46475 => conv_std_logic_vector(98, 8),
46476 => conv_std_logic_vector(98, 8),
46477 => conv_std_logic_vector(99, 8),
46478 => conv_std_logic_vector(100, 8),
46479 => conv_std_logic_vector(101, 8),
46480 => conv_std_logic_vector(101, 8),
46481 => conv_std_logic_vector(102, 8),
46482 => conv_std_logic_vector(103, 8),
46483 => conv_std_logic_vector(103, 8),
46484 => conv_std_logic_vector(104, 8),
46485 => conv_std_logic_vector(105, 8),
46486 => conv_std_logic_vector(106, 8),
46487 => conv_std_logic_vector(106, 8),
46488 => conv_std_logic_vector(107, 8),
46489 => conv_std_logic_vector(108, 8),
46490 => conv_std_logic_vector(108, 8),
46491 => conv_std_logic_vector(109, 8),
46492 => conv_std_logic_vector(110, 8),
46493 => conv_std_logic_vector(111, 8),
46494 => conv_std_logic_vector(111, 8),
46495 => conv_std_logic_vector(112, 8),
46496 => conv_std_logic_vector(113, 8),
46497 => conv_std_logic_vector(113, 8),
46498 => conv_std_logic_vector(114, 8),
46499 => conv_std_logic_vector(115, 8),
46500 => conv_std_logic_vector(115, 8),
46501 => conv_std_logic_vector(116, 8),
46502 => conv_std_logic_vector(117, 8),
46503 => conv_std_logic_vector(118, 8),
46504 => conv_std_logic_vector(118, 8),
46505 => conv_std_logic_vector(119, 8),
46506 => conv_std_logic_vector(120, 8),
46507 => conv_std_logic_vector(120, 8),
46508 => conv_std_logic_vector(121, 8),
46509 => conv_std_logic_vector(122, 8),
46510 => conv_std_logic_vector(123, 8),
46511 => conv_std_logic_vector(123, 8),
46512 => conv_std_logic_vector(124, 8),
46513 => conv_std_logic_vector(125, 8),
46514 => conv_std_logic_vector(125, 8),
46515 => conv_std_logic_vector(126, 8),
46516 => conv_std_logic_vector(127, 8),
46517 => conv_std_logic_vector(127, 8),
46518 => conv_std_logic_vector(128, 8),
46519 => conv_std_logic_vector(129, 8),
46520 => conv_std_logic_vector(130, 8),
46521 => conv_std_logic_vector(130, 8),
46522 => conv_std_logic_vector(131, 8),
46523 => conv_std_logic_vector(132, 8),
46524 => conv_std_logic_vector(132, 8),
46525 => conv_std_logic_vector(133, 8),
46526 => conv_std_logic_vector(134, 8),
46527 => conv_std_logic_vector(135, 8),
46528 => conv_std_logic_vector(135, 8),
46529 => conv_std_logic_vector(136, 8),
46530 => conv_std_logic_vector(137, 8),
46531 => conv_std_logic_vector(137, 8),
46532 => conv_std_logic_vector(138, 8),
46533 => conv_std_logic_vector(139, 8),
46534 => conv_std_logic_vector(139, 8),
46535 => conv_std_logic_vector(140, 8),
46536 => conv_std_logic_vector(141, 8),
46537 => conv_std_logic_vector(142, 8),
46538 => conv_std_logic_vector(142, 8),
46539 => conv_std_logic_vector(143, 8),
46540 => conv_std_logic_vector(144, 8),
46541 => conv_std_logic_vector(144, 8),
46542 => conv_std_logic_vector(145, 8),
46543 => conv_std_logic_vector(146, 8),
46544 => conv_std_logic_vector(147, 8),
46545 => conv_std_logic_vector(147, 8),
46546 => conv_std_logic_vector(148, 8),
46547 => conv_std_logic_vector(149, 8),
46548 => conv_std_logic_vector(149, 8),
46549 => conv_std_logic_vector(150, 8),
46550 => conv_std_logic_vector(151, 8),
46551 => conv_std_logic_vector(152, 8),
46552 => conv_std_logic_vector(152, 8),
46553 => conv_std_logic_vector(153, 8),
46554 => conv_std_logic_vector(154, 8),
46555 => conv_std_logic_vector(154, 8),
46556 => conv_std_logic_vector(155, 8),
46557 => conv_std_logic_vector(156, 8),
46558 => conv_std_logic_vector(156, 8),
46559 => conv_std_logic_vector(157, 8),
46560 => conv_std_logic_vector(158, 8),
46561 => conv_std_logic_vector(159, 8),
46562 => conv_std_logic_vector(159, 8),
46563 => conv_std_logic_vector(160, 8),
46564 => conv_std_logic_vector(161, 8),
46565 => conv_std_logic_vector(161, 8),
46566 => conv_std_logic_vector(162, 8),
46567 => conv_std_logic_vector(163, 8),
46568 => conv_std_logic_vector(164, 8),
46569 => conv_std_logic_vector(164, 8),
46570 => conv_std_logic_vector(165, 8),
46571 => conv_std_logic_vector(166, 8),
46572 => conv_std_logic_vector(166, 8),
46573 => conv_std_logic_vector(167, 8),
46574 => conv_std_logic_vector(168, 8),
46575 => conv_std_logic_vector(168, 8),
46576 => conv_std_logic_vector(169, 8),
46577 => conv_std_logic_vector(170, 8),
46578 => conv_std_logic_vector(171, 8),
46579 => conv_std_logic_vector(171, 8),
46580 => conv_std_logic_vector(172, 8),
46581 => conv_std_logic_vector(173, 8),
46582 => conv_std_logic_vector(173, 8),
46583 => conv_std_logic_vector(174, 8),
46584 => conv_std_logic_vector(175, 8),
46585 => conv_std_logic_vector(176, 8),
46586 => conv_std_logic_vector(176, 8),
46587 => conv_std_logic_vector(177, 8),
46588 => conv_std_logic_vector(178, 8),
46589 => conv_std_logic_vector(178, 8),
46590 => conv_std_logic_vector(179, 8),
46591 => conv_std_logic_vector(180, 8),
46592 => conv_std_logic_vector(0, 8),
46593 => conv_std_logic_vector(0, 8),
46594 => conv_std_logic_vector(1, 8),
46595 => conv_std_logic_vector(2, 8),
46596 => conv_std_logic_vector(2, 8),
46597 => conv_std_logic_vector(3, 8),
46598 => conv_std_logic_vector(4, 8),
46599 => conv_std_logic_vector(4, 8),
46600 => conv_std_logic_vector(5, 8),
46601 => conv_std_logic_vector(6, 8),
46602 => conv_std_logic_vector(7, 8),
46603 => conv_std_logic_vector(7, 8),
46604 => conv_std_logic_vector(8, 8),
46605 => conv_std_logic_vector(9, 8),
46606 => conv_std_logic_vector(9, 8),
46607 => conv_std_logic_vector(10, 8),
46608 => conv_std_logic_vector(11, 8),
46609 => conv_std_logic_vector(12, 8),
46610 => conv_std_logic_vector(12, 8),
46611 => conv_std_logic_vector(13, 8),
46612 => conv_std_logic_vector(14, 8),
46613 => conv_std_logic_vector(14, 8),
46614 => conv_std_logic_vector(15, 8),
46615 => conv_std_logic_vector(16, 8),
46616 => conv_std_logic_vector(17, 8),
46617 => conv_std_logic_vector(17, 8),
46618 => conv_std_logic_vector(18, 8),
46619 => conv_std_logic_vector(19, 8),
46620 => conv_std_logic_vector(19, 8),
46621 => conv_std_logic_vector(20, 8),
46622 => conv_std_logic_vector(21, 8),
46623 => conv_std_logic_vector(22, 8),
46624 => conv_std_logic_vector(22, 8),
46625 => conv_std_logic_vector(23, 8),
46626 => conv_std_logic_vector(24, 8),
46627 => conv_std_logic_vector(24, 8),
46628 => conv_std_logic_vector(25, 8),
46629 => conv_std_logic_vector(26, 8),
46630 => conv_std_logic_vector(27, 8),
46631 => conv_std_logic_vector(27, 8),
46632 => conv_std_logic_vector(28, 8),
46633 => conv_std_logic_vector(29, 8),
46634 => conv_std_logic_vector(29, 8),
46635 => conv_std_logic_vector(30, 8),
46636 => conv_std_logic_vector(31, 8),
46637 => conv_std_logic_vector(31, 8),
46638 => conv_std_logic_vector(32, 8),
46639 => conv_std_logic_vector(33, 8),
46640 => conv_std_logic_vector(34, 8),
46641 => conv_std_logic_vector(34, 8),
46642 => conv_std_logic_vector(35, 8),
46643 => conv_std_logic_vector(36, 8),
46644 => conv_std_logic_vector(36, 8),
46645 => conv_std_logic_vector(37, 8),
46646 => conv_std_logic_vector(38, 8),
46647 => conv_std_logic_vector(39, 8),
46648 => conv_std_logic_vector(39, 8),
46649 => conv_std_logic_vector(40, 8),
46650 => conv_std_logic_vector(41, 8),
46651 => conv_std_logic_vector(41, 8),
46652 => conv_std_logic_vector(42, 8),
46653 => conv_std_logic_vector(43, 8),
46654 => conv_std_logic_vector(44, 8),
46655 => conv_std_logic_vector(44, 8),
46656 => conv_std_logic_vector(45, 8),
46657 => conv_std_logic_vector(46, 8),
46658 => conv_std_logic_vector(46, 8),
46659 => conv_std_logic_vector(47, 8),
46660 => conv_std_logic_vector(48, 8),
46661 => conv_std_logic_vector(49, 8),
46662 => conv_std_logic_vector(49, 8),
46663 => conv_std_logic_vector(50, 8),
46664 => conv_std_logic_vector(51, 8),
46665 => conv_std_logic_vector(51, 8),
46666 => conv_std_logic_vector(52, 8),
46667 => conv_std_logic_vector(53, 8),
46668 => conv_std_logic_vector(54, 8),
46669 => conv_std_logic_vector(54, 8),
46670 => conv_std_logic_vector(55, 8),
46671 => conv_std_logic_vector(56, 8),
46672 => conv_std_logic_vector(56, 8),
46673 => conv_std_logic_vector(57, 8),
46674 => conv_std_logic_vector(58, 8),
46675 => conv_std_logic_vector(59, 8),
46676 => conv_std_logic_vector(59, 8),
46677 => conv_std_logic_vector(60, 8),
46678 => conv_std_logic_vector(61, 8),
46679 => conv_std_logic_vector(61, 8),
46680 => conv_std_logic_vector(62, 8),
46681 => conv_std_logic_vector(63, 8),
46682 => conv_std_logic_vector(63, 8),
46683 => conv_std_logic_vector(64, 8),
46684 => conv_std_logic_vector(65, 8),
46685 => conv_std_logic_vector(66, 8),
46686 => conv_std_logic_vector(66, 8),
46687 => conv_std_logic_vector(67, 8),
46688 => conv_std_logic_vector(68, 8),
46689 => conv_std_logic_vector(68, 8),
46690 => conv_std_logic_vector(69, 8),
46691 => conv_std_logic_vector(70, 8),
46692 => conv_std_logic_vector(71, 8),
46693 => conv_std_logic_vector(71, 8),
46694 => conv_std_logic_vector(72, 8),
46695 => conv_std_logic_vector(73, 8),
46696 => conv_std_logic_vector(73, 8),
46697 => conv_std_logic_vector(74, 8),
46698 => conv_std_logic_vector(75, 8),
46699 => conv_std_logic_vector(76, 8),
46700 => conv_std_logic_vector(76, 8),
46701 => conv_std_logic_vector(77, 8),
46702 => conv_std_logic_vector(78, 8),
46703 => conv_std_logic_vector(78, 8),
46704 => conv_std_logic_vector(79, 8),
46705 => conv_std_logic_vector(80, 8),
46706 => conv_std_logic_vector(81, 8),
46707 => conv_std_logic_vector(81, 8),
46708 => conv_std_logic_vector(82, 8),
46709 => conv_std_logic_vector(83, 8),
46710 => conv_std_logic_vector(83, 8),
46711 => conv_std_logic_vector(84, 8),
46712 => conv_std_logic_vector(85, 8),
46713 => conv_std_logic_vector(86, 8),
46714 => conv_std_logic_vector(86, 8),
46715 => conv_std_logic_vector(87, 8),
46716 => conv_std_logic_vector(88, 8),
46717 => conv_std_logic_vector(88, 8),
46718 => conv_std_logic_vector(89, 8),
46719 => conv_std_logic_vector(90, 8),
46720 => conv_std_logic_vector(91, 8),
46721 => conv_std_logic_vector(91, 8),
46722 => conv_std_logic_vector(92, 8),
46723 => conv_std_logic_vector(93, 8),
46724 => conv_std_logic_vector(93, 8),
46725 => conv_std_logic_vector(94, 8),
46726 => conv_std_logic_vector(95, 8),
46727 => conv_std_logic_vector(95, 8),
46728 => conv_std_logic_vector(96, 8),
46729 => conv_std_logic_vector(97, 8),
46730 => conv_std_logic_vector(98, 8),
46731 => conv_std_logic_vector(98, 8),
46732 => conv_std_logic_vector(99, 8),
46733 => conv_std_logic_vector(100, 8),
46734 => conv_std_logic_vector(100, 8),
46735 => conv_std_logic_vector(101, 8),
46736 => conv_std_logic_vector(102, 8),
46737 => conv_std_logic_vector(103, 8),
46738 => conv_std_logic_vector(103, 8),
46739 => conv_std_logic_vector(104, 8),
46740 => conv_std_logic_vector(105, 8),
46741 => conv_std_logic_vector(105, 8),
46742 => conv_std_logic_vector(106, 8),
46743 => conv_std_logic_vector(107, 8),
46744 => conv_std_logic_vector(108, 8),
46745 => conv_std_logic_vector(108, 8),
46746 => conv_std_logic_vector(109, 8),
46747 => conv_std_logic_vector(110, 8),
46748 => conv_std_logic_vector(110, 8),
46749 => conv_std_logic_vector(111, 8),
46750 => conv_std_logic_vector(112, 8),
46751 => conv_std_logic_vector(113, 8),
46752 => conv_std_logic_vector(113, 8),
46753 => conv_std_logic_vector(114, 8),
46754 => conv_std_logic_vector(115, 8),
46755 => conv_std_logic_vector(115, 8),
46756 => conv_std_logic_vector(116, 8),
46757 => conv_std_logic_vector(117, 8),
46758 => conv_std_logic_vector(118, 8),
46759 => conv_std_logic_vector(118, 8),
46760 => conv_std_logic_vector(119, 8),
46761 => conv_std_logic_vector(120, 8),
46762 => conv_std_logic_vector(120, 8),
46763 => conv_std_logic_vector(121, 8),
46764 => conv_std_logic_vector(122, 8),
46765 => conv_std_logic_vector(122, 8),
46766 => conv_std_logic_vector(123, 8),
46767 => conv_std_logic_vector(124, 8),
46768 => conv_std_logic_vector(125, 8),
46769 => conv_std_logic_vector(125, 8),
46770 => conv_std_logic_vector(126, 8),
46771 => conv_std_logic_vector(127, 8),
46772 => conv_std_logic_vector(127, 8),
46773 => conv_std_logic_vector(128, 8),
46774 => conv_std_logic_vector(129, 8),
46775 => conv_std_logic_vector(130, 8),
46776 => conv_std_logic_vector(130, 8),
46777 => conv_std_logic_vector(131, 8),
46778 => conv_std_logic_vector(132, 8),
46779 => conv_std_logic_vector(132, 8),
46780 => conv_std_logic_vector(133, 8),
46781 => conv_std_logic_vector(134, 8),
46782 => conv_std_logic_vector(135, 8),
46783 => conv_std_logic_vector(135, 8),
46784 => conv_std_logic_vector(136, 8),
46785 => conv_std_logic_vector(137, 8),
46786 => conv_std_logic_vector(137, 8),
46787 => conv_std_logic_vector(138, 8),
46788 => conv_std_logic_vector(139, 8),
46789 => conv_std_logic_vector(140, 8),
46790 => conv_std_logic_vector(140, 8),
46791 => conv_std_logic_vector(141, 8),
46792 => conv_std_logic_vector(142, 8),
46793 => conv_std_logic_vector(142, 8),
46794 => conv_std_logic_vector(143, 8),
46795 => conv_std_logic_vector(144, 8),
46796 => conv_std_logic_vector(145, 8),
46797 => conv_std_logic_vector(145, 8),
46798 => conv_std_logic_vector(146, 8),
46799 => conv_std_logic_vector(147, 8),
46800 => conv_std_logic_vector(147, 8),
46801 => conv_std_logic_vector(148, 8),
46802 => conv_std_logic_vector(149, 8),
46803 => conv_std_logic_vector(150, 8),
46804 => conv_std_logic_vector(150, 8),
46805 => conv_std_logic_vector(151, 8),
46806 => conv_std_logic_vector(152, 8),
46807 => conv_std_logic_vector(152, 8),
46808 => conv_std_logic_vector(153, 8),
46809 => conv_std_logic_vector(154, 8),
46810 => conv_std_logic_vector(154, 8),
46811 => conv_std_logic_vector(155, 8),
46812 => conv_std_logic_vector(156, 8),
46813 => conv_std_logic_vector(157, 8),
46814 => conv_std_logic_vector(157, 8),
46815 => conv_std_logic_vector(158, 8),
46816 => conv_std_logic_vector(159, 8),
46817 => conv_std_logic_vector(159, 8),
46818 => conv_std_logic_vector(160, 8),
46819 => conv_std_logic_vector(161, 8),
46820 => conv_std_logic_vector(162, 8),
46821 => conv_std_logic_vector(162, 8),
46822 => conv_std_logic_vector(163, 8),
46823 => conv_std_logic_vector(164, 8),
46824 => conv_std_logic_vector(164, 8),
46825 => conv_std_logic_vector(165, 8),
46826 => conv_std_logic_vector(166, 8),
46827 => conv_std_logic_vector(167, 8),
46828 => conv_std_logic_vector(167, 8),
46829 => conv_std_logic_vector(168, 8),
46830 => conv_std_logic_vector(169, 8),
46831 => conv_std_logic_vector(169, 8),
46832 => conv_std_logic_vector(170, 8),
46833 => conv_std_logic_vector(171, 8),
46834 => conv_std_logic_vector(172, 8),
46835 => conv_std_logic_vector(172, 8),
46836 => conv_std_logic_vector(173, 8),
46837 => conv_std_logic_vector(174, 8),
46838 => conv_std_logic_vector(174, 8),
46839 => conv_std_logic_vector(175, 8),
46840 => conv_std_logic_vector(176, 8),
46841 => conv_std_logic_vector(177, 8),
46842 => conv_std_logic_vector(177, 8),
46843 => conv_std_logic_vector(178, 8),
46844 => conv_std_logic_vector(179, 8),
46845 => conv_std_logic_vector(179, 8),
46846 => conv_std_logic_vector(180, 8),
46847 => conv_std_logic_vector(181, 8),
46848 => conv_std_logic_vector(0, 8),
46849 => conv_std_logic_vector(0, 8),
46850 => conv_std_logic_vector(1, 8),
46851 => conv_std_logic_vector(2, 8),
46852 => conv_std_logic_vector(2, 8),
46853 => conv_std_logic_vector(3, 8),
46854 => conv_std_logic_vector(4, 8),
46855 => conv_std_logic_vector(5, 8),
46856 => conv_std_logic_vector(5, 8),
46857 => conv_std_logic_vector(6, 8),
46858 => conv_std_logic_vector(7, 8),
46859 => conv_std_logic_vector(7, 8),
46860 => conv_std_logic_vector(8, 8),
46861 => conv_std_logic_vector(9, 8),
46862 => conv_std_logic_vector(10, 8),
46863 => conv_std_logic_vector(10, 8),
46864 => conv_std_logic_vector(11, 8),
46865 => conv_std_logic_vector(12, 8),
46866 => conv_std_logic_vector(12, 8),
46867 => conv_std_logic_vector(13, 8),
46868 => conv_std_logic_vector(14, 8),
46869 => conv_std_logic_vector(15, 8),
46870 => conv_std_logic_vector(15, 8),
46871 => conv_std_logic_vector(16, 8),
46872 => conv_std_logic_vector(17, 8),
46873 => conv_std_logic_vector(17, 8),
46874 => conv_std_logic_vector(18, 8),
46875 => conv_std_logic_vector(19, 8),
46876 => conv_std_logic_vector(20, 8),
46877 => conv_std_logic_vector(20, 8),
46878 => conv_std_logic_vector(21, 8),
46879 => conv_std_logic_vector(22, 8),
46880 => conv_std_logic_vector(22, 8),
46881 => conv_std_logic_vector(23, 8),
46882 => conv_std_logic_vector(24, 8),
46883 => conv_std_logic_vector(25, 8),
46884 => conv_std_logic_vector(25, 8),
46885 => conv_std_logic_vector(26, 8),
46886 => conv_std_logic_vector(27, 8),
46887 => conv_std_logic_vector(27, 8),
46888 => conv_std_logic_vector(28, 8),
46889 => conv_std_logic_vector(29, 8),
46890 => conv_std_logic_vector(30, 8),
46891 => conv_std_logic_vector(30, 8),
46892 => conv_std_logic_vector(31, 8),
46893 => conv_std_logic_vector(32, 8),
46894 => conv_std_logic_vector(32, 8),
46895 => conv_std_logic_vector(33, 8),
46896 => conv_std_logic_vector(34, 8),
46897 => conv_std_logic_vector(35, 8),
46898 => conv_std_logic_vector(35, 8),
46899 => conv_std_logic_vector(36, 8),
46900 => conv_std_logic_vector(37, 8),
46901 => conv_std_logic_vector(37, 8),
46902 => conv_std_logic_vector(38, 8),
46903 => conv_std_logic_vector(39, 8),
46904 => conv_std_logic_vector(40, 8),
46905 => conv_std_logic_vector(40, 8),
46906 => conv_std_logic_vector(41, 8),
46907 => conv_std_logic_vector(42, 8),
46908 => conv_std_logic_vector(42, 8),
46909 => conv_std_logic_vector(43, 8),
46910 => conv_std_logic_vector(44, 8),
46911 => conv_std_logic_vector(45, 8),
46912 => conv_std_logic_vector(45, 8),
46913 => conv_std_logic_vector(46, 8),
46914 => conv_std_logic_vector(47, 8),
46915 => conv_std_logic_vector(47, 8),
46916 => conv_std_logic_vector(48, 8),
46917 => conv_std_logic_vector(49, 8),
46918 => conv_std_logic_vector(50, 8),
46919 => conv_std_logic_vector(50, 8),
46920 => conv_std_logic_vector(51, 8),
46921 => conv_std_logic_vector(52, 8),
46922 => conv_std_logic_vector(52, 8),
46923 => conv_std_logic_vector(53, 8),
46924 => conv_std_logic_vector(54, 8),
46925 => conv_std_logic_vector(55, 8),
46926 => conv_std_logic_vector(55, 8),
46927 => conv_std_logic_vector(56, 8),
46928 => conv_std_logic_vector(57, 8),
46929 => conv_std_logic_vector(57, 8),
46930 => conv_std_logic_vector(58, 8),
46931 => conv_std_logic_vector(59, 8),
46932 => conv_std_logic_vector(60, 8),
46933 => conv_std_logic_vector(60, 8),
46934 => conv_std_logic_vector(61, 8),
46935 => conv_std_logic_vector(62, 8),
46936 => conv_std_logic_vector(62, 8),
46937 => conv_std_logic_vector(63, 8),
46938 => conv_std_logic_vector(64, 8),
46939 => conv_std_logic_vector(65, 8),
46940 => conv_std_logic_vector(65, 8),
46941 => conv_std_logic_vector(66, 8),
46942 => conv_std_logic_vector(67, 8),
46943 => conv_std_logic_vector(67, 8),
46944 => conv_std_logic_vector(68, 8),
46945 => conv_std_logic_vector(69, 8),
46946 => conv_std_logic_vector(70, 8),
46947 => conv_std_logic_vector(70, 8),
46948 => conv_std_logic_vector(71, 8),
46949 => conv_std_logic_vector(72, 8),
46950 => conv_std_logic_vector(72, 8),
46951 => conv_std_logic_vector(73, 8),
46952 => conv_std_logic_vector(74, 8),
46953 => conv_std_logic_vector(75, 8),
46954 => conv_std_logic_vector(75, 8),
46955 => conv_std_logic_vector(76, 8),
46956 => conv_std_logic_vector(77, 8),
46957 => conv_std_logic_vector(77, 8),
46958 => conv_std_logic_vector(78, 8),
46959 => conv_std_logic_vector(79, 8),
46960 => conv_std_logic_vector(80, 8),
46961 => conv_std_logic_vector(80, 8),
46962 => conv_std_logic_vector(81, 8),
46963 => conv_std_logic_vector(82, 8),
46964 => conv_std_logic_vector(82, 8),
46965 => conv_std_logic_vector(83, 8),
46966 => conv_std_logic_vector(84, 8),
46967 => conv_std_logic_vector(85, 8),
46968 => conv_std_logic_vector(85, 8),
46969 => conv_std_logic_vector(86, 8),
46970 => conv_std_logic_vector(87, 8),
46971 => conv_std_logic_vector(87, 8),
46972 => conv_std_logic_vector(88, 8),
46973 => conv_std_logic_vector(89, 8),
46974 => conv_std_logic_vector(90, 8),
46975 => conv_std_logic_vector(90, 8),
46976 => conv_std_logic_vector(91, 8),
46977 => conv_std_logic_vector(92, 8),
46978 => conv_std_logic_vector(92, 8),
46979 => conv_std_logic_vector(93, 8),
46980 => conv_std_logic_vector(94, 8),
46981 => conv_std_logic_vector(95, 8),
46982 => conv_std_logic_vector(95, 8),
46983 => conv_std_logic_vector(96, 8),
46984 => conv_std_logic_vector(97, 8),
46985 => conv_std_logic_vector(97, 8),
46986 => conv_std_logic_vector(98, 8),
46987 => conv_std_logic_vector(99, 8),
46988 => conv_std_logic_vector(100, 8),
46989 => conv_std_logic_vector(100, 8),
46990 => conv_std_logic_vector(101, 8),
46991 => conv_std_logic_vector(102, 8),
46992 => conv_std_logic_vector(102, 8),
46993 => conv_std_logic_vector(103, 8),
46994 => conv_std_logic_vector(104, 8),
46995 => conv_std_logic_vector(105, 8),
46996 => conv_std_logic_vector(105, 8),
46997 => conv_std_logic_vector(106, 8),
46998 => conv_std_logic_vector(107, 8),
46999 => conv_std_logic_vector(107, 8),
47000 => conv_std_logic_vector(108, 8),
47001 => conv_std_logic_vector(109, 8),
47002 => conv_std_logic_vector(110, 8),
47003 => conv_std_logic_vector(110, 8),
47004 => conv_std_logic_vector(111, 8),
47005 => conv_std_logic_vector(112, 8),
47006 => conv_std_logic_vector(112, 8),
47007 => conv_std_logic_vector(113, 8),
47008 => conv_std_logic_vector(114, 8),
47009 => conv_std_logic_vector(115, 8),
47010 => conv_std_logic_vector(115, 8),
47011 => conv_std_logic_vector(116, 8),
47012 => conv_std_logic_vector(117, 8),
47013 => conv_std_logic_vector(117, 8),
47014 => conv_std_logic_vector(118, 8),
47015 => conv_std_logic_vector(119, 8),
47016 => conv_std_logic_vector(120, 8),
47017 => conv_std_logic_vector(120, 8),
47018 => conv_std_logic_vector(121, 8),
47019 => conv_std_logic_vector(122, 8),
47020 => conv_std_logic_vector(122, 8),
47021 => conv_std_logic_vector(123, 8),
47022 => conv_std_logic_vector(124, 8),
47023 => conv_std_logic_vector(125, 8),
47024 => conv_std_logic_vector(125, 8),
47025 => conv_std_logic_vector(126, 8),
47026 => conv_std_logic_vector(127, 8),
47027 => conv_std_logic_vector(127, 8),
47028 => conv_std_logic_vector(128, 8),
47029 => conv_std_logic_vector(129, 8),
47030 => conv_std_logic_vector(130, 8),
47031 => conv_std_logic_vector(130, 8),
47032 => conv_std_logic_vector(131, 8),
47033 => conv_std_logic_vector(132, 8),
47034 => conv_std_logic_vector(132, 8),
47035 => conv_std_logic_vector(133, 8),
47036 => conv_std_logic_vector(134, 8),
47037 => conv_std_logic_vector(135, 8),
47038 => conv_std_logic_vector(135, 8),
47039 => conv_std_logic_vector(136, 8),
47040 => conv_std_logic_vector(137, 8),
47041 => conv_std_logic_vector(137, 8),
47042 => conv_std_logic_vector(138, 8),
47043 => conv_std_logic_vector(139, 8),
47044 => conv_std_logic_vector(140, 8),
47045 => conv_std_logic_vector(140, 8),
47046 => conv_std_logic_vector(141, 8),
47047 => conv_std_logic_vector(142, 8),
47048 => conv_std_logic_vector(142, 8),
47049 => conv_std_logic_vector(143, 8),
47050 => conv_std_logic_vector(144, 8),
47051 => conv_std_logic_vector(145, 8),
47052 => conv_std_logic_vector(145, 8),
47053 => conv_std_logic_vector(146, 8),
47054 => conv_std_logic_vector(147, 8),
47055 => conv_std_logic_vector(147, 8),
47056 => conv_std_logic_vector(148, 8),
47057 => conv_std_logic_vector(149, 8),
47058 => conv_std_logic_vector(150, 8),
47059 => conv_std_logic_vector(150, 8),
47060 => conv_std_logic_vector(151, 8),
47061 => conv_std_logic_vector(152, 8),
47062 => conv_std_logic_vector(152, 8),
47063 => conv_std_logic_vector(153, 8),
47064 => conv_std_logic_vector(154, 8),
47065 => conv_std_logic_vector(155, 8),
47066 => conv_std_logic_vector(155, 8),
47067 => conv_std_logic_vector(156, 8),
47068 => conv_std_logic_vector(157, 8),
47069 => conv_std_logic_vector(157, 8),
47070 => conv_std_logic_vector(158, 8),
47071 => conv_std_logic_vector(159, 8),
47072 => conv_std_logic_vector(160, 8),
47073 => conv_std_logic_vector(160, 8),
47074 => conv_std_logic_vector(161, 8),
47075 => conv_std_logic_vector(162, 8),
47076 => conv_std_logic_vector(162, 8),
47077 => conv_std_logic_vector(163, 8),
47078 => conv_std_logic_vector(164, 8),
47079 => conv_std_logic_vector(165, 8),
47080 => conv_std_logic_vector(165, 8),
47081 => conv_std_logic_vector(166, 8),
47082 => conv_std_logic_vector(167, 8),
47083 => conv_std_logic_vector(167, 8),
47084 => conv_std_logic_vector(168, 8),
47085 => conv_std_logic_vector(169, 8),
47086 => conv_std_logic_vector(170, 8),
47087 => conv_std_logic_vector(170, 8),
47088 => conv_std_logic_vector(171, 8),
47089 => conv_std_logic_vector(172, 8),
47090 => conv_std_logic_vector(172, 8),
47091 => conv_std_logic_vector(173, 8),
47092 => conv_std_logic_vector(174, 8),
47093 => conv_std_logic_vector(175, 8),
47094 => conv_std_logic_vector(175, 8),
47095 => conv_std_logic_vector(176, 8),
47096 => conv_std_logic_vector(177, 8),
47097 => conv_std_logic_vector(177, 8),
47098 => conv_std_logic_vector(178, 8),
47099 => conv_std_logic_vector(179, 8),
47100 => conv_std_logic_vector(180, 8),
47101 => conv_std_logic_vector(180, 8),
47102 => conv_std_logic_vector(181, 8),
47103 => conv_std_logic_vector(182, 8),
47104 => conv_std_logic_vector(0, 8),
47105 => conv_std_logic_vector(0, 8),
47106 => conv_std_logic_vector(1, 8),
47107 => conv_std_logic_vector(2, 8),
47108 => conv_std_logic_vector(2, 8),
47109 => conv_std_logic_vector(3, 8),
47110 => conv_std_logic_vector(4, 8),
47111 => conv_std_logic_vector(5, 8),
47112 => conv_std_logic_vector(5, 8),
47113 => conv_std_logic_vector(6, 8),
47114 => conv_std_logic_vector(7, 8),
47115 => conv_std_logic_vector(7, 8),
47116 => conv_std_logic_vector(8, 8),
47117 => conv_std_logic_vector(9, 8),
47118 => conv_std_logic_vector(10, 8),
47119 => conv_std_logic_vector(10, 8),
47120 => conv_std_logic_vector(11, 8),
47121 => conv_std_logic_vector(12, 8),
47122 => conv_std_logic_vector(12, 8),
47123 => conv_std_logic_vector(13, 8),
47124 => conv_std_logic_vector(14, 8),
47125 => conv_std_logic_vector(15, 8),
47126 => conv_std_logic_vector(15, 8),
47127 => conv_std_logic_vector(16, 8),
47128 => conv_std_logic_vector(17, 8),
47129 => conv_std_logic_vector(17, 8),
47130 => conv_std_logic_vector(18, 8),
47131 => conv_std_logic_vector(19, 8),
47132 => conv_std_logic_vector(20, 8),
47133 => conv_std_logic_vector(20, 8),
47134 => conv_std_logic_vector(21, 8),
47135 => conv_std_logic_vector(22, 8),
47136 => conv_std_logic_vector(23, 8),
47137 => conv_std_logic_vector(23, 8),
47138 => conv_std_logic_vector(24, 8),
47139 => conv_std_logic_vector(25, 8),
47140 => conv_std_logic_vector(25, 8),
47141 => conv_std_logic_vector(26, 8),
47142 => conv_std_logic_vector(27, 8),
47143 => conv_std_logic_vector(28, 8),
47144 => conv_std_logic_vector(28, 8),
47145 => conv_std_logic_vector(29, 8),
47146 => conv_std_logic_vector(30, 8),
47147 => conv_std_logic_vector(30, 8),
47148 => conv_std_logic_vector(31, 8),
47149 => conv_std_logic_vector(32, 8),
47150 => conv_std_logic_vector(33, 8),
47151 => conv_std_logic_vector(33, 8),
47152 => conv_std_logic_vector(34, 8),
47153 => conv_std_logic_vector(35, 8),
47154 => conv_std_logic_vector(35, 8),
47155 => conv_std_logic_vector(36, 8),
47156 => conv_std_logic_vector(37, 8),
47157 => conv_std_logic_vector(38, 8),
47158 => conv_std_logic_vector(38, 8),
47159 => conv_std_logic_vector(39, 8),
47160 => conv_std_logic_vector(40, 8),
47161 => conv_std_logic_vector(40, 8),
47162 => conv_std_logic_vector(41, 8),
47163 => conv_std_logic_vector(42, 8),
47164 => conv_std_logic_vector(43, 8),
47165 => conv_std_logic_vector(43, 8),
47166 => conv_std_logic_vector(44, 8),
47167 => conv_std_logic_vector(45, 8),
47168 => conv_std_logic_vector(46, 8),
47169 => conv_std_logic_vector(46, 8),
47170 => conv_std_logic_vector(47, 8),
47171 => conv_std_logic_vector(48, 8),
47172 => conv_std_logic_vector(48, 8),
47173 => conv_std_logic_vector(49, 8),
47174 => conv_std_logic_vector(50, 8),
47175 => conv_std_logic_vector(51, 8),
47176 => conv_std_logic_vector(51, 8),
47177 => conv_std_logic_vector(52, 8),
47178 => conv_std_logic_vector(53, 8),
47179 => conv_std_logic_vector(53, 8),
47180 => conv_std_logic_vector(54, 8),
47181 => conv_std_logic_vector(55, 8),
47182 => conv_std_logic_vector(56, 8),
47183 => conv_std_logic_vector(56, 8),
47184 => conv_std_logic_vector(57, 8),
47185 => conv_std_logic_vector(58, 8),
47186 => conv_std_logic_vector(58, 8),
47187 => conv_std_logic_vector(59, 8),
47188 => conv_std_logic_vector(60, 8),
47189 => conv_std_logic_vector(61, 8),
47190 => conv_std_logic_vector(61, 8),
47191 => conv_std_logic_vector(62, 8),
47192 => conv_std_logic_vector(63, 8),
47193 => conv_std_logic_vector(63, 8),
47194 => conv_std_logic_vector(64, 8),
47195 => conv_std_logic_vector(65, 8),
47196 => conv_std_logic_vector(66, 8),
47197 => conv_std_logic_vector(66, 8),
47198 => conv_std_logic_vector(67, 8),
47199 => conv_std_logic_vector(68, 8),
47200 => conv_std_logic_vector(69, 8),
47201 => conv_std_logic_vector(69, 8),
47202 => conv_std_logic_vector(70, 8),
47203 => conv_std_logic_vector(71, 8),
47204 => conv_std_logic_vector(71, 8),
47205 => conv_std_logic_vector(72, 8),
47206 => conv_std_logic_vector(73, 8),
47207 => conv_std_logic_vector(74, 8),
47208 => conv_std_logic_vector(74, 8),
47209 => conv_std_logic_vector(75, 8),
47210 => conv_std_logic_vector(76, 8),
47211 => conv_std_logic_vector(76, 8),
47212 => conv_std_logic_vector(77, 8),
47213 => conv_std_logic_vector(78, 8),
47214 => conv_std_logic_vector(79, 8),
47215 => conv_std_logic_vector(79, 8),
47216 => conv_std_logic_vector(80, 8),
47217 => conv_std_logic_vector(81, 8),
47218 => conv_std_logic_vector(81, 8),
47219 => conv_std_logic_vector(82, 8),
47220 => conv_std_logic_vector(83, 8),
47221 => conv_std_logic_vector(84, 8),
47222 => conv_std_logic_vector(84, 8),
47223 => conv_std_logic_vector(85, 8),
47224 => conv_std_logic_vector(86, 8),
47225 => conv_std_logic_vector(86, 8),
47226 => conv_std_logic_vector(87, 8),
47227 => conv_std_logic_vector(88, 8),
47228 => conv_std_logic_vector(89, 8),
47229 => conv_std_logic_vector(89, 8),
47230 => conv_std_logic_vector(90, 8),
47231 => conv_std_logic_vector(91, 8),
47232 => conv_std_logic_vector(92, 8),
47233 => conv_std_logic_vector(92, 8),
47234 => conv_std_logic_vector(93, 8),
47235 => conv_std_logic_vector(94, 8),
47236 => conv_std_logic_vector(94, 8),
47237 => conv_std_logic_vector(95, 8),
47238 => conv_std_logic_vector(96, 8),
47239 => conv_std_logic_vector(97, 8),
47240 => conv_std_logic_vector(97, 8),
47241 => conv_std_logic_vector(98, 8),
47242 => conv_std_logic_vector(99, 8),
47243 => conv_std_logic_vector(99, 8),
47244 => conv_std_logic_vector(100, 8),
47245 => conv_std_logic_vector(101, 8),
47246 => conv_std_logic_vector(102, 8),
47247 => conv_std_logic_vector(102, 8),
47248 => conv_std_logic_vector(103, 8),
47249 => conv_std_logic_vector(104, 8),
47250 => conv_std_logic_vector(104, 8),
47251 => conv_std_logic_vector(105, 8),
47252 => conv_std_logic_vector(106, 8),
47253 => conv_std_logic_vector(107, 8),
47254 => conv_std_logic_vector(107, 8),
47255 => conv_std_logic_vector(108, 8),
47256 => conv_std_logic_vector(109, 8),
47257 => conv_std_logic_vector(109, 8),
47258 => conv_std_logic_vector(110, 8),
47259 => conv_std_logic_vector(111, 8),
47260 => conv_std_logic_vector(112, 8),
47261 => conv_std_logic_vector(112, 8),
47262 => conv_std_logic_vector(113, 8),
47263 => conv_std_logic_vector(114, 8),
47264 => conv_std_logic_vector(115, 8),
47265 => conv_std_logic_vector(115, 8),
47266 => conv_std_logic_vector(116, 8),
47267 => conv_std_logic_vector(117, 8),
47268 => conv_std_logic_vector(117, 8),
47269 => conv_std_logic_vector(118, 8),
47270 => conv_std_logic_vector(119, 8),
47271 => conv_std_logic_vector(120, 8),
47272 => conv_std_logic_vector(120, 8),
47273 => conv_std_logic_vector(121, 8),
47274 => conv_std_logic_vector(122, 8),
47275 => conv_std_logic_vector(122, 8),
47276 => conv_std_logic_vector(123, 8),
47277 => conv_std_logic_vector(124, 8),
47278 => conv_std_logic_vector(125, 8),
47279 => conv_std_logic_vector(125, 8),
47280 => conv_std_logic_vector(126, 8),
47281 => conv_std_logic_vector(127, 8),
47282 => conv_std_logic_vector(127, 8),
47283 => conv_std_logic_vector(128, 8),
47284 => conv_std_logic_vector(129, 8),
47285 => conv_std_logic_vector(130, 8),
47286 => conv_std_logic_vector(130, 8),
47287 => conv_std_logic_vector(131, 8),
47288 => conv_std_logic_vector(132, 8),
47289 => conv_std_logic_vector(132, 8),
47290 => conv_std_logic_vector(133, 8),
47291 => conv_std_logic_vector(134, 8),
47292 => conv_std_logic_vector(135, 8),
47293 => conv_std_logic_vector(135, 8),
47294 => conv_std_logic_vector(136, 8),
47295 => conv_std_logic_vector(137, 8),
47296 => conv_std_logic_vector(138, 8),
47297 => conv_std_logic_vector(138, 8),
47298 => conv_std_logic_vector(139, 8),
47299 => conv_std_logic_vector(140, 8),
47300 => conv_std_logic_vector(140, 8),
47301 => conv_std_logic_vector(141, 8),
47302 => conv_std_logic_vector(142, 8),
47303 => conv_std_logic_vector(143, 8),
47304 => conv_std_logic_vector(143, 8),
47305 => conv_std_logic_vector(144, 8),
47306 => conv_std_logic_vector(145, 8),
47307 => conv_std_logic_vector(145, 8),
47308 => conv_std_logic_vector(146, 8),
47309 => conv_std_logic_vector(147, 8),
47310 => conv_std_logic_vector(148, 8),
47311 => conv_std_logic_vector(148, 8),
47312 => conv_std_logic_vector(149, 8),
47313 => conv_std_logic_vector(150, 8),
47314 => conv_std_logic_vector(150, 8),
47315 => conv_std_logic_vector(151, 8),
47316 => conv_std_logic_vector(152, 8),
47317 => conv_std_logic_vector(153, 8),
47318 => conv_std_logic_vector(153, 8),
47319 => conv_std_logic_vector(154, 8),
47320 => conv_std_logic_vector(155, 8),
47321 => conv_std_logic_vector(155, 8),
47322 => conv_std_logic_vector(156, 8),
47323 => conv_std_logic_vector(157, 8),
47324 => conv_std_logic_vector(158, 8),
47325 => conv_std_logic_vector(158, 8),
47326 => conv_std_logic_vector(159, 8),
47327 => conv_std_logic_vector(160, 8),
47328 => conv_std_logic_vector(161, 8),
47329 => conv_std_logic_vector(161, 8),
47330 => conv_std_logic_vector(162, 8),
47331 => conv_std_logic_vector(163, 8),
47332 => conv_std_logic_vector(163, 8),
47333 => conv_std_logic_vector(164, 8),
47334 => conv_std_logic_vector(165, 8),
47335 => conv_std_logic_vector(166, 8),
47336 => conv_std_logic_vector(166, 8),
47337 => conv_std_logic_vector(167, 8),
47338 => conv_std_logic_vector(168, 8),
47339 => conv_std_logic_vector(168, 8),
47340 => conv_std_logic_vector(169, 8),
47341 => conv_std_logic_vector(170, 8),
47342 => conv_std_logic_vector(171, 8),
47343 => conv_std_logic_vector(171, 8),
47344 => conv_std_logic_vector(172, 8),
47345 => conv_std_logic_vector(173, 8),
47346 => conv_std_logic_vector(173, 8),
47347 => conv_std_logic_vector(174, 8),
47348 => conv_std_logic_vector(175, 8),
47349 => conv_std_logic_vector(176, 8),
47350 => conv_std_logic_vector(176, 8),
47351 => conv_std_logic_vector(177, 8),
47352 => conv_std_logic_vector(178, 8),
47353 => conv_std_logic_vector(178, 8),
47354 => conv_std_logic_vector(179, 8),
47355 => conv_std_logic_vector(180, 8),
47356 => conv_std_logic_vector(181, 8),
47357 => conv_std_logic_vector(181, 8),
47358 => conv_std_logic_vector(182, 8),
47359 => conv_std_logic_vector(183, 8),
47360 => conv_std_logic_vector(0, 8),
47361 => conv_std_logic_vector(0, 8),
47362 => conv_std_logic_vector(1, 8),
47363 => conv_std_logic_vector(2, 8),
47364 => conv_std_logic_vector(2, 8),
47365 => conv_std_logic_vector(3, 8),
47366 => conv_std_logic_vector(4, 8),
47367 => conv_std_logic_vector(5, 8),
47368 => conv_std_logic_vector(5, 8),
47369 => conv_std_logic_vector(6, 8),
47370 => conv_std_logic_vector(7, 8),
47371 => conv_std_logic_vector(7, 8),
47372 => conv_std_logic_vector(8, 8),
47373 => conv_std_logic_vector(9, 8),
47374 => conv_std_logic_vector(10, 8),
47375 => conv_std_logic_vector(10, 8),
47376 => conv_std_logic_vector(11, 8),
47377 => conv_std_logic_vector(12, 8),
47378 => conv_std_logic_vector(13, 8),
47379 => conv_std_logic_vector(13, 8),
47380 => conv_std_logic_vector(14, 8),
47381 => conv_std_logic_vector(15, 8),
47382 => conv_std_logic_vector(15, 8),
47383 => conv_std_logic_vector(16, 8),
47384 => conv_std_logic_vector(17, 8),
47385 => conv_std_logic_vector(18, 8),
47386 => conv_std_logic_vector(18, 8),
47387 => conv_std_logic_vector(19, 8),
47388 => conv_std_logic_vector(20, 8),
47389 => conv_std_logic_vector(20, 8),
47390 => conv_std_logic_vector(21, 8),
47391 => conv_std_logic_vector(22, 8),
47392 => conv_std_logic_vector(23, 8),
47393 => conv_std_logic_vector(23, 8),
47394 => conv_std_logic_vector(24, 8),
47395 => conv_std_logic_vector(25, 8),
47396 => conv_std_logic_vector(26, 8),
47397 => conv_std_logic_vector(26, 8),
47398 => conv_std_logic_vector(27, 8),
47399 => conv_std_logic_vector(28, 8),
47400 => conv_std_logic_vector(28, 8),
47401 => conv_std_logic_vector(29, 8),
47402 => conv_std_logic_vector(30, 8),
47403 => conv_std_logic_vector(31, 8),
47404 => conv_std_logic_vector(31, 8),
47405 => conv_std_logic_vector(32, 8),
47406 => conv_std_logic_vector(33, 8),
47407 => conv_std_logic_vector(33, 8),
47408 => conv_std_logic_vector(34, 8),
47409 => conv_std_logic_vector(35, 8),
47410 => conv_std_logic_vector(36, 8),
47411 => conv_std_logic_vector(36, 8),
47412 => conv_std_logic_vector(37, 8),
47413 => conv_std_logic_vector(38, 8),
47414 => conv_std_logic_vector(39, 8),
47415 => conv_std_logic_vector(39, 8),
47416 => conv_std_logic_vector(40, 8),
47417 => conv_std_logic_vector(41, 8),
47418 => conv_std_logic_vector(41, 8),
47419 => conv_std_logic_vector(42, 8),
47420 => conv_std_logic_vector(43, 8),
47421 => conv_std_logic_vector(44, 8),
47422 => conv_std_logic_vector(44, 8),
47423 => conv_std_logic_vector(45, 8),
47424 => conv_std_logic_vector(46, 8),
47425 => conv_std_logic_vector(46, 8),
47426 => conv_std_logic_vector(47, 8),
47427 => conv_std_logic_vector(48, 8),
47428 => conv_std_logic_vector(49, 8),
47429 => conv_std_logic_vector(49, 8),
47430 => conv_std_logic_vector(50, 8),
47431 => conv_std_logic_vector(51, 8),
47432 => conv_std_logic_vector(52, 8),
47433 => conv_std_logic_vector(52, 8),
47434 => conv_std_logic_vector(53, 8),
47435 => conv_std_logic_vector(54, 8),
47436 => conv_std_logic_vector(54, 8),
47437 => conv_std_logic_vector(55, 8),
47438 => conv_std_logic_vector(56, 8),
47439 => conv_std_logic_vector(57, 8),
47440 => conv_std_logic_vector(57, 8),
47441 => conv_std_logic_vector(58, 8),
47442 => conv_std_logic_vector(59, 8),
47443 => conv_std_logic_vector(59, 8),
47444 => conv_std_logic_vector(60, 8),
47445 => conv_std_logic_vector(61, 8),
47446 => conv_std_logic_vector(62, 8),
47447 => conv_std_logic_vector(62, 8),
47448 => conv_std_logic_vector(63, 8),
47449 => conv_std_logic_vector(64, 8),
47450 => conv_std_logic_vector(65, 8),
47451 => conv_std_logic_vector(65, 8),
47452 => conv_std_logic_vector(66, 8),
47453 => conv_std_logic_vector(67, 8),
47454 => conv_std_logic_vector(67, 8),
47455 => conv_std_logic_vector(68, 8),
47456 => conv_std_logic_vector(69, 8),
47457 => conv_std_logic_vector(70, 8),
47458 => conv_std_logic_vector(70, 8),
47459 => conv_std_logic_vector(71, 8),
47460 => conv_std_logic_vector(72, 8),
47461 => conv_std_logic_vector(72, 8),
47462 => conv_std_logic_vector(73, 8),
47463 => conv_std_logic_vector(74, 8),
47464 => conv_std_logic_vector(75, 8),
47465 => conv_std_logic_vector(75, 8),
47466 => conv_std_logic_vector(76, 8),
47467 => conv_std_logic_vector(77, 8),
47468 => conv_std_logic_vector(78, 8),
47469 => conv_std_logic_vector(78, 8),
47470 => conv_std_logic_vector(79, 8),
47471 => conv_std_logic_vector(80, 8),
47472 => conv_std_logic_vector(80, 8),
47473 => conv_std_logic_vector(81, 8),
47474 => conv_std_logic_vector(82, 8),
47475 => conv_std_logic_vector(83, 8),
47476 => conv_std_logic_vector(83, 8),
47477 => conv_std_logic_vector(84, 8),
47478 => conv_std_logic_vector(85, 8),
47479 => conv_std_logic_vector(85, 8),
47480 => conv_std_logic_vector(86, 8),
47481 => conv_std_logic_vector(87, 8),
47482 => conv_std_logic_vector(88, 8),
47483 => conv_std_logic_vector(88, 8),
47484 => conv_std_logic_vector(89, 8),
47485 => conv_std_logic_vector(90, 8),
47486 => conv_std_logic_vector(91, 8),
47487 => conv_std_logic_vector(91, 8),
47488 => conv_std_logic_vector(92, 8),
47489 => conv_std_logic_vector(93, 8),
47490 => conv_std_logic_vector(93, 8),
47491 => conv_std_logic_vector(94, 8),
47492 => conv_std_logic_vector(95, 8),
47493 => conv_std_logic_vector(96, 8),
47494 => conv_std_logic_vector(96, 8),
47495 => conv_std_logic_vector(97, 8),
47496 => conv_std_logic_vector(98, 8),
47497 => conv_std_logic_vector(99, 8),
47498 => conv_std_logic_vector(99, 8),
47499 => conv_std_logic_vector(100, 8),
47500 => conv_std_logic_vector(101, 8),
47501 => conv_std_logic_vector(101, 8),
47502 => conv_std_logic_vector(102, 8),
47503 => conv_std_logic_vector(103, 8),
47504 => conv_std_logic_vector(104, 8),
47505 => conv_std_logic_vector(104, 8),
47506 => conv_std_logic_vector(105, 8),
47507 => conv_std_logic_vector(106, 8),
47508 => conv_std_logic_vector(106, 8),
47509 => conv_std_logic_vector(107, 8),
47510 => conv_std_logic_vector(108, 8),
47511 => conv_std_logic_vector(109, 8),
47512 => conv_std_logic_vector(109, 8),
47513 => conv_std_logic_vector(110, 8),
47514 => conv_std_logic_vector(111, 8),
47515 => conv_std_logic_vector(112, 8),
47516 => conv_std_logic_vector(112, 8),
47517 => conv_std_logic_vector(113, 8),
47518 => conv_std_logic_vector(114, 8),
47519 => conv_std_logic_vector(114, 8),
47520 => conv_std_logic_vector(115, 8),
47521 => conv_std_logic_vector(116, 8),
47522 => conv_std_logic_vector(117, 8),
47523 => conv_std_logic_vector(117, 8),
47524 => conv_std_logic_vector(118, 8),
47525 => conv_std_logic_vector(119, 8),
47526 => conv_std_logic_vector(119, 8),
47527 => conv_std_logic_vector(120, 8),
47528 => conv_std_logic_vector(121, 8),
47529 => conv_std_logic_vector(122, 8),
47530 => conv_std_logic_vector(122, 8),
47531 => conv_std_logic_vector(123, 8),
47532 => conv_std_logic_vector(124, 8),
47533 => conv_std_logic_vector(125, 8),
47534 => conv_std_logic_vector(125, 8),
47535 => conv_std_logic_vector(126, 8),
47536 => conv_std_logic_vector(127, 8),
47537 => conv_std_logic_vector(127, 8),
47538 => conv_std_logic_vector(128, 8),
47539 => conv_std_logic_vector(129, 8),
47540 => conv_std_logic_vector(130, 8),
47541 => conv_std_logic_vector(130, 8),
47542 => conv_std_logic_vector(131, 8),
47543 => conv_std_logic_vector(132, 8),
47544 => conv_std_logic_vector(132, 8),
47545 => conv_std_logic_vector(133, 8),
47546 => conv_std_logic_vector(134, 8),
47547 => conv_std_logic_vector(135, 8),
47548 => conv_std_logic_vector(135, 8),
47549 => conv_std_logic_vector(136, 8),
47550 => conv_std_logic_vector(137, 8),
47551 => conv_std_logic_vector(138, 8),
47552 => conv_std_logic_vector(138, 8),
47553 => conv_std_logic_vector(139, 8),
47554 => conv_std_logic_vector(140, 8),
47555 => conv_std_logic_vector(140, 8),
47556 => conv_std_logic_vector(141, 8),
47557 => conv_std_logic_vector(142, 8),
47558 => conv_std_logic_vector(143, 8),
47559 => conv_std_logic_vector(143, 8),
47560 => conv_std_logic_vector(144, 8),
47561 => conv_std_logic_vector(145, 8),
47562 => conv_std_logic_vector(145, 8),
47563 => conv_std_logic_vector(146, 8),
47564 => conv_std_logic_vector(147, 8),
47565 => conv_std_logic_vector(148, 8),
47566 => conv_std_logic_vector(148, 8),
47567 => conv_std_logic_vector(149, 8),
47568 => conv_std_logic_vector(150, 8),
47569 => conv_std_logic_vector(151, 8),
47570 => conv_std_logic_vector(151, 8),
47571 => conv_std_logic_vector(152, 8),
47572 => conv_std_logic_vector(153, 8),
47573 => conv_std_logic_vector(153, 8),
47574 => conv_std_logic_vector(154, 8),
47575 => conv_std_logic_vector(155, 8),
47576 => conv_std_logic_vector(156, 8),
47577 => conv_std_logic_vector(156, 8),
47578 => conv_std_logic_vector(157, 8),
47579 => conv_std_logic_vector(158, 8),
47580 => conv_std_logic_vector(158, 8),
47581 => conv_std_logic_vector(159, 8),
47582 => conv_std_logic_vector(160, 8),
47583 => conv_std_logic_vector(161, 8),
47584 => conv_std_logic_vector(161, 8),
47585 => conv_std_logic_vector(162, 8),
47586 => conv_std_logic_vector(163, 8),
47587 => conv_std_logic_vector(164, 8),
47588 => conv_std_logic_vector(164, 8),
47589 => conv_std_logic_vector(165, 8),
47590 => conv_std_logic_vector(166, 8),
47591 => conv_std_logic_vector(166, 8),
47592 => conv_std_logic_vector(167, 8),
47593 => conv_std_logic_vector(168, 8),
47594 => conv_std_logic_vector(169, 8),
47595 => conv_std_logic_vector(169, 8),
47596 => conv_std_logic_vector(170, 8),
47597 => conv_std_logic_vector(171, 8),
47598 => conv_std_logic_vector(171, 8),
47599 => conv_std_logic_vector(172, 8),
47600 => conv_std_logic_vector(173, 8),
47601 => conv_std_logic_vector(174, 8),
47602 => conv_std_logic_vector(174, 8),
47603 => conv_std_logic_vector(175, 8),
47604 => conv_std_logic_vector(176, 8),
47605 => conv_std_logic_vector(177, 8),
47606 => conv_std_logic_vector(177, 8),
47607 => conv_std_logic_vector(178, 8),
47608 => conv_std_logic_vector(179, 8),
47609 => conv_std_logic_vector(179, 8),
47610 => conv_std_logic_vector(180, 8),
47611 => conv_std_logic_vector(181, 8),
47612 => conv_std_logic_vector(182, 8),
47613 => conv_std_logic_vector(182, 8),
47614 => conv_std_logic_vector(183, 8),
47615 => conv_std_logic_vector(184, 8),
47616 => conv_std_logic_vector(0, 8),
47617 => conv_std_logic_vector(0, 8),
47618 => conv_std_logic_vector(1, 8),
47619 => conv_std_logic_vector(2, 8),
47620 => conv_std_logic_vector(2, 8),
47621 => conv_std_logic_vector(3, 8),
47622 => conv_std_logic_vector(4, 8),
47623 => conv_std_logic_vector(5, 8),
47624 => conv_std_logic_vector(5, 8),
47625 => conv_std_logic_vector(6, 8),
47626 => conv_std_logic_vector(7, 8),
47627 => conv_std_logic_vector(7, 8),
47628 => conv_std_logic_vector(8, 8),
47629 => conv_std_logic_vector(9, 8),
47630 => conv_std_logic_vector(10, 8),
47631 => conv_std_logic_vector(10, 8),
47632 => conv_std_logic_vector(11, 8),
47633 => conv_std_logic_vector(12, 8),
47634 => conv_std_logic_vector(13, 8),
47635 => conv_std_logic_vector(13, 8),
47636 => conv_std_logic_vector(14, 8),
47637 => conv_std_logic_vector(15, 8),
47638 => conv_std_logic_vector(15, 8),
47639 => conv_std_logic_vector(16, 8),
47640 => conv_std_logic_vector(17, 8),
47641 => conv_std_logic_vector(18, 8),
47642 => conv_std_logic_vector(18, 8),
47643 => conv_std_logic_vector(19, 8),
47644 => conv_std_logic_vector(20, 8),
47645 => conv_std_logic_vector(21, 8),
47646 => conv_std_logic_vector(21, 8),
47647 => conv_std_logic_vector(22, 8),
47648 => conv_std_logic_vector(23, 8),
47649 => conv_std_logic_vector(23, 8),
47650 => conv_std_logic_vector(24, 8),
47651 => conv_std_logic_vector(25, 8),
47652 => conv_std_logic_vector(26, 8),
47653 => conv_std_logic_vector(26, 8),
47654 => conv_std_logic_vector(27, 8),
47655 => conv_std_logic_vector(28, 8),
47656 => conv_std_logic_vector(29, 8),
47657 => conv_std_logic_vector(29, 8),
47658 => conv_std_logic_vector(30, 8),
47659 => conv_std_logic_vector(31, 8),
47660 => conv_std_logic_vector(31, 8),
47661 => conv_std_logic_vector(32, 8),
47662 => conv_std_logic_vector(33, 8),
47663 => conv_std_logic_vector(34, 8),
47664 => conv_std_logic_vector(34, 8),
47665 => conv_std_logic_vector(35, 8),
47666 => conv_std_logic_vector(36, 8),
47667 => conv_std_logic_vector(37, 8),
47668 => conv_std_logic_vector(37, 8),
47669 => conv_std_logic_vector(38, 8),
47670 => conv_std_logic_vector(39, 8),
47671 => conv_std_logic_vector(39, 8),
47672 => conv_std_logic_vector(40, 8),
47673 => conv_std_logic_vector(41, 8),
47674 => conv_std_logic_vector(42, 8),
47675 => conv_std_logic_vector(42, 8),
47676 => conv_std_logic_vector(43, 8),
47677 => conv_std_logic_vector(44, 8),
47678 => conv_std_logic_vector(45, 8),
47679 => conv_std_logic_vector(45, 8),
47680 => conv_std_logic_vector(46, 8),
47681 => conv_std_logic_vector(47, 8),
47682 => conv_std_logic_vector(47, 8),
47683 => conv_std_logic_vector(48, 8),
47684 => conv_std_logic_vector(49, 8),
47685 => conv_std_logic_vector(50, 8),
47686 => conv_std_logic_vector(50, 8),
47687 => conv_std_logic_vector(51, 8),
47688 => conv_std_logic_vector(52, 8),
47689 => conv_std_logic_vector(53, 8),
47690 => conv_std_logic_vector(53, 8),
47691 => conv_std_logic_vector(54, 8),
47692 => conv_std_logic_vector(55, 8),
47693 => conv_std_logic_vector(55, 8),
47694 => conv_std_logic_vector(56, 8),
47695 => conv_std_logic_vector(57, 8),
47696 => conv_std_logic_vector(58, 8),
47697 => conv_std_logic_vector(58, 8),
47698 => conv_std_logic_vector(59, 8),
47699 => conv_std_logic_vector(60, 8),
47700 => conv_std_logic_vector(61, 8),
47701 => conv_std_logic_vector(61, 8),
47702 => conv_std_logic_vector(62, 8),
47703 => conv_std_logic_vector(63, 8),
47704 => conv_std_logic_vector(63, 8),
47705 => conv_std_logic_vector(64, 8),
47706 => conv_std_logic_vector(65, 8),
47707 => conv_std_logic_vector(66, 8),
47708 => conv_std_logic_vector(66, 8),
47709 => conv_std_logic_vector(67, 8),
47710 => conv_std_logic_vector(68, 8),
47711 => conv_std_logic_vector(69, 8),
47712 => conv_std_logic_vector(69, 8),
47713 => conv_std_logic_vector(70, 8),
47714 => conv_std_logic_vector(71, 8),
47715 => conv_std_logic_vector(71, 8),
47716 => conv_std_logic_vector(72, 8),
47717 => conv_std_logic_vector(73, 8),
47718 => conv_std_logic_vector(74, 8),
47719 => conv_std_logic_vector(74, 8),
47720 => conv_std_logic_vector(75, 8),
47721 => conv_std_logic_vector(76, 8),
47722 => conv_std_logic_vector(77, 8),
47723 => conv_std_logic_vector(77, 8),
47724 => conv_std_logic_vector(78, 8),
47725 => conv_std_logic_vector(79, 8),
47726 => conv_std_logic_vector(79, 8),
47727 => conv_std_logic_vector(80, 8),
47728 => conv_std_logic_vector(81, 8),
47729 => conv_std_logic_vector(82, 8),
47730 => conv_std_logic_vector(82, 8),
47731 => conv_std_logic_vector(83, 8),
47732 => conv_std_logic_vector(84, 8),
47733 => conv_std_logic_vector(85, 8),
47734 => conv_std_logic_vector(85, 8),
47735 => conv_std_logic_vector(86, 8),
47736 => conv_std_logic_vector(87, 8),
47737 => conv_std_logic_vector(87, 8),
47738 => conv_std_logic_vector(88, 8),
47739 => conv_std_logic_vector(89, 8),
47740 => conv_std_logic_vector(90, 8),
47741 => conv_std_logic_vector(90, 8),
47742 => conv_std_logic_vector(91, 8),
47743 => conv_std_logic_vector(92, 8),
47744 => conv_std_logic_vector(93, 8),
47745 => conv_std_logic_vector(93, 8),
47746 => conv_std_logic_vector(94, 8),
47747 => conv_std_logic_vector(95, 8),
47748 => conv_std_logic_vector(95, 8),
47749 => conv_std_logic_vector(96, 8),
47750 => conv_std_logic_vector(97, 8),
47751 => conv_std_logic_vector(98, 8),
47752 => conv_std_logic_vector(98, 8),
47753 => conv_std_logic_vector(99, 8),
47754 => conv_std_logic_vector(100, 8),
47755 => conv_std_logic_vector(100, 8),
47756 => conv_std_logic_vector(101, 8),
47757 => conv_std_logic_vector(102, 8),
47758 => conv_std_logic_vector(103, 8),
47759 => conv_std_logic_vector(103, 8),
47760 => conv_std_logic_vector(104, 8),
47761 => conv_std_logic_vector(105, 8),
47762 => conv_std_logic_vector(106, 8),
47763 => conv_std_logic_vector(106, 8),
47764 => conv_std_logic_vector(107, 8),
47765 => conv_std_logic_vector(108, 8),
47766 => conv_std_logic_vector(108, 8),
47767 => conv_std_logic_vector(109, 8),
47768 => conv_std_logic_vector(110, 8),
47769 => conv_std_logic_vector(111, 8),
47770 => conv_std_logic_vector(111, 8),
47771 => conv_std_logic_vector(112, 8),
47772 => conv_std_logic_vector(113, 8),
47773 => conv_std_logic_vector(114, 8),
47774 => conv_std_logic_vector(114, 8),
47775 => conv_std_logic_vector(115, 8),
47776 => conv_std_logic_vector(116, 8),
47777 => conv_std_logic_vector(116, 8),
47778 => conv_std_logic_vector(117, 8),
47779 => conv_std_logic_vector(118, 8),
47780 => conv_std_logic_vector(119, 8),
47781 => conv_std_logic_vector(119, 8),
47782 => conv_std_logic_vector(120, 8),
47783 => conv_std_logic_vector(121, 8),
47784 => conv_std_logic_vector(122, 8),
47785 => conv_std_logic_vector(122, 8),
47786 => conv_std_logic_vector(123, 8),
47787 => conv_std_logic_vector(124, 8),
47788 => conv_std_logic_vector(124, 8),
47789 => conv_std_logic_vector(125, 8),
47790 => conv_std_logic_vector(126, 8),
47791 => conv_std_logic_vector(127, 8),
47792 => conv_std_logic_vector(127, 8),
47793 => conv_std_logic_vector(128, 8),
47794 => conv_std_logic_vector(129, 8),
47795 => conv_std_logic_vector(130, 8),
47796 => conv_std_logic_vector(130, 8),
47797 => conv_std_logic_vector(131, 8),
47798 => conv_std_logic_vector(132, 8),
47799 => conv_std_logic_vector(132, 8),
47800 => conv_std_logic_vector(133, 8),
47801 => conv_std_logic_vector(134, 8),
47802 => conv_std_logic_vector(135, 8),
47803 => conv_std_logic_vector(135, 8),
47804 => conv_std_logic_vector(136, 8),
47805 => conv_std_logic_vector(137, 8),
47806 => conv_std_logic_vector(138, 8),
47807 => conv_std_logic_vector(138, 8),
47808 => conv_std_logic_vector(139, 8),
47809 => conv_std_logic_vector(140, 8),
47810 => conv_std_logic_vector(140, 8),
47811 => conv_std_logic_vector(141, 8),
47812 => conv_std_logic_vector(142, 8),
47813 => conv_std_logic_vector(143, 8),
47814 => conv_std_logic_vector(143, 8),
47815 => conv_std_logic_vector(144, 8),
47816 => conv_std_logic_vector(145, 8),
47817 => conv_std_logic_vector(146, 8),
47818 => conv_std_logic_vector(146, 8),
47819 => conv_std_logic_vector(147, 8),
47820 => conv_std_logic_vector(148, 8),
47821 => conv_std_logic_vector(148, 8),
47822 => conv_std_logic_vector(149, 8),
47823 => conv_std_logic_vector(150, 8),
47824 => conv_std_logic_vector(151, 8),
47825 => conv_std_logic_vector(151, 8),
47826 => conv_std_logic_vector(152, 8),
47827 => conv_std_logic_vector(153, 8),
47828 => conv_std_logic_vector(154, 8),
47829 => conv_std_logic_vector(154, 8),
47830 => conv_std_logic_vector(155, 8),
47831 => conv_std_logic_vector(156, 8),
47832 => conv_std_logic_vector(156, 8),
47833 => conv_std_logic_vector(157, 8),
47834 => conv_std_logic_vector(158, 8),
47835 => conv_std_logic_vector(159, 8),
47836 => conv_std_logic_vector(159, 8),
47837 => conv_std_logic_vector(160, 8),
47838 => conv_std_logic_vector(161, 8),
47839 => conv_std_logic_vector(162, 8),
47840 => conv_std_logic_vector(162, 8),
47841 => conv_std_logic_vector(163, 8),
47842 => conv_std_logic_vector(164, 8),
47843 => conv_std_logic_vector(164, 8),
47844 => conv_std_logic_vector(165, 8),
47845 => conv_std_logic_vector(166, 8),
47846 => conv_std_logic_vector(167, 8),
47847 => conv_std_logic_vector(167, 8),
47848 => conv_std_logic_vector(168, 8),
47849 => conv_std_logic_vector(169, 8),
47850 => conv_std_logic_vector(170, 8),
47851 => conv_std_logic_vector(170, 8),
47852 => conv_std_logic_vector(171, 8),
47853 => conv_std_logic_vector(172, 8),
47854 => conv_std_logic_vector(172, 8),
47855 => conv_std_logic_vector(173, 8),
47856 => conv_std_logic_vector(174, 8),
47857 => conv_std_logic_vector(175, 8),
47858 => conv_std_logic_vector(175, 8),
47859 => conv_std_logic_vector(176, 8),
47860 => conv_std_logic_vector(177, 8),
47861 => conv_std_logic_vector(178, 8),
47862 => conv_std_logic_vector(178, 8),
47863 => conv_std_logic_vector(179, 8),
47864 => conv_std_logic_vector(180, 8),
47865 => conv_std_logic_vector(180, 8),
47866 => conv_std_logic_vector(181, 8),
47867 => conv_std_logic_vector(182, 8),
47868 => conv_std_logic_vector(183, 8),
47869 => conv_std_logic_vector(183, 8),
47870 => conv_std_logic_vector(184, 8),
47871 => conv_std_logic_vector(185, 8),
47872 => conv_std_logic_vector(0, 8),
47873 => conv_std_logic_vector(0, 8),
47874 => conv_std_logic_vector(1, 8),
47875 => conv_std_logic_vector(2, 8),
47876 => conv_std_logic_vector(2, 8),
47877 => conv_std_logic_vector(3, 8),
47878 => conv_std_logic_vector(4, 8),
47879 => conv_std_logic_vector(5, 8),
47880 => conv_std_logic_vector(5, 8),
47881 => conv_std_logic_vector(6, 8),
47882 => conv_std_logic_vector(7, 8),
47883 => conv_std_logic_vector(8, 8),
47884 => conv_std_logic_vector(8, 8),
47885 => conv_std_logic_vector(9, 8),
47886 => conv_std_logic_vector(10, 8),
47887 => conv_std_logic_vector(10, 8),
47888 => conv_std_logic_vector(11, 8),
47889 => conv_std_logic_vector(12, 8),
47890 => conv_std_logic_vector(13, 8),
47891 => conv_std_logic_vector(13, 8),
47892 => conv_std_logic_vector(14, 8),
47893 => conv_std_logic_vector(15, 8),
47894 => conv_std_logic_vector(16, 8),
47895 => conv_std_logic_vector(16, 8),
47896 => conv_std_logic_vector(17, 8),
47897 => conv_std_logic_vector(18, 8),
47898 => conv_std_logic_vector(18, 8),
47899 => conv_std_logic_vector(19, 8),
47900 => conv_std_logic_vector(20, 8),
47901 => conv_std_logic_vector(21, 8),
47902 => conv_std_logic_vector(21, 8),
47903 => conv_std_logic_vector(22, 8),
47904 => conv_std_logic_vector(23, 8),
47905 => conv_std_logic_vector(24, 8),
47906 => conv_std_logic_vector(24, 8),
47907 => conv_std_logic_vector(25, 8),
47908 => conv_std_logic_vector(26, 8),
47909 => conv_std_logic_vector(27, 8),
47910 => conv_std_logic_vector(27, 8),
47911 => conv_std_logic_vector(28, 8),
47912 => conv_std_logic_vector(29, 8),
47913 => conv_std_logic_vector(29, 8),
47914 => conv_std_logic_vector(30, 8),
47915 => conv_std_logic_vector(31, 8),
47916 => conv_std_logic_vector(32, 8),
47917 => conv_std_logic_vector(32, 8),
47918 => conv_std_logic_vector(33, 8),
47919 => conv_std_logic_vector(34, 8),
47920 => conv_std_logic_vector(35, 8),
47921 => conv_std_logic_vector(35, 8),
47922 => conv_std_logic_vector(36, 8),
47923 => conv_std_logic_vector(37, 8),
47924 => conv_std_logic_vector(37, 8),
47925 => conv_std_logic_vector(38, 8),
47926 => conv_std_logic_vector(39, 8),
47927 => conv_std_logic_vector(40, 8),
47928 => conv_std_logic_vector(40, 8),
47929 => conv_std_logic_vector(41, 8),
47930 => conv_std_logic_vector(42, 8),
47931 => conv_std_logic_vector(43, 8),
47932 => conv_std_logic_vector(43, 8),
47933 => conv_std_logic_vector(44, 8),
47934 => conv_std_logic_vector(45, 8),
47935 => conv_std_logic_vector(46, 8),
47936 => conv_std_logic_vector(46, 8),
47937 => conv_std_logic_vector(47, 8),
47938 => conv_std_logic_vector(48, 8),
47939 => conv_std_logic_vector(48, 8),
47940 => conv_std_logic_vector(49, 8),
47941 => conv_std_logic_vector(50, 8),
47942 => conv_std_logic_vector(51, 8),
47943 => conv_std_logic_vector(51, 8),
47944 => conv_std_logic_vector(52, 8),
47945 => conv_std_logic_vector(53, 8),
47946 => conv_std_logic_vector(54, 8),
47947 => conv_std_logic_vector(54, 8),
47948 => conv_std_logic_vector(55, 8),
47949 => conv_std_logic_vector(56, 8),
47950 => conv_std_logic_vector(56, 8),
47951 => conv_std_logic_vector(57, 8),
47952 => conv_std_logic_vector(58, 8),
47953 => conv_std_logic_vector(59, 8),
47954 => conv_std_logic_vector(59, 8),
47955 => conv_std_logic_vector(60, 8),
47956 => conv_std_logic_vector(61, 8),
47957 => conv_std_logic_vector(62, 8),
47958 => conv_std_logic_vector(62, 8),
47959 => conv_std_logic_vector(63, 8),
47960 => conv_std_logic_vector(64, 8),
47961 => conv_std_logic_vector(65, 8),
47962 => conv_std_logic_vector(65, 8),
47963 => conv_std_logic_vector(66, 8),
47964 => conv_std_logic_vector(67, 8),
47965 => conv_std_logic_vector(67, 8),
47966 => conv_std_logic_vector(68, 8),
47967 => conv_std_logic_vector(69, 8),
47968 => conv_std_logic_vector(70, 8),
47969 => conv_std_logic_vector(70, 8),
47970 => conv_std_logic_vector(71, 8),
47971 => conv_std_logic_vector(72, 8),
47972 => conv_std_logic_vector(73, 8),
47973 => conv_std_logic_vector(73, 8),
47974 => conv_std_logic_vector(74, 8),
47975 => conv_std_logic_vector(75, 8),
47976 => conv_std_logic_vector(75, 8),
47977 => conv_std_logic_vector(76, 8),
47978 => conv_std_logic_vector(77, 8),
47979 => conv_std_logic_vector(78, 8),
47980 => conv_std_logic_vector(78, 8),
47981 => conv_std_logic_vector(79, 8),
47982 => conv_std_logic_vector(80, 8),
47983 => conv_std_logic_vector(81, 8),
47984 => conv_std_logic_vector(81, 8),
47985 => conv_std_logic_vector(82, 8),
47986 => conv_std_logic_vector(83, 8),
47987 => conv_std_logic_vector(84, 8),
47988 => conv_std_logic_vector(84, 8),
47989 => conv_std_logic_vector(85, 8),
47990 => conv_std_logic_vector(86, 8),
47991 => conv_std_logic_vector(86, 8),
47992 => conv_std_logic_vector(87, 8),
47993 => conv_std_logic_vector(88, 8),
47994 => conv_std_logic_vector(89, 8),
47995 => conv_std_logic_vector(89, 8),
47996 => conv_std_logic_vector(90, 8),
47997 => conv_std_logic_vector(91, 8),
47998 => conv_std_logic_vector(92, 8),
47999 => conv_std_logic_vector(92, 8),
48000 => conv_std_logic_vector(93, 8),
48001 => conv_std_logic_vector(94, 8),
48002 => conv_std_logic_vector(94, 8),
48003 => conv_std_logic_vector(95, 8),
48004 => conv_std_logic_vector(96, 8),
48005 => conv_std_logic_vector(97, 8),
48006 => conv_std_logic_vector(97, 8),
48007 => conv_std_logic_vector(98, 8),
48008 => conv_std_logic_vector(99, 8),
48009 => conv_std_logic_vector(100, 8),
48010 => conv_std_logic_vector(100, 8),
48011 => conv_std_logic_vector(101, 8),
48012 => conv_std_logic_vector(102, 8),
48013 => conv_std_logic_vector(102, 8),
48014 => conv_std_logic_vector(103, 8),
48015 => conv_std_logic_vector(104, 8),
48016 => conv_std_logic_vector(105, 8),
48017 => conv_std_logic_vector(105, 8),
48018 => conv_std_logic_vector(106, 8),
48019 => conv_std_logic_vector(107, 8),
48020 => conv_std_logic_vector(108, 8),
48021 => conv_std_logic_vector(108, 8),
48022 => conv_std_logic_vector(109, 8),
48023 => conv_std_logic_vector(110, 8),
48024 => conv_std_logic_vector(111, 8),
48025 => conv_std_logic_vector(111, 8),
48026 => conv_std_logic_vector(112, 8),
48027 => conv_std_logic_vector(113, 8),
48028 => conv_std_logic_vector(113, 8),
48029 => conv_std_logic_vector(114, 8),
48030 => conv_std_logic_vector(115, 8),
48031 => conv_std_logic_vector(116, 8),
48032 => conv_std_logic_vector(116, 8),
48033 => conv_std_logic_vector(117, 8),
48034 => conv_std_logic_vector(118, 8),
48035 => conv_std_logic_vector(119, 8),
48036 => conv_std_logic_vector(119, 8),
48037 => conv_std_logic_vector(120, 8),
48038 => conv_std_logic_vector(121, 8),
48039 => conv_std_logic_vector(121, 8),
48040 => conv_std_logic_vector(122, 8),
48041 => conv_std_logic_vector(123, 8),
48042 => conv_std_logic_vector(124, 8),
48043 => conv_std_logic_vector(124, 8),
48044 => conv_std_logic_vector(125, 8),
48045 => conv_std_logic_vector(126, 8),
48046 => conv_std_logic_vector(127, 8),
48047 => conv_std_logic_vector(127, 8),
48048 => conv_std_logic_vector(128, 8),
48049 => conv_std_logic_vector(129, 8),
48050 => conv_std_logic_vector(130, 8),
48051 => conv_std_logic_vector(130, 8),
48052 => conv_std_logic_vector(131, 8),
48053 => conv_std_logic_vector(132, 8),
48054 => conv_std_logic_vector(132, 8),
48055 => conv_std_logic_vector(133, 8),
48056 => conv_std_logic_vector(134, 8),
48057 => conv_std_logic_vector(135, 8),
48058 => conv_std_logic_vector(135, 8),
48059 => conv_std_logic_vector(136, 8),
48060 => conv_std_logic_vector(137, 8),
48061 => conv_std_logic_vector(138, 8),
48062 => conv_std_logic_vector(138, 8),
48063 => conv_std_logic_vector(139, 8),
48064 => conv_std_logic_vector(140, 8),
48065 => conv_std_logic_vector(140, 8),
48066 => conv_std_logic_vector(141, 8),
48067 => conv_std_logic_vector(142, 8),
48068 => conv_std_logic_vector(143, 8),
48069 => conv_std_logic_vector(143, 8),
48070 => conv_std_logic_vector(144, 8),
48071 => conv_std_logic_vector(145, 8),
48072 => conv_std_logic_vector(146, 8),
48073 => conv_std_logic_vector(146, 8),
48074 => conv_std_logic_vector(147, 8),
48075 => conv_std_logic_vector(148, 8),
48076 => conv_std_logic_vector(149, 8),
48077 => conv_std_logic_vector(149, 8),
48078 => conv_std_logic_vector(150, 8),
48079 => conv_std_logic_vector(151, 8),
48080 => conv_std_logic_vector(151, 8),
48081 => conv_std_logic_vector(152, 8),
48082 => conv_std_logic_vector(153, 8),
48083 => conv_std_logic_vector(154, 8),
48084 => conv_std_logic_vector(154, 8),
48085 => conv_std_logic_vector(155, 8),
48086 => conv_std_logic_vector(156, 8),
48087 => conv_std_logic_vector(157, 8),
48088 => conv_std_logic_vector(157, 8),
48089 => conv_std_logic_vector(158, 8),
48090 => conv_std_logic_vector(159, 8),
48091 => conv_std_logic_vector(159, 8),
48092 => conv_std_logic_vector(160, 8),
48093 => conv_std_logic_vector(161, 8),
48094 => conv_std_logic_vector(162, 8),
48095 => conv_std_logic_vector(162, 8),
48096 => conv_std_logic_vector(163, 8),
48097 => conv_std_logic_vector(164, 8),
48098 => conv_std_logic_vector(165, 8),
48099 => conv_std_logic_vector(165, 8),
48100 => conv_std_logic_vector(166, 8),
48101 => conv_std_logic_vector(167, 8),
48102 => conv_std_logic_vector(168, 8),
48103 => conv_std_logic_vector(168, 8),
48104 => conv_std_logic_vector(169, 8),
48105 => conv_std_logic_vector(170, 8),
48106 => conv_std_logic_vector(170, 8),
48107 => conv_std_logic_vector(171, 8),
48108 => conv_std_logic_vector(172, 8),
48109 => conv_std_logic_vector(173, 8),
48110 => conv_std_logic_vector(173, 8),
48111 => conv_std_logic_vector(174, 8),
48112 => conv_std_logic_vector(175, 8),
48113 => conv_std_logic_vector(176, 8),
48114 => conv_std_logic_vector(176, 8),
48115 => conv_std_logic_vector(177, 8),
48116 => conv_std_logic_vector(178, 8),
48117 => conv_std_logic_vector(178, 8),
48118 => conv_std_logic_vector(179, 8),
48119 => conv_std_logic_vector(180, 8),
48120 => conv_std_logic_vector(181, 8),
48121 => conv_std_logic_vector(181, 8),
48122 => conv_std_logic_vector(182, 8),
48123 => conv_std_logic_vector(183, 8),
48124 => conv_std_logic_vector(184, 8),
48125 => conv_std_logic_vector(184, 8),
48126 => conv_std_logic_vector(185, 8),
48127 => conv_std_logic_vector(186, 8),
48128 => conv_std_logic_vector(0, 8),
48129 => conv_std_logic_vector(0, 8),
48130 => conv_std_logic_vector(1, 8),
48131 => conv_std_logic_vector(2, 8),
48132 => conv_std_logic_vector(2, 8),
48133 => conv_std_logic_vector(3, 8),
48134 => conv_std_logic_vector(4, 8),
48135 => conv_std_logic_vector(5, 8),
48136 => conv_std_logic_vector(5, 8),
48137 => conv_std_logic_vector(6, 8),
48138 => conv_std_logic_vector(7, 8),
48139 => conv_std_logic_vector(8, 8),
48140 => conv_std_logic_vector(8, 8),
48141 => conv_std_logic_vector(9, 8),
48142 => conv_std_logic_vector(10, 8),
48143 => conv_std_logic_vector(11, 8),
48144 => conv_std_logic_vector(11, 8),
48145 => conv_std_logic_vector(12, 8),
48146 => conv_std_logic_vector(13, 8),
48147 => conv_std_logic_vector(13, 8),
48148 => conv_std_logic_vector(14, 8),
48149 => conv_std_logic_vector(15, 8),
48150 => conv_std_logic_vector(16, 8),
48151 => conv_std_logic_vector(16, 8),
48152 => conv_std_logic_vector(17, 8),
48153 => conv_std_logic_vector(18, 8),
48154 => conv_std_logic_vector(19, 8),
48155 => conv_std_logic_vector(19, 8),
48156 => conv_std_logic_vector(20, 8),
48157 => conv_std_logic_vector(21, 8),
48158 => conv_std_logic_vector(22, 8),
48159 => conv_std_logic_vector(22, 8),
48160 => conv_std_logic_vector(23, 8),
48161 => conv_std_logic_vector(24, 8),
48162 => conv_std_logic_vector(24, 8),
48163 => conv_std_logic_vector(25, 8),
48164 => conv_std_logic_vector(26, 8),
48165 => conv_std_logic_vector(27, 8),
48166 => conv_std_logic_vector(27, 8),
48167 => conv_std_logic_vector(28, 8),
48168 => conv_std_logic_vector(29, 8),
48169 => conv_std_logic_vector(30, 8),
48170 => conv_std_logic_vector(30, 8),
48171 => conv_std_logic_vector(31, 8),
48172 => conv_std_logic_vector(32, 8),
48173 => conv_std_logic_vector(33, 8),
48174 => conv_std_logic_vector(33, 8),
48175 => conv_std_logic_vector(34, 8),
48176 => conv_std_logic_vector(35, 8),
48177 => conv_std_logic_vector(35, 8),
48178 => conv_std_logic_vector(36, 8),
48179 => conv_std_logic_vector(37, 8),
48180 => conv_std_logic_vector(38, 8),
48181 => conv_std_logic_vector(38, 8),
48182 => conv_std_logic_vector(39, 8),
48183 => conv_std_logic_vector(40, 8),
48184 => conv_std_logic_vector(41, 8),
48185 => conv_std_logic_vector(41, 8),
48186 => conv_std_logic_vector(42, 8),
48187 => conv_std_logic_vector(43, 8),
48188 => conv_std_logic_vector(44, 8),
48189 => conv_std_logic_vector(44, 8),
48190 => conv_std_logic_vector(45, 8),
48191 => conv_std_logic_vector(46, 8),
48192 => conv_std_logic_vector(47, 8),
48193 => conv_std_logic_vector(47, 8),
48194 => conv_std_logic_vector(48, 8),
48195 => conv_std_logic_vector(49, 8),
48196 => conv_std_logic_vector(49, 8),
48197 => conv_std_logic_vector(50, 8),
48198 => conv_std_logic_vector(51, 8),
48199 => conv_std_logic_vector(52, 8),
48200 => conv_std_logic_vector(52, 8),
48201 => conv_std_logic_vector(53, 8),
48202 => conv_std_logic_vector(54, 8),
48203 => conv_std_logic_vector(55, 8),
48204 => conv_std_logic_vector(55, 8),
48205 => conv_std_logic_vector(56, 8),
48206 => conv_std_logic_vector(57, 8),
48207 => conv_std_logic_vector(58, 8),
48208 => conv_std_logic_vector(58, 8),
48209 => conv_std_logic_vector(59, 8),
48210 => conv_std_logic_vector(60, 8),
48211 => conv_std_logic_vector(60, 8),
48212 => conv_std_logic_vector(61, 8),
48213 => conv_std_logic_vector(62, 8),
48214 => conv_std_logic_vector(63, 8),
48215 => conv_std_logic_vector(63, 8),
48216 => conv_std_logic_vector(64, 8),
48217 => conv_std_logic_vector(65, 8),
48218 => conv_std_logic_vector(66, 8),
48219 => conv_std_logic_vector(66, 8),
48220 => conv_std_logic_vector(67, 8),
48221 => conv_std_logic_vector(68, 8),
48222 => conv_std_logic_vector(69, 8),
48223 => conv_std_logic_vector(69, 8),
48224 => conv_std_logic_vector(70, 8),
48225 => conv_std_logic_vector(71, 8),
48226 => conv_std_logic_vector(71, 8),
48227 => conv_std_logic_vector(72, 8),
48228 => conv_std_logic_vector(73, 8),
48229 => conv_std_logic_vector(74, 8),
48230 => conv_std_logic_vector(74, 8),
48231 => conv_std_logic_vector(75, 8),
48232 => conv_std_logic_vector(76, 8),
48233 => conv_std_logic_vector(77, 8),
48234 => conv_std_logic_vector(77, 8),
48235 => conv_std_logic_vector(78, 8),
48236 => conv_std_logic_vector(79, 8),
48237 => conv_std_logic_vector(80, 8),
48238 => conv_std_logic_vector(80, 8),
48239 => conv_std_logic_vector(81, 8),
48240 => conv_std_logic_vector(82, 8),
48241 => conv_std_logic_vector(82, 8),
48242 => conv_std_logic_vector(83, 8),
48243 => conv_std_logic_vector(84, 8),
48244 => conv_std_logic_vector(85, 8),
48245 => conv_std_logic_vector(85, 8),
48246 => conv_std_logic_vector(86, 8),
48247 => conv_std_logic_vector(87, 8),
48248 => conv_std_logic_vector(88, 8),
48249 => conv_std_logic_vector(88, 8),
48250 => conv_std_logic_vector(89, 8),
48251 => conv_std_logic_vector(90, 8),
48252 => conv_std_logic_vector(91, 8),
48253 => conv_std_logic_vector(91, 8),
48254 => conv_std_logic_vector(92, 8),
48255 => conv_std_logic_vector(93, 8),
48256 => conv_std_logic_vector(94, 8),
48257 => conv_std_logic_vector(94, 8),
48258 => conv_std_logic_vector(95, 8),
48259 => conv_std_logic_vector(96, 8),
48260 => conv_std_logic_vector(96, 8),
48261 => conv_std_logic_vector(97, 8),
48262 => conv_std_logic_vector(98, 8),
48263 => conv_std_logic_vector(99, 8),
48264 => conv_std_logic_vector(99, 8),
48265 => conv_std_logic_vector(100, 8),
48266 => conv_std_logic_vector(101, 8),
48267 => conv_std_logic_vector(102, 8),
48268 => conv_std_logic_vector(102, 8),
48269 => conv_std_logic_vector(103, 8),
48270 => conv_std_logic_vector(104, 8),
48271 => conv_std_logic_vector(105, 8),
48272 => conv_std_logic_vector(105, 8),
48273 => conv_std_logic_vector(106, 8),
48274 => conv_std_logic_vector(107, 8),
48275 => conv_std_logic_vector(107, 8),
48276 => conv_std_logic_vector(108, 8),
48277 => conv_std_logic_vector(109, 8),
48278 => conv_std_logic_vector(110, 8),
48279 => conv_std_logic_vector(110, 8),
48280 => conv_std_logic_vector(111, 8),
48281 => conv_std_logic_vector(112, 8),
48282 => conv_std_logic_vector(113, 8),
48283 => conv_std_logic_vector(113, 8),
48284 => conv_std_logic_vector(114, 8),
48285 => conv_std_logic_vector(115, 8),
48286 => conv_std_logic_vector(116, 8),
48287 => conv_std_logic_vector(116, 8),
48288 => conv_std_logic_vector(117, 8),
48289 => conv_std_logic_vector(118, 8),
48290 => conv_std_logic_vector(118, 8),
48291 => conv_std_logic_vector(119, 8),
48292 => conv_std_logic_vector(120, 8),
48293 => conv_std_logic_vector(121, 8),
48294 => conv_std_logic_vector(121, 8),
48295 => conv_std_logic_vector(122, 8),
48296 => conv_std_logic_vector(123, 8),
48297 => conv_std_logic_vector(124, 8),
48298 => conv_std_logic_vector(124, 8),
48299 => conv_std_logic_vector(125, 8),
48300 => conv_std_logic_vector(126, 8),
48301 => conv_std_logic_vector(127, 8),
48302 => conv_std_logic_vector(127, 8),
48303 => conv_std_logic_vector(128, 8),
48304 => conv_std_logic_vector(129, 8),
48305 => conv_std_logic_vector(129, 8),
48306 => conv_std_logic_vector(130, 8),
48307 => conv_std_logic_vector(131, 8),
48308 => conv_std_logic_vector(132, 8),
48309 => conv_std_logic_vector(132, 8),
48310 => conv_std_logic_vector(133, 8),
48311 => conv_std_logic_vector(134, 8),
48312 => conv_std_logic_vector(135, 8),
48313 => conv_std_logic_vector(135, 8),
48314 => conv_std_logic_vector(136, 8),
48315 => conv_std_logic_vector(137, 8),
48316 => conv_std_logic_vector(138, 8),
48317 => conv_std_logic_vector(138, 8),
48318 => conv_std_logic_vector(139, 8),
48319 => conv_std_logic_vector(140, 8),
48320 => conv_std_logic_vector(141, 8),
48321 => conv_std_logic_vector(141, 8),
48322 => conv_std_logic_vector(142, 8),
48323 => conv_std_logic_vector(143, 8),
48324 => conv_std_logic_vector(143, 8),
48325 => conv_std_logic_vector(144, 8),
48326 => conv_std_logic_vector(145, 8),
48327 => conv_std_logic_vector(146, 8),
48328 => conv_std_logic_vector(146, 8),
48329 => conv_std_logic_vector(147, 8),
48330 => conv_std_logic_vector(148, 8),
48331 => conv_std_logic_vector(149, 8),
48332 => conv_std_logic_vector(149, 8),
48333 => conv_std_logic_vector(150, 8),
48334 => conv_std_logic_vector(151, 8),
48335 => conv_std_logic_vector(152, 8),
48336 => conv_std_logic_vector(152, 8),
48337 => conv_std_logic_vector(153, 8),
48338 => conv_std_logic_vector(154, 8),
48339 => conv_std_logic_vector(154, 8),
48340 => conv_std_logic_vector(155, 8),
48341 => conv_std_logic_vector(156, 8),
48342 => conv_std_logic_vector(157, 8),
48343 => conv_std_logic_vector(157, 8),
48344 => conv_std_logic_vector(158, 8),
48345 => conv_std_logic_vector(159, 8),
48346 => conv_std_logic_vector(160, 8),
48347 => conv_std_logic_vector(160, 8),
48348 => conv_std_logic_vector(161, 8),
48349 => conv_std_logic_vector(162, 8),
48350 => conv_std_logic_vector(163, 8),
48351 => conv_std_logic_vector(163, 8),
48352 => conv_std_logic_vector(164, 8),
48353 => conv_std_logic_vector(165, 8),
48354 => conv_std_logic_vector(165, 8),
48355 => conv_std_logic_vector(166, 8),
48356 => conv_std_logic_vector(167, 8),
48357 => conv_std_logic_vector(168, 8),
48358 => conv_std_logic_vector(168, 8),
48359 => conv_std_logic_vector(169, 8),
48360 => conv_std_logic_vector(170, 8),
48361 => conv_std_logic_vector(171, 8),
48362 => conv_std_logic_vector(171, 8),
48363 => conv_std_logic_vector(172, 8),
48364 => conv_std_logic_vector(173, 8),
48365 => conv_std_logic_vector(174, 8),
48366 => conv_std_logic_vector(174, 8),
48367 => conv_std_logic_vector(175, 8),
48368 => conv_std_logic_vector(176, 8),
48369 => conv_std_logic_vector(176, 8),
48370 => conv_std_logic_vector(177, 8),
48371 => conv_std_logic_vector(178, 8),
48372 => conv_std_logic_vector(179, 8),
48373 => conv_std_logic_vector(179, 8),
48374 => conv_std_logic_vector(180, 8),
48375 => conv_std_logic_vector(181, 8),
48376 => conv_std_logic_vector(182, 8),
48377 => conv_std_logic_vector(182, 8),
48378 => conv_std_logic_vector(183, 8),
48379 => conv_std_logic_vector(184, 8),
48380 => conv_std_logic_vector(185, 8),
48381 => conv_std_logic_vector(185, 8),
48382 => conv_std_logic_vector(186, 8),
48383 => conv_std_logic_vector(187, 8),
48384 => conv_std_logic_vector(0, 8),
48385 => conv_std_logic_vector(0, 8),
48386 => conv_std_logic_vector(1, 8),
48387 => conv_std_logic_vector(2, 8),
48388 => conv_std_logic_vector(2, 8),
48389 => conv_std_logic_vector(3, 8),
48390 => conv_std_logic_vector(4, 8),
48391 => conv_std_logic_vector(5, 8),
48392 => conv_std_logic_vector(5, 8),
48393 => conv_std_logic_vector(6, 8),
48394 => conv_std_logic_vector(7, 8),
48395 => conv_std_logic_vector(8, 8),
48396 => conv_std_logic_vector(8, 8),
48397 => conv_std_logic_vector(9, 8),
48398 => conv_std_logic_vector(10, 8),
48399 => conv_std_logic_vector(11, 8),
48400 => conv_std_logic_vector(11, 8),
48401 => conv_std_logic_vector(12, 8),
48402 => conv_std_logic_vector(13, 8),
48403 => conv_std_logic_vector(14, 8),
48404 => conv_std_logic_vector(14, 8),
48405 => conv_std_logic_vector(15, 8),
48406 => conv_std_logic_vector(16, 8),
48407 => conv_std_logic_vector(16, 8),
48408 => conv_std_logic_vector(17, 8),
48409 => conv_std_logic_vector(18, 8),
48410 => conv_std_logic_vector(19, 8),
48411 => conv_std_logic_vector(19, 8),
48412 => conv_std_logic_vector(20, 8),
48413 => conv_std_logic_vector(21, 8),
48414 => conv_std_logic_vector(22, 8),
48415 => conv_std_logic_vector(22, 8),
48416 => conv_std_logic_vector(23, 8),
48417 => conv_std_logic_vector(24, 8),
48418 => conv_std_logic_vector(25, 8),
48419 => conv_std_logic_vector(25, 8),
48420 => conv_std_logic_vector(26, 8),
48421 => conv_std_logic_vector(27, 8),
48422 => conv_std_logic_vector(28, 8),
48423 => conv_std_logic_vector(28, 8),
48424 => conv_std_logic_vector(29, 8),
48425 => conv_std_logic_vector(30, 8),
48426 => conv_std_logic_vector(31, 8),
48427 => conv_std_logic_vector(31, 8),
48428 => conv_std_logic_vector(32, 8),
48429 => conv_std_logic_vector(33, 8),
48430 => conv_std_logic_vector(33, 8),
48431 => conv_std_logic_vector(34, 8),
48432 => conv_std_logic_vector(35, 8),
48433 => conv_std_logic_vector(36, 8),
48434 => conv_std_logic_vector(36, 8),
48435 => conv_std_logic_vector(37, 8),
48436 => conv_std_logic_vector(38, 8),
48437 => conv_std_logic_vector(39, 8),
48438 => conv_std_logic_vector(39, 8),
48439 => conv_std_logic_vector(40, 8),
48440 => conv_std_logic_vector(41, 8),
48441 => conv_std_logic_vector(42, 8),
48442 => conv_std_logic_vector(42, 8),
48443 => conv_std_logic_vector(43, 8),
48444 => conv_std_logic_vector(44, 8),
48445 => conv_std_logic_vector(45, 8),
48446 => conv_std_logic_vector(45, 8),
48447 => conv_std_logic_vector(46, 8),
48448 => conv_std_logic_vector(47, 8),
48449 => conv_std_logic_vector(47, 8),
48450 => conv_std_logic_vector(48, 8),
48451 => conv_std_logic_vector(49, 8),
48452 => conv_std_logic_vector(50, 8),
48453 => conv_std_logic_vector(50, 8),
48454 => conv_std_logic_vector(51, 8),
48455 => conv_std_logic_vector(52, 8),
48456 => conv_std_logic_vector(53, 8),
48457 => conv_std_logic_vector(53, 8),
48458 => conv_std_logic_vector(54, 8),
48459 => conv_std_logic_vector(55, 8),
48460 => conv_std_logic_vector(56, 8),
48461 => conv_std_logic_vector(56, 8),
48462 => conv_std_logic_vector(57, 8),
48463 => conv_std_logic_vector(58, 8),
48464 => conv_std_logic_vector(59, 8),
48465 => conv_std_logic_vector(59, 8),
48466 => conv_std_logic_vector(60, 8),
48467 => conv_std_logic_vector(61, 8),
48468 => conv_std_logic_vector(62, 8),
48469 => conv_std_logic_vector(62, 8),
48470 => conv_std_logic_vector(63, 8),
48471 => conv_std_logic_vector(64, 8),
48472 => conv_std_logic_vector(64, 8),
48473 => conv_std_logic_vector(65, 8),
48474 => conv_std_logic_vector(66, 8),
48475 => conv_std_logic_vector(67, 8),
48476 => conv_std_logic_vector(67, 8),
48477 => conv_std_logic_vector(68, 8),
48478 => conv_std_logic_vector(69, 8),
48479 => conv_std_logic_vector(70, 8),
48480 => conv_std_logic_vector(70, 8),
48481 => conv_std_logic_vector(71, 8),
48482 => conv_std_logic_vector(72, 8),
48483 => conv_std_logic_vector(73, 8),
48484 => conv_std_logic_vector(73, 8),
48485 => conv_std_logic_vector(74, 8),
48486 => conv_std_logic_vector(75, 8),
48487 => conv_std_logic_vector(76, 8),
48488 => conv_std_logic_vector(76, 8),
48489 => conv_std_logic_vector(77, 8),
48490 => conv_std_logic_vector(78, 8),
48491 => conv_std_logic_vector(78, 8),
48492 => conv_std_logic_vector(79, 8),
48493 => conv_std_logic_vector(80, 8),
48494 => conv_std_logic_vector(81, 8),
48495 => conv_std_logic_vector(81, 8),
48496 => conv_std_logic_vector(82, 8),
48497 => conv_std_logic_vector(83, 8),
48498 => conv_std_logic_vector(84, 8),
48499 => conv_std_logic_vector(84, 8),
48500 => conv_std_logic_vector(85, 8),
48501 => conv_std_logic_vector(86, 8),
48502 => conv_std_logic_vector(87, 8),
48503 => conv_std_logic_vector(87, 8),
48504 => conv_std_logic_vector(88, 8),
48505 => conv_std_logic_vector(89, 8),
48506 => conv_std_logic_vector(90, 8),
48507 => conv_std_logic_vector(90, 8),
48508 => conv_std_logic_vector(91, 8),
48509 => conv_std_logic_vector(92, 8),
48510 => conv_std_logic_vector(93, 8),
48511 => conv_std_logic_vector(93, 8),
48512 => conv_std_logic_vector(94, 8),
48513 => conv_std_logic_vector(95, 8),
48514 => conv_std_logic_vector(95, 8),
48515 => conv_std_logic_vector(96, 8),
48516 => conv_std_logic_vector(97, 8),
48517 => conv_std_logic_vector(98, 8),
48518 => conv_std_logic_vector(98, 8),
48519 => conv_std_logic_vector(99, 8),
48520 => conv_std_logic_vector(100, 8),
48521 => conv_std_logic_vector(101, 8),
48522 => conv_std_logic_vector(101, 8),
48523 => conv_std_logic_vector(102, 8),
48524 => conv_std_logic_vector(103, 8),
48525 => conv_std_logic_vector(104, 8),
48526 => conv_std_logic_vector(104, 8),
48527 => conv_std_logic_vector(105, 8),
48528 => conv_std_logic_vector(106, 8),
48529 => conv_std_logic_vector(107, 8),
48530 => conv_std_logic_vector(107, 8),
48531 => conv_std_logic_vector(108, 8),
48532 => conv_std_logic_vector(109, 8),
48533 => conv_std_logic_vector(110, 8),
48534 => conv_std_logic_vector(110, 8),
48535 => conv_std_logic_vector(111, 8),
48536 => conv_std_logic_vector(112, 8),
48537 => conv_std_logic_vector(112, 8),
48538 => conv_std_logic_vector(113, 8),
48539 => conv_std_logic_vector(114, 8),
48540 => conv_std_logic_vector(115, 8),
48541 => conv_std_logic_vector(115, 8),
48542 => conv_std_logic_vector(116, 8),
48543 => conv_std_logic_vector(117, 8),
48544 => conv_std_logic_vector(118, 8),
48545 => conv_std_logic_vector(118, 8),
48546 => conv_std_logic_vector(119, 8),
48547 => conv_std_logic_vector(120, 8),
48548 => conv_std_logic_vector(121, 8),
48549 => conv_std_logic_vector(121, 8),
48550 => conv_std_logic_vector(122, 8),
48551 => conv_std_logic_vector(123, 8),
48552 => conv_std_logic_vector(124, 8),
48553 => conv_std_logic_vector(124, 8),
48554 => conv_std_logic_vector(125, 8),
48555 => conv_std_logic_vector(126, 8),
48556 => conv_std_logic_vector(126, 8),
48557 => conv_std_logic_vector(127, 8),
48558 => conv_std_logic_vector(128, 8),
48559 => conv_std_logic_vector(129, 8),
48560 => conv_std_logic_vector(129, 8),
48561 => conv_std_logic_vector(130, 8),
48562 => conv_std_logic_vector(131, 8),
48563 => conv_std_logic_vector(132, 8),
48564 => conv_std_logic_vector(132, 8),
48565 => conv_std_logic_vector(133, 8),
48566 => conv_std_logic_vector(134, 8),
48567 => conv_std_logic_vector(135, 8),
48568 => conv_std_logic_vector(135, 8),
48569 => conv_std_logic_vector(136, 8),
48570 => conv_std_logic_vector(137, 8),
48571 => conv_std_logic_vector(138, 8),
48572 => conv_std_logic_vector(138, 8),
48573 => conv_std_logic_vector(139, 8),
48574 => conv_std_logic_vector(140, 8),
48575 => conv_std_logic_vector(141, 8),
48576 => conv_std_logic_vector(141, 8),
48577 => conv_std_logic_vector(142, 8),
48578 => conv_std_logic_vector(143, 8),
48579 => conv_std_logic_vector(143, 8),
48580 => conv_std_logic_vector(144, 8),
48581 => conv_std_logic_vector(145, 8),
48582 => conv_std_logic_vector(146, 8),
48583 => conv_std_logic_vector(146, 8),
48584 => conv_std_logic_vector(147, 8),
48585 => conv_std_logic_vector(148, 8),
48586 => conv_std_logic_vector(149, 8),
48587 => conv_std_logic_vector(149, 8),
48588 => conv_std_logic_vector(150, 8),
48589 => conv_std_logic_vector(151, 8),
48590 => conv_std_logic_vector(152, 8),
48591 => conv_std_logic_vector(152, 8),
48592 => conv_std_logic_vector(153, 8),
48593 => conv_std_logic_vector(154, 8),
48594 => conv_std_logic_vector(155, 8),
48595 => conv_std_logic_vector(155, 8),
48596 => conv_std_logic_vector(156, 8),
48597 => conv_std_logic_vector(157, 8),
48598 => conv_std_logic_vector(157, 8),
48599 => conv_std_logic_vector(158, 8),
48600 => conv_std_logic_vector(159, 8),
48601 => conv_std_logic_vector(160, 8),
48602 => conv_std_logic_vector(160, 8),
48603 => conv_std_logic_vector(161, 8),
48604 => conv_std_logic_vector(162, 8),
48605 => conv_std_logic_vector(163, 8),
48606 => conv_std_logic_vector(163, 8),
48607 => conv_std_logic_vector(164, 8),
48608 => conv_std_logic_vector(165, 8),
48609 => conv_std_logic_vector(166, 8),
48610 => conv_std_logic_vector(166, 8),
48611 => conv_std_logic_vector(167, 8),
48612 => conv_std_logic_vector(168, 8),
48613 => conv_std_logic_vector(169, 8),
48614 => conv_std_logic_vector(169, 8),
48615 => conv_std_logic_vector(170, 8),
48616 => conv_std_logic_vector(171, 8),
48617 => conv_std_logic_vector(172, 8),
48618 => conv_std_logic_vector(172, 8),
48619 => conv_std_logic_vector(173, 8),
48620 => conv_std_logic_vector(174, 8),
48621 => conv_std_logic_vector(174, 8),
48622 => conv_std_logic_vector(175, 8),
48623 => conv_std_logic_vector(176, 8),
48624 => conv_std_logic_vector(177, 8),
48625 => conv_std_logic_vector(177, 8),
48626 => conv_std_logic_vector(178, 8),
48627 => conv_std_logic_vector(179, 8),
48628 => conv_std_logic_vector(180, 8),
48629 => conv_std_logic_vector(180, 8),
48630 => conv_std_logic_vector(181, 8),
48631 => conv_std_logic_vector(182, 8),
48632 => conv_std_logic_vector(183, 8),
48633 => conv_std_logic_vector(183, 8),
48634 => conv_std_logic_vector(184, 8),
48635 => conv_std_logic_vector(185, 8),
48636 => conv_std_logic_vector(186, 8),
48637 => conv_std_logic_vector(186, 8),
48638 => conv_std_logic_vector(187, 8),
48639 => conv_std_logic_vector(188, 8),
48640 => conv_std_logic_vector(0, 8),
48641 => conv_std_logic_vector(0, 8),
48642 => conv_std_logic_vector(1, 8),
48643 => conv_std_logic_vector(2, 8),
48644 => conv_std_logic_vector(2, 8),
48645 => conv_std_logic_vector(3, 8),
48646 => conv_std_logic_vector(4, 8),
48647 => conv_std_logic_vector(5, 8),
48648 => conv_std_logic_vector(5, 8),
48649 => conv_std_logic_vector(6, 8),
48650 => conv_std_logic_vector(7, 8),
48651 => conv_std_logic_vector(8, 8),
48652 => conv_std_logic_vector(8, 8),
48653 => conv_std_logic_vector(9, 8),
48654 => conv_std_logic_vector(10, 8),
48655 => conv_std_logic_vector(11, 8),
48656 => conv_std_logic_vector(11, 8),
48657 => conv_std_logic_vector(12, 8),
48658 => conv_std_logic_vector(13, 8),
48659 => conv_std_logic_vector(14, 8),
48660 => conv_std_logic_vector(14, 8),
48661 => conv_std_logic_vector(15, 8),
48662 => conv_std_logic_vector(16, 8),
48663 => conv_std_logic_vector(17, 8),
48664 => conv_std_logic_vector(17, 8),
48665 => conv_std_logic_vector(18, 8),
48666 => conv_std_logic_vector(19, 8),
48667 => conv_std_logic_vector(20, 8),
48668 => conv_std_logic_vector(20, 8),
48669 => conv_std_logic_vector(21, 8),
48670 => conv_std_logic_vector(22, 8),
48671 => conv_std_logic_vector(23, 8),
48672 => conv_std_logic_vector(23, 8),
48673 => conv_std_logic_vector(24, 8),
48674 => conv_std_logic_vector(25, 8),
48675 => conv_std_logic_vector(25, 8),
48676 => conv_std_logic_vector(26, 8),
48677 => conv_std_logic_vector(27, 8),
48678 => conv_std_logic_vector(28, 8),
48679 => conv_std_logic_vector(28, 8),
48680 => conv_std_logic_vector(29, 8),
48681 => conv_std_logic_vector(30, 8),
48682 => conv_std_logic_vector(31, 8),
48683 => conv_std_logic_vector(31, 8),
48684 => conv_std_logic_vector(32, 8),
48685 => conv_std_logic_vector(33, 8),
48686 => conv_std_logic_vector(34, 8),
48687 => conv_std_logic_vector(34, 8),
48688 => conv_std_logic_vector(35, 8),
48689 => conv_std_logic_vector(36, 8),
48690 => conv_std_logic_vector(37, 8),
48691 => conv_std_logic_vector(37, 8),
48692 => conv_std_logic_vector(38, 8),
48693 => conv_std_logic_vector(39, 8),
48694 => conv_std_logic_vector(40, 8),
48695 => conv_std_logic_vector(40, 8),
48696 => conv_std_logic_vector(41, 8),
48697 => conv_std_logic_vector(42, 8),
48698 => conv_std_logic_vector(43, 8),
48699 => conv_std_logic_vector(43, 8),
48700 => conv_std_logic_vector(44, 8),
48701 => conv_std_logic_vector(45, 8),
48702 => conv_std_logic_vector(46, 8),
48703 => conv_std_logic_vector(46, 8),
48704 => conv_std_logic_vector(47, 8),
48705 => conv_std_logic_vector(48, 8),
48706 => conv_std_logic_vector(48, 8),
48707 => conv_std_logic_vector(49, 8),
48708 => conv_std_logic_vector(50, 8),
48709 => conv_std_logic_vector(51, 8),
48710 => conv_std_logic_vector(51, 8),
48711 => conv_std_logic_vector(52, 8),
48712 => conv_std_logic_vector(53, 8),
48713 => conv_std_logic_vector(54, 8),
48714 => conv_std_logic_vector(54, 8),
48715 => conv_std_logic_vector(55, 8),
48716 => conv_std_logic_vector(56, 8),
48717 => conv_std_logic_vector(57, 8),
48718 => conv_std_logic_vector(57, 8),
48719 => conv_std_logic_vector(58, 8),
48720 => conv_std_logic_vector(59, 8),
48721 => conv_std_logic_vector(60, 8),
48722 => conv_std_logic_vector(60, 8),
48723 => conv_std_logic_vector(61, 8),
48724 => conv_std_logic_vector(62, 8),
48725 => conv_std_logic_vector(63, 8),
48726 => conv_std_logic_vector(63, 8),
48727 => conv_std_logic_vector(64, 8),
48728 => conv_std_logic_vector(65, 8),
48729 => conv_std_logic_vector(66, 8),
48730 => conv_std_logic_vector(66, 8),
48731 => conv_std_logic_vector(67, 8),
48732 => conv_std_logic_vector(68, 8),
48733 => conv_std_logic_vector(69, 8),
48734 => conv_std_logic_vector(69, 8),
48735 => conv_std_logic_vector(70, 8),
48736 => conv_std_logic_vector(71, 8),
48737 => conv_std_logic_vector(71, 8),
48738 => conv_std_logic_vector(72, 8),
48739 => conv_std_logic_vector(73, 8),
48740 => conv_std_logic_vector(74, 8),
48741 => conv_std_logic_vector(74, 8),
48742 => conv_std_logic_vector(75, 8),
48743 => conv_std_logic_vector(76, 8),
48744 => conv_std_logic_vector(77, 8),
48745 => conv_std_logic_vector(77, 8),
48746 => conv_std_logic_vector(78, 8),
48747 => conv_std_logic_vector(79, 8),
48748 => conv_std_logic_vector(80, 8),
48749 => conv_std_logic_vector(80, 8),
48750 => conv_std_logic_vector(81, 8),
48751 => conv_std_logic_vector(82, 8),
48752 => conv_std_logic_vector(83, 8),
48753 => conv_std_logic_vector(83, 8),
48754 => conv_std_logic_vector(84, 8),
48755 => conv_std_logic_vector(85, 8),
48756 => conv_std_logic_vector(86, 8),
48757 => conv_std_logic_vector(86, 8),
48758 => conv_std_logic_vector(87, 8),
48759 => conv_std_logic_vector(88, 8),
48760 => conv_std_logic_vector(89, 8),
48761 => conv_std_logic_vector(89, 8),
48762 => conv_std_logic_vector(90, 8),
48763 => conv_std_logic_vector(91, 8),
48764 => conv_std_logic_vector(92, 8),
48765 => conv_std_logic_vector(92, 8),
48766 => conv_std_logic_vector(93, 8),
48767 => conv_std_logic_vector(94, 8),
48768 => conv_std_logic_vector(95, 8),
48769 => conv_std_logic_vector(95, 8),
48770 => conv_std_logic_vector(96, 8),
48771 => conv_std_logic_vector(97, 8),
48772 => conv_std_logic_vector(97, 8),
48773 => conv_std_logic_vector(98, 8),
48774 => conv_std_logic_vector(99, 8),
48775 => conv_std_logic_vector(100, 8),
48776 => conv_std_logic_vector(100, 8),
48777 => conv_std_logic_vector(101, 8),
48778 => conv_std_logic_vector(102, 8),
48779 => conv_std_logic_vector(103, 8),
48780 => conv_std_logic_vector(103, 8),
48781 => conv_std_logic_vector(104, 8),
48782 => conv_std_logic_vector(105, 8),
48783 => conv_std_logic_vector(106, 8),
48784 => conv_std_logic_vector(106, 8),
48785 => conv_std_logic_vector(107, 8),
48786 => conv_std_logic_vector(108, 8),
48787 => conv_std_logic_vector(109, 8),
48788 => conv_std_logic_vector(109, 8),
48789 => conv_std_logic_vector(110, 8),
48790 => conv_std_logic_vector(111, 8),
48791 => conv_std_logic_vector(112, 8),
48792 => conv_std_logic_vector(112, 8),
48793 => conv_std_logic_vector(113, 8),
48794 => conv_std_logic_vector(114, 8),
48795 => conv_std_logic_vector(115, 8),
48796 => conv_std_logic_vector(115, 8),
48797 => conv_std_logic_vector(116, 8),
48798 => conv_std_logic_vector(117, 8),
48799 => conv_std_logic_vector(118, 8),
48800 => conv_std_logic_vector(118, 8),
48801 => conv_std_logic_vector(119, 8),
48802 => conv_std_logic_vector(120, 8),
48803 => conv_std_logic_vector(120, 8),
48804 => conv_std_logic_vector(121, 8),
48805 => conv_std_logic_vector(122, 8),
48806 => conv_std_logic_vector(123, 8),
48807 => conv_std_logic_vector(123, 8),
48808 => conv_std_logic_vector(124, 8),
48809 => conv_std_logic_vector(125, 8),
48810 => conv_std_logic_vector(126, 8),
48811 => conv_std_logic_vector(126, 8),
48812 => conv_std_logic_vector(127, 8),
48813 => conv_std_logic_vector(128, 8),
48814 => conv_std_logic_vector(129, 8),
48815 => conv_std_logic_vector(129, 8),
48816 => conv_std_logic_vector(130, 8),
48817 => conv_std_logic_vector(131, 8),
48818 => conv_std_logic_vector(132, 8),
48819 => conv_std_logic_vector(132, 8),
48820 => conv_std_logic_vector(133, 8),
48821 => conv_std_logic_vector(134, 8),
48822 => conv_std_logic_vector(135, 8),
48823 => conv_std_logic_vector(135, 8),
48824 => conv_std_logic_vector(136, 8),
48825 => conv_std_logic_vector(137, 8),
48826 => conv_std_logic_vector(138, 8),
48827 => conv_std_logic_vector(138, 8),
48828 => conv_std_logic_vector(139, 8),
48829 => conv_std_logic_vector(140, 8),
48830 => conv_std_logic_vector(141, 8),
48831 => conv_std_logic_vector(141, 8),
48832 => conv_std_logic_vector(142, 8),
48833 => conv_std_logic_vector(143, 8),
48834 => conv_std_logic_vector(143, 8),
48835 => conv_std_logic_vector(144, 8),
48836 => conv_std_logic_vector(145, 8),
48837 => conv_std_logic_vector(146, 8),
48838 => conv_std_logic_vector(146, 8),
48839 => conv_std_logic_vector(147, 8),
48840 => conv_std_logic_vector(148, 8),
48841 => conv_std_logic_vector(149, 8),
48842 => conv_std_logic_vector(149, 8),
48843 => conv_std_logic_vector(150, 8),
48844 => conv_std_logic_vector(151, 8),
48845 => conv_std_logic_vector(152, 8),
48846 => conv_std_logic_vector(152, 8),
48847 => conv_std_logic_vector(153, 8),
48848 => conv_std_logic_vector(154, 8),
48849 => conv_std_logic_vector(155, 8),
48850 => conv_std_logic_vector(155, 8),
48851 => conv_std_logic_vector(156, 8),
48852 => conv_std_logic_vector(157, 8),
48853 => conv_std_logic_vector(158, 8),
48854 => conv_std_logic_vector(158, 8),
48855 => conv_std_logic_vector(159, 8),
48856 => conv_std_logic_vector(160, 8),
48857 => conv_std_logic_vector(161, 8),
48858 => conv_std_logic_vector(161, 8),
48859 => conv_std_logic_vector(162, 8),
48860 => conv_std_logic_vector(163, 8),
48861 => conv_std_logic_vector(164, 8),
48862 => conv_std_logic_vector(164, 8),
48863 => conv_std_logic_vector(165, 8),
48864 => conv_std_logic_vector(166, 8),
48865 => conv_std_logic_vector(166, 8),
48866 => conv_std_logic_vector(167, 8),
48867 => conv_std_logic_vector(168, 8),
48868 => conv_std_logic_vector(169, 8),
48869 => conv_std_logic_vector(169, 8),
48870 => conv_std_logic_vector(170, 8),
48871 => conv_std_logic_vector(171, 8),
48872 => conv_std_logic_vector(172, 8),
48873 => conv_std_logic_vector(172, 8),
48874 => conv_std_logic_vector(173, 8),
48875 => conv_std_logic_vector(174, 8),
48876 => conv_std_logic_vector(175, 8),
48877 => conv_std_logic_vector(175, 8),
48878 => conv_std_logic_vector(176, 8),
48879 => conv_std_logic_vector(177, 8),
48880 => conv_std_logic_vector(178, 8),
48881 => conv_std_logic_vector(178, 8),
48882 => conv_std_logic_vector(179, 8),
48883 => conv_std_logic_vector(180, 8),
48884 => conv_std_logic_vector(181, 8),
48885 => conv_std_logic_vector(181, 8),
48886 => conv_std_logic_vector(182, 8),
48887 => conv_std_logic_vector(183, 8),
48888 => conv_std_logic_vector(184, 8),
48889 => conv_std_logic_vector(184, 8),
48890 => conv_std_logic_vector(185, 8),
48891 => conv_std_logic_vector(186, 8),
48892 => conv_std_logic_vector(187, 8),
48893 => conv_std_logic_vector(187, 8),
48894 => conv_std_logic_vector(188, 8),
48895 => conv_std_logic_vector(189, 8),
48896 => conv_std_logic_vector(0, 8),
48897 => conv_std_logic_vector(0, 8),
48898 => conv_std_logic_vector(1, 8),
48899 => conv_std_logic_vector(2, 8),
48900 => conv_std_logic_vector(2, 8),
48901 => conv_std_logic_vector(3, 8),
48902 => conv_std_logic_vector(4, 8),
48903 => conv_std_logic_vector(5, 8),
48904 => conv_std_logic_vector(5, 8),
48905 => conv_std_logic_vector(6, 8),
48906 => conv_std_logic_vector(7, 8),
48907 => conv_std_logic_vector(8, 8),
48908 => conv_std_logic_vector(8, 8),
48909 => conv_std_logic_vector(9, 8),
48910 => conv_std_logic_vector(10, 8),
48911 => conv_std_logic_vector(11, 8),
48912 => conv_std_logic_vector(11, 8),
48913 => conv_std_logic_vector(12, 8),
48914 => conv_std_logic_vector(13, 8),
48915 => conv_std_logic_vector(14, 8),
48916 => conv_std_logic_vector(14, 8),
48917 => conv_std_logic_vector(15, 8),
48918 => conv_std_logic_vector(16, 8),
48919 => conv_std_logic_vector(17, 8),
48920 => conv_std_logic_vector(17, 8),
48921 => conv_std_logic_vector(18, 8),
48922 => conv_std_logic_vector(19, 8),
48923 => conv_std_logic_vector(20, 8),
48924 => conv_std_logic_vector(20, 8),
48925 => conv_std_logic_vector(21, 8),
48926 => conv_std_logic_vector(22, 8),
48927 => conv_std_logic_vector(23, 8),
48928 => conv_std_logic_vector(23, 8),
48929 => conv_std_logic_vector(24, 8),
48930 => conv_std_logic_vector(25, 8),
48931 => conv_std_logic_vector(26, 8),
48932 => conv_std_logic_vector(26, 8),
48933 => conv_std_logic_vector(27, 8),
48934 => conv_std_logic_vector(28, 8),
48935 => conv_std_logic_vector(29, 8),
48936 => conv_std_logic_vector(29, 8),
48937 => conv_std_logic_vector(30, 8),
48938 => conv_std_logic_vector(31, 8),
48939 => conv_std_logic_vector(32, 8),
48940 => conv_std_logic_vector(32, 8),
48941 => conv_std_logic_vector(33, 8),
48942 => conv_std_logic_vector(34, 8),
48943 => conv_std_logic_vector(35, 8),
48944 => conv_std_logic_vector(35, 8),
48945 => conv_std_logic_vector(36, 8),
48946 => conv_std_logic_vector(37, 8),
48947 => conv_std_logic_vector(38, 8),
48948 => conv_std_logic_vector(38, 8),
48949 => conv_std_logic_vector(39, 8),
48950 => conv_std_logic_vector(40, 8),
48951 => conv_std_logic_vector(41, 8),
48952 => conv_std_logic_vector(41, 8),
48953 => conv_std_logic_vector(42, 8),
48954 => conv_std_logic_vector(43, 8),
48955 => conv_std_logic_vector(44, 8),
48956 => conv_std_logic_vector(44, 8),
48957 => conv_std_logic_vector(45, 8),
48958 => conv_std_logic_vector(46, 8),
48959 => conv_std_logic_vector(47, 8),
48960 => conv_std_logic_vector(47, 8),
48961 => conv_std_logic_vector(48, 8),
48962 => conv_std_logic_vector(49, 8),
48963 => conv_std_logic_vector(49, 8),
48964 => conv_std_logic_vector(50, 8),
48965 => conv_std_logic_vector(51, 8),
48966 => conv_std_logic_vector(52, 8),
48967 => conv_std_logic_vector(52, 8),
48968 => conv_std_logic_vector(53, 8),
48969 => conv_std_logic_vector(54, 8),
48970 => conv_std_logic_vector(55, 8),
48971 => conv_std_logic_vector(55, 8),
48972 => conv_std_logic_vector(56, 8),
48973 => conv_std_logic_vector(57, 8),
48974 => conv_std_logic_vector(58, 8),
48975 => conv_std_logic_vector(58, 8),
48976 => conv_std_logic_vector(59, 8),
48977 => conv_std_logic_vector(60, 8),
48978 => conv_std_logic_vector(61, 8),
48979 => conv_std_logic_vector(61, 8),
48980 => conv_std_logic_vector(62, 8),
48981 => conv_std_logic_vector(63, 8),
48982 => conv_std_logic_vector(64, 8),
48983 => conv_std_logic_vector(64, 8),
48984 => conv_std_logic_vector(65, 8),
48985 => conv_std_logic_vector(66, 8),
48986 => conv_std_logic_vector(67, 8),
48987 => conv_std_logic_vector(67, 8),
48988 => conv_std_logic_vector(68, 8),
48989 => conv_std_logic_vector(69, 8),
48990 => conv_std_logic_vector(70, 8),
48991 => conv_std_logic_vector(70, 8),
48992 => conv_std_logic_vector(71, 8),
48993 => conv_std_logic_vector(72, 8),
48994 => conv_std_logic_vector(73, 8),
48995 => conv_std_logic_vector(73, 8),
48996 => conv_std_logic_vector(74, 8),
48997 => conv_std_logic_vector(75, 8),
48998 => conv_std_logic_vector(76, 8),
48999 => conv_std_logic_vector(76, 8),
49000 => conv_std_logic_vector(77, 8),
49001 => conv_std_logic_vector(78, 8),
49002 => conv_std_logic_vector(79, 8),
49003 => conv_std_logic_vector(79, 8),
49004 => conv_std_logic_vector(80, 8),
49005 => conv_std_logic_vector(81, 8),
49006 => conv_std_logic_vector(82, 8),
49007 => conv_std_logic_vector(82, 8),
49008 => conv_std_logic_vector(83, 8),
49009 => conv_std_logic_vector(84, 8),
49010 => conv_std_logic_vector(85, 8),
49011 => conv_std_logic_vector(85, 8),
49012 => conv_std_logic_vector(86, 8),
49013 => conv_std_logic_vector(87, 8),
49014 => conv_std_logic_vector(88, 8),
49015 => conv_std_logic_vector(88, 8),
49016 => conv_std_logic_vector(89, 8),
49017 => conv_std_logic_vector(90, 8),
49018 => conv_std_logic_vector(91, 8),
49019 => conv_std_logic_vector(91, 8),
49020 => conv_std_logic_vector(92, 8),
49021 => conv_std_logic_vector(93, 8),
49022 => conv_std_logic_vector(94, 8),
49023 => conv_std_logic_vector(94, 8),
49024 => conv_std_logic_vector(95, 8),
49025 => conv_std_logic_vector(96, 8),
49026 => conv_std_logic_vector(96, 8),
49027 => conv_std_logic_vector(97, 8),
49028 => conv_std_logic_vector(98, 8),
49029 => conv_std_logic_vector(99, 8),
49030 => conv_std_logic_vector(99, 8),
49031 => conv_std_logic_vector(100, 8),
49032 => conv_std_logic_vector(101, 8),
49033 => conv_std_logic_vector(102, 8),
49034 => conv_std_logic_vector(102, 8),
49035 => conv_std_logic_vector(103, 8),
49036 => conv_std_logic_vector(104, 8),
49037 => conv_std_logic_vector(105, 8),
49038 => conv_std_logic_vector(105, 8),
49039 => conv_std_logic_vector(106, 8),
49040 => conv_std_logic_vector(107, 8),
49041 => conv_std_logic_vector(108, 8),
49042 => conv_std_logic_vector(108, 8),
49043 => conv_std_logic_vector(109, 8),
49044 => conv_std_logic_vector(110, 8),
49045 => conv_std_logic_vector(111, 8),
49046 => conv_std_logic_vector(111, 8),
49047 => conv_std_logic_vector(112, 8),
49048 => conv_std_logic_vector(113, 8),
49049 => conv_std_logic_vector(114, 8),
49050 => conv_std_logic_vector(114, 8),
49051 => conv_std_logic_vector(115, 8),
49052 => conv_std_logic_vector(116, 8),
49053 => conv_std_logic_vector(117, 8),
49054 => conv_std_logic_vector(117, 8),
49055 => conv_std_logic_vector(118, 8),
49056 => conv_std_logic_vector(119, 8),
49057 => conv_std_logic_vector(120, 8),
49058 => conv_std_logic_vector(120, 8),
49059 => conv_std_logic_vector(121, 8),
49060 => conv_std_logic_vector(122, 8),
49061 => conv_std_logic_vector(123, 8),
49062 => conv_std_logic_vector(123, 8),
49063 => conv_std_logic_vector(124, 8),
49064 => conv_std_logic_vector(125, 8),
49065 => conv_std_logic_vector(126, 8),
49066 => conv_std_logic_vector(126, 8),
49067 => conv_std_logic_vector(127, 8),
49068 => conv_std_logic_vector(128, 8),
49069 => conv_std_logic_vector(129, 8),
49070 => conv_std_logic_vector(129, 8),
49071 => conv_std_logic_vector(130, 8),
49072 => conv_std_logic_vector(131, 8),
49073 => conv_std_logic_vector(132, 8),
49074 => conv_std_logic_vector(132, 8),
49075 => conv_std_logic_vector(133, 8),
49076 => conv_std_logic_vector(134, 8),
49077 => conv_std_logic_vector(135, 8),
49078 => conv_std_logic_vector(135, 8),
49079 => conv_std_logic_vector(136, 8),
49080 => conv_std_logic_vector(137, 8),
49081 => conv_std_logic_vector(138, 8),
49082 => conv_std_logic_vector(138, 8),
49083 => conv_std_logic_vector(139, 8),
49084 => conv_std_logic_vector(140, 8),
49085 => conv_std_logic_vector(141, 8),
49086 => conv_std_logic_vector(141, 8),
49087 => conv_std_logic_vector(142, 8),
49088 => conv_std_logic_vector(143, 8),
49089 => conv_std_logic_vector(143, 8),
49090 => conv_std_logic_vector(144, 8),
49091 => conv_std_logic_vector(145, 8),
49092 => conv_std_logic_vector(146, 8),
49093 => conv_std_logic_vector(146, 8),
49094 => conv_std_logic_vector(147, 8),
49095 => conv_std_logic_vector(148, 8),
49096 => conv_std_logic_vector(149, 8),
49097 => conv_std_logic_vector(149, 8),
49098 => conv_std_logic_vector(150, 8),
49099 => conv_std_logic_vector(151, 8),
49100 => conv_std_logic_vector(152, 8),
49101 => conv_std_logic_vector(152, 8),
49102 => conv_std_logic_vector(153, 8),
49103 => conv_std_logic_vector(154, 8),
49104 => conv_std_logic_vector(155, 8),
49105 => conv_std_logic_vector(155, 8),
49106 => conv_std_logic_vector(156, 8),
49107 => conv_std_logic_vector(157, 8),
49108 => conv_std_logic_vector(158, 8),
49109 => conv_std_logic_vector(158, 8),
49110 => conv_std_logic_vector(159, 8),
49111 => conv_std_logic_vector(160, 8),
49112 => conv_std_logic_vector(161, 8),
49113 => conv_std_logic_vector(161, 8),
49114 => conv_std_logic_vector(162, 8),
49115 => conv_std_logic_vector(163, 8),
49116 => conv_std_logic_vector(164, 8),
49117 => conv_std_logic_vector(164, 8),
49118 => conv_std_logic_vector(165, 8),
49119 => conv_std_logic_vector(166, 8),
49120 => conv_std_logic_vector(167, 8),
49121 => conv_std_logic_vector(167, 8),
49122 => conv_std_logic_vector(168, 8),
49123 => conv_std_logic_vector(169, 8),
49124 => conv_std_logic_vector(170, 8),
49125 => conv_std_logic_vector(170, 8),
49126 => conv_std_logic_vector(171, 8),
49127 => conv_std_logic_vector(172, 8),
49128 => conv_std_logic_vector(173, 8),
49129 => conv_std_logic_vector(173, 8),
49130 => conv_std_logic_vector(174, 8),
49131 => conv_std_logic_vector(175, 8),
49132 => conv_std_logic_vector(176, 8),
49133 => conv_std_logic_vector(176, 8),
49134 => conv_std_logic_vector(177, 8),
49135 => conv_std_logic_vector(178, 8),
49136 => conv_std_logic_vector(179, 8),
49137 => conv_std_logic_vector(179, 8),
49138 => conv_std_logic_vector(180, 8),
49139 => conv_std_logic_vector(181, 8),
49140 => conv_std_logic_vector(182, 8),
49141 => conv_std_logic_vector(182, 8),
49142 => conv_std_logic_vector(183, 8),
49143 => conv_std_logic_vector(184, 8),
49144 => conv_std_logic_vector(185, 8),
49145 => conv_std_logic_vector(185, 8),
49146 => conv_std_logic_vector(186, 8),
49147 => conv_std_logic_vector(187, 8),
49148 => conv_std_logic_vector(188, 8),
49149 => conv_std_logic_vector(188, 8),
49150 => conv_std_logic_vector(189, 8),
49151 => conv_std_logic_vector(190, 8),
49152 => conv_std_logic_vector(0, 8),
49153 => conv_std_logic_vector(0, 8),
49154 => conv_std_logic_vector(1, 8),
49155 => conv_std_logic_vector(2, 8),
49156 => conv_std_logic_vector(3, 8),
49157 => conv_std_logic_vector(3, 8),
49158 => conv_std_logic_vector(4, 8),
49159 => conv_std_logic_vector(5, 8),
49160 => conv_std_logic_vector(6, 8),
49161 => conv_std_logic_vector(6, 8),
49162 => conv_std_logic_vector(7, 8),
49163 => conv_std_logic_vector(8, 8),
49164 => conv_std_logic_vector(9, 8),
49165 => conv_std_logic_vector(9, 8),
49166 => conv_std_logic_vector(10, 8),
49167 => conv_std_logic_vector(11, 8),
49168 => conv_std_logic_vector(12, 8),
49169 => conv_std_logic_vector(12, 8),
49170 => conv_std_logic_vector(13, 8),
49171 => conv_std_logic_vector(14, 8),
49172 => conv_std_logic_vector(15, 8),
49173 => conv_std_logic_vector(15, 8),
49174 => conv_std_logic_vector(16, 8),
49175 => conv_std_logic_vector(17, 8),
49176 => conv_std_logic_vector(18, 8),
49177 => conv_std_logic_vector(18, 8),
49178 => conv_std_logic_vector(19, 8),
49179 => conv_std_logic_vector(20, 8),
49180 => conv_std_logic_vector(21, 8),
49181 => conv_std_logic_vector(21, 8),
49182 => conv_std_logic_vector(22, 8),
49183 => conv_std_logic_vector(23, 8),
49184 => conv_std_logic_vector(24, 8),
49185 => conv_std_logic_vector(24, 8),
49186 => conv_std_logic_vector(25, 8),
49187 => conv_std_logic_vector(26, 8),
49188 => conv_std_logic_vector(27, 8),
49189 => conv_std_logic_vector(27, 8),
49190 => conv_std_logic_vector(28, 8),
49191 => conv_std_logic_vector(29, 8),
49192 => conv_std_logic_vector(30, 8),
49193 => conv_std_logic_vector(30, 8),
49194 => conv_std_logic_vector(31, 8),
49195 => conv_std_logic_vector(32, 8),
49196 => conv_std_logic_vector(33, 8),
49197 => conv_std_logic_vector(33, 8),
49198 => conv_std_logic_vector(34, 8),
49199 => conv_std_logic_vector(35, 8),
49200 => conv_std_logic_vector(36, 8),
49201 => conv_std_logic_vector(36, 8),
49202 => conv_std_logic_vector(37, 8),
49203 => conv_std_logic_vector(38, 8),
49204 => conv_std_logic_vector(39, 8),
49205 => conv_std_logic_vector(39, 8),
49206 => conv_std_logic_vector(40, 8),
49207 => conv_std_logic_vector(41, 8),
49208 => conv_std_logic_vector(42, 8),
49209 => conv_std_logic_vector(42, 8),
49210 => conv_std_logic_vector(43, 8),
49211 => conv_std_logic_vector(44, 8),
49212 => conv_std_logic_vector(45, 8),
49213 => conv_std_logic_vector(45, 8),
49214 => conv_std_logic_vector(46, 8),
49215 => conv_std_logic_vector(47, 8),
49216 => conv_std_logic_vector(48, 8),
49217 => conv_std_logic_vector(48, 8),
49218 => conv_std_logic_vector(49, 8),
49219 => conv_std_logic_vector(50, 8),
49220 => conv_std_logic_vector(51, 8),
49221 => conv_std_logic_vector(51, 8),
49222 => conv_std_logic_vector(52, 8),
49223 => conv_std_logic_vector(53, 8),
49224 => conv_std_logic_vector(54, 8),
49225 => conv_std_logic_vector(54, 8),
49226 => conv_std_logic_vector(55, 8),
49227 => conv_std_logic_vector(56, 8),
49228 => conv_std_logic_vector(57, 8),
49229 => conv_std_logic_vector(57, 8),
49230 => conv_std_logic_vector(58, 8),
49231 => conv_std_logic_vector(59, 8),
49232 => conv_std_logic_vector(60, 8),
49233 => conv_std_logic_vector(60, 8),
49234 => conv_std_logic_vector(61, 8),
49235 => conv_std_logic_vector(62, 8),
49236 => conv_std_logic_vector(63, 8),
49237 => conv_std_logic_vector(63, 8),
49238 => conv_std_logic_vector(64, 8),
49239 => conv_std_logic_vector(65, 8),
49240 => conv_std_logic_vector(66, 8),
49241 => conv_std_logic_vector(66, 8),
49242 => conv_std_logic_vector(67, 8),
49243 => conv_std_logic_vector(68, 8),
49244 => conv_std_logic_vector(69, 8),
49245 => conv_std_logic_vector(69, 8),
49246 => conv_std_logic_vector(70, 8),
49247 => conv_std_logic_vector(71, 8),
49248 => conv_std_logic_vector(72, 8),
49249 => conv_std_logic_vector(72, 8),
49250 => conv_std_logic_vector(73, 8),
49251 => conv_std_logic_vector(74, 8),
49252 => conv_std_logic_vector(75, 8),
49253 => conv_std_logic_vector(75, 8),
49254 => conv_std_logic_vector(76, 8),
49255 => conv_std_logic_vector(77, 8),
49256 => conv_std_logic_vector(78, 8),
49257 => conv_std_logic_vector(78, 8),
49258 => conv_std_logic_vector(79, 8),
49259 => conv_std_logic_vector(80, 8),
49260 => conv_std_logic_vector(81, 8),
49261 => conv_std_logic_vector(81, 8),
49262 => conv_std_logic_vector(82, 8),
49263 => conv_std_logic_vector(83, 8),
49264 => conv_std_logic_vector(84, 8),
49265 => conv_std_logic_vector(84, 8),
49266 => conv_std_logic_vector(85, 8),
49267 => conv_std_logic_vector(86, 8),
49268 => conv_std_logic_vector(87, 8),
49269 => conv_std_logic_vector(87, 8),
49270 => conv_std_logic_vector(88, 8),
49271 => conv_std_logic_vector(89, 8),
49272 => conv_std_logic_vector(90, 8),
49273 => conv_std_logic_vector(90, 8),
49274 => conv_std_logic_vector(91, 8),
49275 => conv_std_logic_vector(92, 8),
49276 => conv_std_logic_vector(93, 8),
49277 => conv_std_logic_vector(93, 8),
49278 => conv_std_logic_vector(94, 8),
49279 => conv_std_logic_vector(95, 8),
49280 => conv_std_logic_vector(96, 8),
49281 => conv_std_logic_vector(96, 8),
49282 => conv_std_logic_vector(97, 8),
49283 => conv_std_logic_vector(98, 8),
49284 => conv_std_logic_vector(99, 8),
49285 => conv_std_logic_vector(99, 8),
49286 => conv_std_logic_vector(100, 8),
49287 => conv_std_logic_vector(101, 8),
49288 => conv_std_logic_vector(102, 8),
49289 => conv_std_logic_vector(102, 8),
49290 => conv_std_logic_vector(103, 8),
49291 => conv_std_logic_vector(104, 8),
49292 => conv_std_logic_vector(105, 8),
49293 => conv_std_logic_vector(105, 8),
49294 => conv_std_logic_vector(106, 8),
49295 => conv_std_logic_vector(107, 8),
49296 => conv_std_logic_vector(108, 8),
49297 => conv_std_logic_vector(108, 8),
49298 => conv_std_logic_vector(109, 8),
49299 => conv_std_logic_vector(110, 8),
49300 => conv_std_logic_vector(111, 8),
49301 => conv_std_logic_vector(111, 8),
49302 => conv_std_logic_vector(112, 8),
49303 => conv_std_logic_vector(113, 8),
49304 => conv_std_logic_vector(114, 8),
49305 => conv_std_logic_vector(114, 8),
49306 => conv_std_logic_vector(115, 8),
49307 => conv_std_logic_vector(116, 8),
49308 => conv_std_logic_vector(117, 8),
49309 => conv_std_logic_vector(117, 8),
49310 => conv_std_logic_vector(118, 8),
49311 => conv_std_logic_vector(119, 8),
49312 => conv_std_logic_vector(120, 8),
49313 => conv_std_logic_vector(120, 8),
49314 => conv_std_logic_vector(121, 8),
49315 => conv_std_logic_vector(122, 8),
49316 => conv_std_logic_vector(123, 8),
49317 => conv_std_logic_vector(123, 8),
49318 => conv_std_logic_vector(124, 8),
49319 => conv_std_logic_vector(125, 8),
49320 => conv_std_logic_vector(126, 8),
49321 => conv_std_logic_vector(126, 8),
49322 => conv_std_logic_vector(127, 8),
49323 => conv_std_logic_vector(128, 8),
49324 => conv_std_logic_vector(129, 8),
49325 => conv_std_logic_vector(129, 8),
49326 => conv_std_logic_vector(130, 8),
49327 => conv_std_logic_vector(131, 8),
49328 => conv_std_logic_vector(132, 8),
49329 => conv_std_logic_vector(132, 8),
49330 => conv_std_logic_vector(133, 8),
49331 => conv_std_logic_vector(134, 8),
49332 => conv_std_logic_vector(135, 8),
49333 => conv_std_logic_vector(135, 8),
49334 => conv_std_logic_vector(136, 8),
49335 => conv_std_logic_vector(137, 8),
49336 => conv_std_logic_vector(138, 8),
49337 => conv_std_logic_vector(138, 8),
49338 => conv_std_logic_vector(139, 8),
49339 => conv_std_logic_vector(140, 8),
49340 => conv_std_logic_vector(141, 8),
49341 => conv_std_logic_vector(141, 8),
49342 => conv_std_logic_vector(142, 8),
49343 => conv_std_logic_vector(143, 8),
49344 => conv_std_logic_vector(144, 8),
49345 => conv_std_logic_vector(144, 8),
49346 => conv_std_logic_vector(145, 8),
49347 => conv_std_logic_vector(146, 8),
49348 => conv_std_logic_vector(147, 8),
49349 => conv_std_logic_vector(147, 8),
49350 => conv_std_logic_vector(148, 8),
49351 => conv_std_logic_vector(149, 8),
49352 => conv_std_logic_vector(150, 8),
49353 => conv_std_logic_vector(150, 8),
49354 => conv_std_logic_vector(151, 8),
49355 => conv_std_logic_vector(152, 8),
49356 => conv_std_logic_vector(153, 8),
49357 => conv_std_logic_vector(153, 8),
49358 => conv_std_logic_vector(154, 8),
49359 => conv_std_logic_vector(155, 8),
49360 => conv_std_logic_vector(156, 8),
49361 => conv_std_logic_vector(156, 8),
49362 => conv_std_logic_vector(157, 8),
49363 => conv_std_logic_vector(158, 8),
49364 => conv_std_logic_vector(159, 8),
49365 => conv_std_logic_vector(159, 8),
49366 => conv_std_logic_vector(160, 8),
49367 => conv_std_logic_vector(161, 8),
49368 => conv_std_logic_vector(162, 8),
49369 => conv_std_logic_vector(162, 8),
49370 => conv_std_logic_vector(163, 8),
49371 => conv_std_logic_vector(164, 8),
49372 => conv_std_logic_vector(165, 8),
49373 => conv_std_logic_vector(165, 8),
49374 => conv_std_logic_vector(166, 8),
49375 => conv_std_logic_vector(167, 8),
49376 => conv_std_logic_vector(168, 8),
49377 => conv_std_logic_vector(168, 8),
49378 => conv_std_logic_vector(169, 8),
49379 => conv_std_logic_vector(170, 8),
49380 => conv_std_logic_vector(171, 8),
49381 => conv_std_logic_vector(171, 8),
49382 => conv_std_logic_vector(172, 8),
49383 => conv_std_logic_vector(173, 8),
49384 => conv_std_logic_vector(174, 8),
49385 => conv_std_logic_vector(174, 8),
49386 => conv_std_logic_vector(175, 8),
49387 => conv_std_logic_vector(176, 8),
49388 => conv_std_logic_vector(177, 8),
49389 => conv_std_logic_vector(177, 8),
49390 => conv_std_logic_vector(178, 8),
49391 => conv_std_logic_vector(179, 8),
49392 => conv_std_logic_vector(180, 8),
49393 => conv_std_logic_vector(180, 8),
49394 => conv_std_logic_vector(181, 8),
49395 => conv_std_logic_vector(182, 8),
49396 => conv_std_logic_vector(183, 8),
49397 => conv_std_logic_vector(183, 8),
49398 => conv_std_logic_vector(184, 8),
49399 => conv_std_logic_vector(185, 8),
49400 => conv_std_logic_vector(186, 8),
49401 => conv_std_logic_vector(186, 8),
49402 => conv_std_logic_vector(187, 8),
49403 => conv_std_logic_vector(188, 8),
49404 => conv_std_logic_vector(189, 8),
49405 => conv_std_logic_vector(189, 8),
49406 => conv_std_logic_vector(190, 8),
49407 => conv_std_logic_vector(191, 8),
49408 => conv_std_logic_vector(0, 8),
49409 => conv_std_logic_vector(0, 8),
49410 => conv_std_logic_vector(1, 8),
49411 => conv_std_logic_vector(2, 8),
49412 => conv_std_logic_vector(3, 8),
49413 => conv_std_logic_vector(3, 8),
49414 => conv_std_logic_vector(4, 8),
49415 => conv_std_logic_vector(5, 8),
49416 => conv_std_logic_vector(6, 8),
49417 => conv_std_logic_vector(6, 8),
49418 => conv_std_logic_vector(7, 8),
49419 => conv_std_logic_vector(8, 8),
49420 => conv_std_logic_vector(9, 8),
49421 => conv_std_logic_vector(9, 8),
49422 => conv_std_logic_vector(10, 8),
49423 => conv_std_logic_vector(11, 8),
49424 => conv_std_logic_vector(12, 8),
49425 => conv_std_logic_vector(12, 8),
49426 => conv_std_logic_vector(13, 8),
49427 => conv_std_logic_vector(14, 8),
49428 => conv_std_logic_vector(15, 8),
49429 => conv_std_logic_vector(15, 8),
49430 => conv_std_logic_vector(16, 8),
49431 => conv_std_logic_vector(17, 8),
49432 => conv_std_logic_vector(18, 8),
49433 => conv_std_logic_vector(18, 8),
49434 => conv_std_logic_vector(19, 8),
49435 => conv_std_logic_vector(20, 8),
49436 => conv_std_logic_vector(21, 8),
49437 => conv_std_logic_vector(21, 8),
49438 => conv_std_logic_vector(22, 8),
49439 => conv_std_logic_vector(23, 8),
49440 => conv_std_logic_vector(24, 8),
49441 => conv_std_logic_vector(24, 8),
49442 => conv_std_logic_vector(25, 8),
49443 => conv_std_logic_vector(26, 8),
49444 => conv_std_logic_vector(27, 8),
49445 => conv_std_logic_vector(27, 8),
49446 => conv_std_logic_vector(28, 8),
49447 => conv_std_logic_vector(29, 8),
49448 => conv_std_logic_vector(30, 8),
49449 => conv_std_logic_vector(30, 8),
49450 => conv_std_logic_vector(31, 8),
49451 => conv_std_logic_vector(32, 8),
49452 => conv_std_logic_vector(33, 8),
49453 => conv_std_logic_vector(33, 8),
49454 => conv_std_logic_vector(34, 8),
49455 => conv_std_logic_vector(35, 8),
49456 => conv_std_logic_vector(36, 8),
49457 => conv_std_logic_vector(36, 8),
49458 => conv_std_logic_vector(37, 8),
49459 => conv_std_logic_vector(38, 8),
49460 => conv_std_logic_vector(39, 8),
49461 => conv_std_logic_vector(39, 8),
49462 => conv_std_logic_vector(40, 8),
49463 => conv_std_logic_vector(41, 8),
49464 => conv_std_logic_vector(42, 8),
49465 => conv_std_logic_vector(42, 8),
49466 => conv_std_logic_vector(43, 8),
49467 => conv_std_logic_vector(44, 8),
49468 => conv_std_logic_vector(45, 8),
49469 => conv_std_logic_vector(45, 8),
49470 => conv_std_logic_vector(46, 8),
49471 => conv_std_logic_vector(47, 8),
49472 => conv_std_logic_vector(48, 8),
49473 => conv_std_logic_vector(49, 8),
49474 => conv_std_logic_vector(49, 8),
49475 => conv_std_logic_vector(50, 8),
49476 => conv_std_logic_vector(51, 8),
49477 => conv_std_logic_vector(52, 8),
49478 => conv_std_logic_vector(52, 8),
49479 => conv_std_logic_vector(53, 8),
49480 => conv_std_logic_vector(54, 8),
49481 => conv_std_logic_vector(55, 8),
49482 => conv_std_logic_vector(55, 8),
49483 => conv_std_logic_vector(56, 8),
49484 => conv_std_logic_vector(57, 8),
49485 => conv_std_logic_vector(58, 8),
49486 => conv_std_logic_vector(58, 8),
49487 => conv_std_logic_vector(59, 8),
49488 => conv_std_logic_vector(60, 8),
49489 => conv_std_logic_vector(61, 8),
49490 => conv_std_logic_vector(61, 8),
49491 => conv_std_logic_vector(62, 8),
49492 => conv_std_logic_vector(63, 8),
49493 => conv_std_logic_vector(64, 8),
49494 => conv_std_logic_vector(64, 8),
49495 => conv_std_logic_vector(65, 8),
49496 => conv_std_logic_vector(66, 8),
49497 => conv_std_logic_vector(67, 8),
49498 => conv_std_logic_vector(67, 8),
49499 => conv_std_logic_vector(68, 8),
49500 => conv_std_logic_vector(69, 8),
49501 => conv_std_logic_vector(70, 8),
49502 => conv_std_logic_vector(70, 8),
49503 => conv_std_logic_vector(71, 8),
49504 => conv_std_logic_vector(72, 8),
49505 => conv_std_logic_vector(73, 8),
49506 => conv_std_logic_vector(73, 8),
49507 => conv_std_logic_vector(74, 8),
49508 => conv_std_logic_vector(75, 8),
49509 => conv_std_logic_vector(76, 8),
49510 => conv_std_logic_vector(76, 8),
49511 => conv_std_logic_vector(77, 8),
49512 => conv_std_logic_vector(78, 8),
49513 => conv_std_logic_vector(79, 8),
49514 => conv_std_logic_vector(79, 8),
49515 => conv_std_logic_vector(80, 8),
49516 => conv_std_logic_vector(81, 8),
49517 => conv_std_logic_vector(82, 8),
49518 => conv_std_logic_vector(82, 8),
49519 => conv_std_logic_vector(83, 8),
49520 => conv_std_logic_vector(84, 8),
49521 => conv_std_logic_vector(85, 8),
49522 => conv_std_logic_vector(85, 8),
49523 => conv_std_logic_vector(86, 8),
49524 => conv_std_logic_vector(87, 8),
49525 => conv_std_logic_vector(88, 8),
49526 => conv_std_logic_vector(88, 8),
49527 => conv_std_logic_vector(89, 8),
49528 => conv_std_logic_vector(90, 8),
49529 => conv_std_logic_vector(91, 8),
49530 => conv_std_logic_vector(91, 8),
49531 => conv_std_logic_vector(92, 8),
49532 => conv_std_logic_vector(93, 8),
49533 => conv_std_logic_vector(94, 8),
49534 => conv_std_logic_vector(94, 8),
49535 => conv_std_logic_vector(95, 8),
49536 => conv_std_logic_vector(96, 8),
49537 => conv_std_logic_vector(97, 8),
49538 => conv_std_logic_vector(98, 8),
49539 => conv_std_logic_vector(98, 8),
49540 => conv_std_logic_vector(99, 8),
49541 => conv_std_logic_vector(100, 8),
49542 => conv_std_logic_vector(101, 8),
49543 => conv_std_logic_vector(101, 8),
49544 => conv_std_logic_vector(102, 8),
49545 => conv_std_logic_vector(103, 8),
49546 => conv_std_logic_vector(104, 8),
49547 => conv_std_logic_vector(104, 8),
49548 => conv_std_logic_vector(105, 8),
49549 => conv_std_logic_vector(106, 8),
49550 => conv_std_logic_vector(107, 8),
49551 => conv_std_logic_vector(107, 8),
49552 => conv_std_logic_vector(108, 8),
49553 => conv_std_logic_vector(109, 8),
49554 => conv_std_logic_vector(110, 8),
49555 => conv_std_logic_vector(110, 8),
49556 => conv_std_logic_vector(111, 8),
49557 => conv_std_logic_vector(112, 8),
49558 => conv_std_logic_vector(113, 8),
49559 => conv_std_logic_vector(113, 8),
49560 => conv_std_logic_vector(114, 8),
49561 => conv_std_logic_vector(115, 8),
49562 => conv_std_logic_vector(116, 8),
49563 => conv_std_logic_vector(116, 8),
49564 => conv_std_logic_vector(117, 8),
49565 => conv_std_logic_vector(118, 8),
49566 => conv_std_logic_vector(119, 8),
49567 => conv_std_logic_vector(119, 8),
49568 => conv_std_logic_vector(120, 8),
49569 => conv_std_logic_vector(121, 8),
49570 => conv_std_logic_vector(122, 8),
49571 => conv_std_logic_vector(122, 8),
49572 => conv_std_logic_vector(123, 8),
49573 => conv_std_logic_vector(124, 8),
49574 => conv_std_logic_vector(125, 8),
49575 => conv_std_logic_vector(125, 8),
49576 => conv_std_logic_vector(126, 8),
49577 => conv_std_logic_vector(127, 8),
49578 => conv_std_logic_vector(128, 8),
49579 => conv_std_logic_vector(128, 8),
49580 => conv_std_logic_vector(129, 8),
49581 => conv_std_logic_vector(130, 8),
49582 => conv_std_logic_vector(131, 8),
49583 => conv_std_logic_vector(131, 8),
49584 => conv_std_logic_vector(132, 8),
49585 => conv_std_logic_vector(133, 8),
49586 => conv_std_logic_vector(134, 8),
49587 => conv_std_logic_vector(134, 8),
49588 => conv_std_logic_vector(135, 8),
49589 => conv_std_logic_vector(136, 8),
49590 => conv_std_logic_vector(137, 8),
49591 => conv_std_logic_vector(137, 8),
49592 => conv_std_logic_vector(138, 8),
49593 => conv_std_logic_vector(139, 8),
49594 => conv_std_logic_vector(140, 8),
49595 => conv_std_logic_vector(140, 8),
49596 => conv_std_logic_vector(141, 8),
49597 => conv_std_logic_vector(142, 8),
49598 => conv_std_logic_vector(143, 8),
49599 => conv_std_logic_vector(143, 8),
49600 => conv_std_logic_vector(144, 8),
49601 => conv_std_logic_vector(145, 8),
49602 => conv_std_logic_vector(146, 8),
49603 => conv_std_logic_vector(147, 8),
49604 => conv_std_logic_vector(147, 8),
49605 => conv_std_logic_vector(148, 8),
49606 => conv_std_logic_vector(149, 8),
49607 => conv_std_logic_vector(150, 8),
49608 => conv_std_logic_vector(150, 8),
49609 => conv_std_logic_vector(151, 8),
49610 => conv_std_logic_vector(152, 8),
49611 => conv_std_logic_vector(153, 8),
49612 => conv_std_logic_vector(153, 8),
49613 => conv_std_logic_vector(154, 8),
49614 => conv_std_logic_vector(155, 8),
49615 => conv_std_logic_vector(156, 8),
49616 => conv_std_logic_vector(156, 8),
49617 => conv_std_logic_vector(157, 8),
49618 => conv_std_logic_vector(158, 8),
49619 => conv_std_logic_vector(159, 8),
49620 => conv_std_logic_vector(159, 8),
49621 => conv_std_logic_vector(160, 8),
49622 => conv_std_logic_vector(161, 8),
49623 => conv_std_logic_vector(162, 8),
49624 => conv_std_logic_vector(162, 8),
49625 => conv_std_logic_vector(163, 8),
49626 => conv_std_logic_vector(164, 8),
49627 => conv_std_logic_vector(165, 8),
49628 => conv_std_logic_vector(165, 8),
49629 => conv_std_logic_vector(166, 8),
49630 => conv_std_logic_vector(167, 8),
49631 => conv_std_logic_vector(168, 8),
49632 => conv_std_logic_vector(168, 8),
49633 => conv_std_logic_vector(169, 8),
49634 => conv_std_logic_vector(170, 8),
49635 => conv_std_logic_vector(171, 8),
49636 => conv_std_logic_vector(171, 8),
49637 => conv_std_logic_vector(172, 8),
49638 => conv_std_logic_vector(173, 8),
49639 => conv_std_logic_vector(174, 8),
49640 => conv_std_logic_vector(174, 8),
49641 => conv_std_logic_vector(175, 8),
49642 => conv_std_logic_vector(176, 8),
49643 => conv_std_logic_vector(177, 8),
49644 => conv_std_logic_vector(177, 8),
49645 => conv_std_logic_vector(178, 8),
49646 => conv_std_logic_vector(179, 8),
49647 => conv_std_logic_vector(180, 8),
49648 => conv_std_logic_vector(180, 8),
49649 => conv_std_logic_vector(181, 8),
49650 => conv_std_logic_vector(182, 8),
49651 => conv_std_logic_vector(183, 8),
49652 => conv_std_logic_vector(183, 8),
49653 => conv_std_logic_vector(184, 8),
49654 => conv_std_logic_vector(185, 8),
49655 => conv_std_logic_vector(186, 8),
49656 => conv_std_logic_vector(186, 8),
49657 => conv_std_logic_vector(187, 8),
49658 => conv_std_logic_vector(188, 8),
49659 => conv_std_logic_vector(189, 8),
49660 => conv_std_logic_vector(189, 8),
49661 => conv_std_logic_vector(190, 8),
49662 => conv_std_logic_vector(191, 8),
49663 => conv_std_logic_vector(192, 8),
49664 => conv_std_logic_vector(0, 8),
49665 => conv_std_logic_vector(0, 8),
49666 => conv_std_logic_vector(1, 8),
49667 => conv_std_logic_vector(2, 8),
49668 => conv_std_logic_vector(3, 8),
49669 => conv_std_logic_vector(3, 8),
49670 => conv_std_logic_vector(4, 8),
49671 => conv_std_logic_vector(5, 8),
49672 => conv_std_logic_vector(6, 8),
49673 => conv_std_logic_vector(6, 8),
49674 => conv_std_logic_vector(7, 8),
49675 => conv_std_logic_vector(8, 8),
49676 => conv_std_logic_vector(9, 8),
49677 => conv_std_logic_vector(9, 8),
49678 => conv_std_logic_vector(10, 8),
49679 => conv_std_logic_vector(11, 8),
49680 => conv_std_logic_vector(12, 8),
49681 => conv_std_logic_vector(12, 8),
49682 => conv_std_logic_vector(13, 8),
49683 => conv_std_logic_vector(14, 8),
49684 => conv_std_logic_vector(15, 8),
49685 => conv_std_logic_vector(15, 8),
49686 => conv_std_logic_vector(16, 8),
49687 => conv_std_logic_vector(17, 8),
49688 => conv_std_logic_vector(18, 8),
49689 => conv_std_logic_vector(18, 8),
49690 => conv_std_logic_vector(19, 8),
49691 => conv_std_logic_vector(20, 8),
49692 => conv_std_logic_vector(21, 8),
49693 => conv_std_logic_vector(21, 8),
49694 => conv_std_logic_vector(22, 8),
49695 => conv_std_logic_vector(23, 8),
49696 => conv_std_logic_vector(24, 8),
49697 => conv_std_logic_vector(25, 8),
49698 => conv_std_logic_vector(25, 8),
49699 => conv_std_logic_vector(26, 8),
49700 => conv_std_logic_vector(27, 8),
49701 => conv_std_logic_vector(28, 8),
49702 => conv_std_logic_vector(28, 8),
49703 => conv_std_logic_vector(29, 8),
49704 => conv_std_logic_vector(30, 8),
49705 => conv_std_logic_vector(31, 8),
49706 => conv_std_logic_vector(31, 8),
49707 => conv_std_logic_vector(32, 8),
49708 => conv_std_logic_vector(33, 8),
49709 => conv_std_logic_vector(34, 8),
49710 => conv_std_logic_vector(34, 8),
49711 => conv_std_logic_vector(35, 8),
49712 => conv_std_logic_vector(36, 8),
49713 => conv_std_logic_vector(37, 8),
49714 => conv_std_logic_vector(37, 8),
49715 => conv_std_logic_vector(38, 8),
49716 => conv_std_logic_vector(39, 8),
49717 => conv_std_logic_vector(40, 8),
49718 => conv_std_logic_vector(40, 8),
49719 => conv_std_logic_vector(41, 8),
49720 => conv_std_logic_vector(42, 8),
49721 => conv_std_logic_vector(43, 8),
49722 => conv_std_logic_vector(43, 8),
49723 => conv_std_logic_vector(44, 8),
49724 => conv_std_logic_vector(45, 8),
49725 => conv_std_logic_vector(46, 8),
49726 => conv_std_logic_vector(46, 8),
49727 => conv_std_logic_vector(47, 8),
49728 => conv_std_logic_vector(48, 8),
49729 => conv_std_logic_vector(49, 8),
49730 => conv_std_logic_vector(50, 8),
49731 => conv_std_logic_vector(50, 8),
49732 => conv_std_logic_vector(51, 8),
49733 => conv_std_logic_vector(52, 8),
49734 => conv_std_logic_vector(53, 8),
49735 => conv_std_logic_vector(53, 8),
49736 => conv_std_logic_vector(54, 8),
49737 => conv_std_logic_vector(55, 8),
49738 => conv_std_logic_vector(56, 8),
49739 => conv_std_logic_vector(56, 8),
49740 => conv_std_logic_vector(57, 8),
49741 => conv_std_logic_vector(58, 8),
49742 => conv_std_logic_vector(59, 8),
49743 => conv_std_logic_vector(59, 8),
49744 => conv_std_logic_vector(60, 8),
49745 => conv_std_logic_vector(61, 8),
49746 => conv_std_logic_vector(62, 8),
49747 => conv_std_logic_vector(62, 8),
49748 => conv_std_logic_vector(63, 8),
49749 => conv_std_logic_vector(64, 8),
49750 => conv_std_logic_vector(65, 8),
49751 => conv_std_logic_vector(65, 8),
49752 => conv_std_logic_vector(66, 8),
49753 => conv_std_logic_vector(67, 8),
49754 => conv_std_logic_vector(68, 8),
49755 => conv_std_logic_vector(68, 8),
49756 => conv_std_logic_vector(69, 8),
49757 => conv_std_logic_vector(70, 8),
49758 => conv_std_logic_vector(71, 8),
49759 => conv_std_logic_vector(71, 8),
49760 => conv_std_logic_vector(72, 8),
49761 => conv_std_logic_vector(73, 8),
49762 => conv_std_logic_vector(74, 8),
49763 => conv_std_logic_vector(75, 8),
49764 => conv_std_logic_vector(75, 8),
49765 => conv_std_logic_vector(76, 8),
49766 => conv_std_logic_vector(77, 8),
49767 => conv_std_logic_vector(78, 8),
49768 => conv_std_logic_vector(78, 8),
49769 => conv_std_logic_vector(79, 8),
49770 => conv_std_logic_vector(80, 8),
49771 => conv_std_logic_vector(81, 8),
49772 => conv_std_logic_vector(81, 8),
49773 => conv_std_logic_vector(82, 8),
49774 => conv_std_logic_vector(83, 8),
49775 => conv_std_logic_vector(84, 8),
49776 => conv_std_logic_vector(84, 8),
49777 => conv_std_logic_vector(85, 8),
49778 => conv_std_logic_vector(86, 8),
49779 => conv_std_logic_vector(87, 8),
49780 => conv_std_logic_vector(87, 8),
49781 => conv_std_logic_vector(88, 8),
49782 => conv_std_logic_vector(89, 8),
49783 => conv_std_logic_vector(90, 8),
49784 => conv_std_logic_vector(90, 8),
49785 => conv_std_logic_vector(91, 8),
49786 => conv_std_logic_vector(92, 8),
49787 => conv_std_logic_vector(93, 8),
49788 => conv_std_logic_vector(93, 8),
49789 => conv_std_logic_vector(94, 8),
49790 => conv_std_logic_vector(95, 8),
49791 => conv_std_logic_vector(96, 8),
49792 => conv_std_logic_vector(97, 8),
49793 => conv_std_logic_vector(97, 8),
49794 => conv_std_logic_vector(98, 8),
49795 => conv_std_logic_vector(99, 8),
49796 => conv_std_logic_vector(100, 8),
49797 => conv_std_logic_vector(100, 8),
49798 => conv_std_logic_vector(101, 8),
49799 => conv_std_logic_vector(102, 8),
49800 => conv_std_logic_vector(103, 8),
49801 => conv_std_logic_vector(103, 8),
49802 => conv_std_logic_vector(104, 8),
49803 => conv_std_logic_vector(105, 8),
49804 => conv_std_logic_vector(106, 8),
49805 => conv_std_logic_vector(106, 8),
49806 => conv_std_logic_vector(107, 8),
49807 => conv_std_logic_vector(108, 8),
49808 => conv_std_logic_vector(109, 8),
49809 => conv_std_logic_vector(109, 8),
49810 => conv_std_logic_vector(110, 8),
49811 => conv_std_logic_vector(111, 8),
49812 => conv_std_logic_vector(112, 8),
49813 => conv_std_logic_vector(112, 8),
49814 => conv_std_logic_vector(113, 8),
49815 => conv_std_logic_vector(114, 8),
49816 => conv_std_logic_vector(115, 8),
49817 => conv_std_logic_vector(115, 8),
49818 => conv_std_logic_vector(116, 8),
49819 => conv_std_logic_vector(117, 8),
49820 => conv_std_logic_vector(118, 8),
49821 => conv_std_logic_vector(118, 8),
49822 => conv_std_logic_vector(119, 8),
49823 => conv_std_logic_vector(120, 8),
49824 => conv_std_logic_vector(121, 8),
49825 => conv_std_logic_vector(122, 8),
49826 => conv_std_logic_vector(122, 8),
49827 => conv_std_logic_vector(123, 8),
49828 => conv_std_logic_vector(124, 8),
49829 => conv_std_logic_vector(125, 8),
49830 => conv_std_logic_vector(125, 8),
49831 => conv_std_logic_vector(126, 8),
49832 => conv_std_logic_vector(127, 8),
49833 => conv_std_logic_vector(128, 8),
49834 => conv_std_logic_vector(128, 8),
49835 => conv_std_logic_vector(129, 8),
49836 => conv_std_logic_vector(130, 8),
49837 => conv_std_logic_vector(131, 8),
49838 => conv_std_logic_vector(131, 8),
49839 => conv_std_logic_vector(132, 8),
49840 => conv_std_logic_vector(133, 8),
49841 => conv_std_logic_vector(134, 8),
49842 => conv_std_logic_vector(134, 8),
49843 => conv_std_logic_vector(135, 8),
49844 => conv_std_logic_vector(136, 8),
49845 => conv_std_logic_vector(137, 8),
49846 => conv_std_logic_vector(137, 8),
49847 => conv_std_logic_vector(138, 8),
49848 => conv_std_logic_vector(139, 8),
49849 => conv_std_logic_vector(140, 8),
49850 => conv_std_logic_vector(140, 8),
49851 => conv_std_logic_vector(141, 8),
49852 => conv_std_logic_vector(142, 8),
49853 => conv_std_logic_vector(143, 8),
49854 => conv_std_logic_vector(143, 8),
49855 => conv_std_logic_vector(144, 8),
49856 => conv_std_logic_vector(145, 8),
49857 => conv_std_logic_vector(146, 8),
49858 => conv_std_logic_vector(147, 8),
49859 => conv_std_logic_vector(147, 8),
49860 => conv_std_logic_vector(148, 8),
49861 => conv_std_logic_vector(149, 8),
49862 => conv_std_logic_vector(150, 8),
49863 => conv_std_logic_vector(150, 8),
49864 => conv_std_logic_vector(151, 8),
49865 => conv_std_logic_vector(152, 8),
49866 => conv_std_logic_vector(153, 8),
49867 => conv_std_logic_vector(153, 8),
49868 => conv_std_logic_vector(154, 8),
49869 => conv_std_logic_vector(155, 8),
49870 => conv_std_logic_vector(156, 8),
49871 => conv_std_logic_vector(156, 8),
49872 => conv_std_logic_vector(157, 8),
49873 => conv_std_logic_vector(158, 8),
49874 => conv_std_logic_vector(159, 8),
49875 => conv_std_logic_vector(159, 8),
49876 => conv_std_logic_vector(160, 8),
49877 => conv_std_logic_vector(161, 8),
49878 => conv_std_logic_vector(162, 8),
49879 => conv_std_logic_vector(162, 8),
49880 => conv_std_logic_vector(163, 8),
49881 => conv_std_logic_vector(164, 8),
49882 => conv_std_logic_vector(165, 8),
49883 => conv_std_logic_vector(165, 8),
49884 => conv_std_logic_vector(166, 8),
49885 => conv_std_logic_vector(167, 8),
49886 => conv_std_logic_vector(168, 8),
49887 => conv_std_logic_vector(168, 8),
49888 => conv_std_logic_vector(169, 8),
49889 => conv_std_logic_vector(170, 8),
49890 => conv_std_logic_vector(171, 8),
49891 => conv_std_logic_vector(172, 8),
49892 => conv_std_logic_vector(172, 8),
49893 => conv_std_logic_vector(173, 8),
49894 => conv_std_logic_vector(174, 8),
49895 => conv_std_logic_vector(175, 8),
49896 => conv_std_logic_vector(175, 8),
49897 => conv_std_logic_vector(176, 8),
49898 => conv_std_logic_vector(177, 8),
49899 => conv_std_logic_vector(178, 8),
49900 => conv_std_logic_vector(178, 8),
49901 => conv_std_logic_vector(179, 8),
49902 => conv_std_logic_vector(180, 8),
49903 => conv_std_logic_vector(181, 8),
49904 => conv_std_logic_vector(181, 8),
49905 => conv_std_logic_vector(182, 8),
49906 => conv_std_logic_vector(183, 8),
49907 => conv_std_logic_vector(184, 8),
49908 => conv_std_logic_vector(184, 8),
49909 => conv_std_logic_vector(185, 8),
49910 => conv_std_logic_vector(186, 8),
49911 => conv_std_logic_vector(187, 8),
49912 => conv_std_logic_vector(187, 8),
49913 => conv_std_logic_vector(188, 8),
49914 => conv_std_logic_vector(189, 8),
49915 => conv_std_logic_vector(190, 8),
49916 => conv_std_logic_vector(190, 8),
49917 => conv_std_logic_vector(191, 8),
49918 => conv_std_logic_vector(192, 8),
49919 => conv_std_logic_vector(193, 8),
49920 => conv_std_logic_vector(0, 8),
49921 => conv_std_logic_vector(0, 8),
49922 => conv_std_logic_vector(1, 8),
49923 => conv_std_logic_vector(2, 8),
49924 => conv_std_logic_vector(3, 8),
49925 => conv_std_logic_vector(3, 8),
49926 => conv_std_logic_vector(4, 8),
49927 => conv_std_logic_vector(5, 8),
49928 => conv_std_logic_vector(6, 8),
49929 => conv_std_logic_vector(6, 8),
49930 => conv_std_logic_vector(7, 8),
49931 => conv_std_logic_vector(8, 8),
49932 => conv_std_logic_vector(9, 8),
49933 => conv_std_logic_vector(9, 8),
49934 => conv_std_logic_vector(10, 8),
49935 => conv_std_logic_vector(11, 8),
49936 => conv_std_logic_vector(12, 8),
49937 => conv_std_logic_vector(12, 8),
49938 => conv_std_logic_vector(13, 8),
49939 => conv_std_logic_vector(14, 8),
49940 => conv_std_logic_vector(15, 8),
49941 => conv_std_logic_vector(15, 8),
49942 => conv_std_logic_vector(16, 8),
49943 => conv_std_logic_vector(17, 8),
49944 => conv_std_logic_vector(18, 8),
49945 => conv_std_logic_vector(19, 8),
49946 => conv_std_logic_vector(19, 8),
49947 => conv_std_logic_vector(20, 8),
49948 => conv_std_logic_vector(21, 8),
49949 => conv_std_logic_vector(22, 8),
49950 => conv_std_logic_vector(22, 8),
49951 => conv_std_logic_vector(23, 8),
49952 => conv_std_logic_vector(24, 8),
49953 => conv_std_logic_vector(25, 8),
49954 => conv_std_logic_vector(25, 8),
49955 => conv_std_logic_vector(26, 8),
49956 => conv_std_logic_vector(27, 8),
49957 => conv_std_logic_vector(28, 8),
49958 => conv_std_logic_vector(28, 8),
49959 => conv_std_logic_vector(29, 8),
49960 => conv_std_logic_vector(30, 8),
49961 => conv_std_logic_vector(31, 8),
49962 => conv_std_logic_vector(31, 8),
49963 => conv_std_logic_vector(32, 8),
49964 => conv_std_logic_vector(33, 8),
49965 => conv_std_logic_vector(34, 8),
49966 => conv_std_logic_vector(35, 8),
49967 => conv_std_logic_vector(35, 8),
49968 => conv_std_logic_vector(36, 8),
49969 => conv_std_logic_vector(37, 8),
49970 => conv_std_logic_vector(38, 8),
49971 => conv_std_logic_vector(38, 8),
49972 => conv_std_logic_vector(39, 8),
49973 => conv_std_logic_vector(40, 8),
49974 => conv_std_logic_vector(41, 8),
49975 => conv_std_logic_vector(41, 8),
49976 => conv_std_logic_vector(42, 8),
49977 => conv_std_logic_vector(43, 8),
49978 => conv_std_logic_vector(44, 8),
49979 => conv_std_logic_vector(44, 8),
49980 => conv_std_logic_vector(45, 8),
49981 => conv_std_logic_vector(46, 8),
49982 => conv_std_logic_vector(47, 8),
49983 => conv_std_logic_vector(47, 8),
49984 => conv_std_logic_vector(48, 8),
49985 => conv_std_logic_vector(49, 8),
49986 => conv_std_logic_vector(50, 8),
49987 => conv_std_logic_vector(51, 8),
49988 => conv_std_logic_vector(51, 8),
49989 => conv_std_logic_vector(52, 8),
49990 => conv_std_logic_vector(53, 8),
49991 => conv_std_logic_vector(54, 8),
49992 => conv_std_logic_vector(54, 8),
49993 => conv_std_logic_vector(55, 8),
49994 => conv_std_logic_vector(56, 8),
49995 => conv_std_logic_vector(57, 8),
49996 => conv_std_logic_vector(57, 8),
49997 => conv_std_logic_vector(58, 8),
49998 => conv_std_logic_vector(59, 8),
49999 => conv_std_logic_vector(60, 8),
50000 => conv_std_logic_vector(60, 8),
50001 => conv_std_logic_vector(61, 8),
50002 => conv_std_logic_vector(62, 8),
50003 => conv_std_logic_vector(63, 8),
50004 => conv_std_logic_vector(63, 8),
50005 => conv_std_logic_vector(64, 8),
50006 => conv_std_logic_vector(65, 8),
50007 => conv_std_logic_vector(66, 8),
50008 => conv_std_logic_vector(67, 8),
50009 => conv_std_logic_vector(67, 8),
50010 => conv_std_logic_vector(68, 8),
50011 => conv_std_logic_vector(69, 8),
50012 => conv_std_logic_vector(70, 8),
50013 => conv_std_logic_vector(70, 8),
50014 => conv_std_logic_vector(71, 8),
50015 => conv_std_logic_vector(72, 8),
50016 => conv_std_logic_vector(73, 8),
50017 => conv_std_logic_vector(73, 8),
50018 => conv_std_logic_vector(74, 8),
50019 => conv_std_logic_vector(75, 8),
50020 => conv_std_logic_vector(76, 8),
50021 => conv_std_logic_vector(76, 8),
50022 => conv_std_logic_vector(77, 8),
50023 => conv_std_logic_vector(78, 8),
50024 => conv_std_logic_vector(79, 8),
50025 => conv_std_logic_vector(79, 8),
50026 => conv_std_logic_vector(80, 8),
50027 => conv_std_logic_vector(81, 8),
50028 => conv_std_logic_vector(82, 8),
50029 => conv_std_logic_vector(83, 8),
50030 => conv_std_logic_vector(83, 8),
50031 => conv_std_logic_vector(84, 8),
50032 => conv_std_logic_vector(85, 8),
50033 => conv_std_logic_vector(86, 8),
50034 => conv_std_logic_vector(86, 8),
50035 => conv_std_logic_vector(87, 8),
50036 => conv_std_logic_vector(88, 8),
50037 => conv_std_logic_vector(89, 8),
50038 => conv_std_logic_vector(89, 8),
50039 => conv_std_logic_vector(90, 8),
50040 => conv_std_logic_vector(91, 8),
50041 => conv_std_logic_vector(92, 8),
50042 => conv_std_logic_vector(92, 8),
50043 => conv_std_logic_vector(93, 8),
50044 => conv_std_logic_vector(94, 8),
50045 => conv_std_logic_vector(95, 8),
50046 => conv_std_logic_vector(95, 8),
50047 => conv_std_logic_vector(96, 8),
50048 => conv_std_logic_vector(97, 8),
50049 => conv_std_logic_vector(98, 8),
50050 => conv_std_logic_vector(99, 8),
50051 => conv_std_logic_vector(99, 8),
50052 => conv_std_logic_vector(100, 8),
50053 => conv_std_logic_vector(101, 8),
50054 => conv_std_logic_vector(102, 8),
50055 => conv_std_logic_vector(102, 8),
50056 => conv_std_logic_vector(103, 8),
50057 => conv_std_logic_vector(104, 8),
50058 => conv_std_logic_vector(105, 8),
50059 => conv_std_logic_vector(105, 8),
50060 => conv_std_logic_vector(106, 8),
50061 => conv_std_logic_vector(107, 8),
50062 => conv_std_logic_vector(108, 8),
50063 => conv_std_logic_vector(108, 8),
50064 => conv_std_logic_vector(109, 8),
50065 => conv_std_logic_vector(110, 8),
50066 => conv_std_logic_vector(111, 8),
50067 => conv_std_logic_vector(111, 8),
50068 => conv_std_logic_vector(112, 8),
50069 => conv_std_logic_vector(113, 8),
50070 => conv_std_logic_vector(114, 8),
50071 => conv_std_logic_vector(115, 8),
50072 => conv_std_logic_vector(115, 8),
50073 => conv_std_logic_vector(116, 8),
50074 => conv_std_logic_vector(117, 8),
50075 => conv_std_logic_vector(118, 8),
50076 => conv_std_logic_vector(118, 8),
50077 => conv_std_logic_vector(119, 8),
50078 => conv_std_logic_vector(120, 8),
50079 => conv_std_logic_vector(121, 8),
50080 => conv_std_logic_vector(121, 8),
50081 => conv_std_logic_vector(122, 8),
50082 => conv_std_logic_vector(123, 8),
50083 => conv_std_logic_vector(124, 8),
50084 => conv_std_logic_vector(124, 8),
50085 => conv_std_logic_vector(125, 8),
50086 => conv_std_logic_vector(126, 8),
50087 => conv_std_logic_vector(127, 8),
50088 => conv_std_logic_vector(127, 8),
50089 => conv_std_logic_vector(128, 8),
50090 => conv_std_logic_vector(129, 8),
50091 => conv_std_logic_vector(130, 8),
50092 => conv_std_logic_vector(131, 8),
50093 => conv_std_logic_vector(131, 8),
50094 => conv_std_logic_vector(132, 8),
50095 => conv_std_logic_vector(133, 8),
50096 => conv_std_logic_vector(134, 8),
50097 => conv_std_logic_vector(134, 8),
50098 => conv_std_logic_vector(135, 8),
50099 => conv_std_logic_vector(136, 8),
50100 => conv_std_logic_vector(137, 8),
50101 => conv_std_logic_vector(137, 8),
50102 => conv_std_logic_vector(138, 8),
50103 => conv_std_logic_vector(139, 8),
50104 => conv_std_logic_vector(140, 8),
50105 => conv_std_logic_vector(140, 8),
50106 => conv_std_logic_vector(141, 8),
50107 => conv_std_logic_vector(142, 8),
50108 => conv_std_logic_vector(143, 8),
50109 => conv_std_logic_vector(143, 8),
50110 => conv_std_logic_vector(144, 8),
50111 => conv_std_logic_vector(145, 8),
50112 => conv_std_logic_vector(146, 8),
50113 => conv_std_logic_vector(147, 8),
50114 => conv_std_logic_vector(147, 8),
50115 => conv_std_logic_vector(148, 8),
50116 => conv_std_logic_vector(149, 8),
50117 => conv_std_logic_vector(150, 8),
50118 => conv_std_logic_vector(150, 8),
50119 => conv_std_logic_vector(151, 8),
50120 => conv_std_logic_vector(152, 8),
50121 => conv_std_logic_vector(153, 8),
50122 => conv_std_logic_vector(153, 8),
50123 => conv_std_logic_vector(154, 8),
50124 => conv_std_logic_vector(155, 8),
50125 => conv_std_logic_vector(156, 8),
50126 => conv_std_logic_vector(156, 8),
50127 => conv_std_logic_vector(157, 8),
50128 => conv_std_logic_vector(158, 8),
50129 => conv_std_logic_vector(159, 8),
50130 => conv_std_logic_vector(159, 8),
50131 => conv_std_logic_vector(160, 8),
50132 => conv_std_logic_vector(161, 8),
50133 => conv_std_logic_vector(162, 8),
50134 => conv_std_logic_vector(163, 8),
50135 => conv_std_logic_vector(163, 8),
50136 => conv_std_logic_vector(164, 8),
50137 => conv_std_logic_vector(165, 8),
50138 => conv_std_logic_vector(166, 8),
50139 => conv_std_logic_vector(166, 8),
50140 => conv_std_logic_vector(167, 8),
50141 => conv_std_logic_vector(168, 8),
50142 => conv_std_logic_vector(169, 8),
50143 => conv_std_logic_vector(169, 8),
50144 => conv_std_logic_vector(170, 8),
50145 => conv_std_logic_vector(171, 8),
50146 => conv_std_logic_vector(172, 8),
50147 => conv_std_logic_vector(172, 8),
50148 => conv_std_logic_vector(173, 8),
50149 => conv_std_logic_vector(174, 8),
50150 => conv_std_logic_vector(175, 8),
50151 => conv_std_logic_vector(175, 8),
50152 => conv_std_logic_vector(176, 8),
50153 => conv_std_logic_vector(177, 8),
50154 => conv_std_logic_vector(178, 8),
50155 => conv_std_logic_vector(179, 8),
50156 => conv_std_logic_vector(179, 8),
50157 => conv_std_logic_vector(180, 8),
50158 => conv_std_logic_vector(181, 8),
50159 => conv_std_logic_vector(182, 8),
50160 => conv_std_logic_vector(182, 8),
50161 => conv_std_logic_vector(183, 8),
50162 => conv_std_logic_vector(184, 8),
50163 => conv_std_logic_vector(185, 8),
50164 => conv_std_logic_vector(185, 8),
50165 => conv_std_logic_vector(186, 8),
50166 => conv_std_logic_vector(187, 8),
50167 => conv_std_logic_vector(188, 8),
50168 => conv_std_logic_vector(188, 8),
50169 => conv_std_logic_vector(189, 8),
50170 => conv_std_logic_vector(190, 8),
50171 => conv_std_logic_vector(191, 8),
50172 => conv_std_logic_vector(191, 8),
50173 => conv_std_logic_vector(192, 8),
50174 => conv_std_logic_vector(193, 8),
50175 => conv_std_logic_vector(194, 8),
50176 => conv_std_logic_vector(0, 8),
50177 => conv_std_logic_vector(0, 8),
50178 => conv_std_logic_vector(1, 8),
50179 => conv_std_logic_vector(2, 8),
50180 => conv_std_logic_vector(3, 8),
50181 => conv_std_logic_vector(3, 8),
50182 => conv_std_logic_vector(4, 8),
50183 => conv_std_logic_vector(5, 8),
50184 => conv_std_logic_vector(6, 8),
50185 => conv_std_logic_vector(6, 8),
50186 => conv_std_logic_vector(7, 8),
50187 => conv_std_logic_vector(8, 8),
50188 => conv_std_logic_vector(9, 8),
50189 => conv_std_logic_vector(9, 8),
50190 => conv_std_logic_vector(10, 8),
50191 => conv_std_logic_vector(11, 8),
50192 => conv_std_logic_vector(12, 8),
50193 => conv_std_logic_vector(13, 8),
50194 => conv_std_logic_vector(13, 8),
50195 => conv_std_logic_vector(14, 8),
50196 => conv_std_logic_vector(15, 8),
50197 => conv_std_logic_vector(16, 8),
50198 => conv_std_logic_vector(16, 8),
50199 => conv_std_logic_vector(17, 8),
50200 => conv_std_logic_vector(18, 8),
50201 => conv_std_logic_vector(19, 8),
50202 => conv_std_logic_vector(19, 8),
50203 => conv_std_logic_vector(20, 8),
50204 => conv_std_logic_vector(21, 8),
50205 => conv_std_logic_vector(22, 8),
50206 => conv_std_logic_vector(22, 8),
50207 => conv_std_logic_vector(23, 8),
50208 => conv_std_logic_vector(24, 8),
50209 => conv_std_logic_vector(25, 8),
50210 => conv_std_logic_vector(26, 8),
50211 => conv_std_logic_vector(26, 8),
50212 => conv_std_logic_vector(27, 8),
50213 => conv_std_logic_vector(28, 8),
50214 => conv_std_logic_vector(29, 8),
50215 => conv_std_logic_vector(29, 8),
50216 => conv_std_logic_vector(30, 8),
50217 => conv_std_logic_vector(31, 8),
50218 => conv_std_logic_vector(32, 8),
50219 => conv_std_logic_vector(32, 8),
50220 => conv_std_logic_vector(33, 8),
50221 => conv_std_logic_vector(34, 8),
50222 => conv_std_logic_vector(35, 8),
50223 => conv_std_logic_vector(35, 8),
50224 => conv_std_logic_vector(36, 8),
50225 => conv_std_logic_vector(37, 8),
50226 => conv_std_logic_vector(38, 8),
50227 => conv_std_logic_vector(39, 8),
50228 => conv_std_logic_vector(39, 8),
50229 => conv_std_logic_vector(40, 8),
50230 => conv_std_logic_vector(41, 8),
50231 => conv_std_logic_vector(42, 8),
50232 => conv_std_logic_vector(42, 8),
50233 => conv_std_logic_vector(43, 8),
50234 => conv_std_logic_vector(44, 8),
50235 => conv_std_logic_vector(45, 8),
50236 => conv_std_logic_vector(45, 8),
50237 => conv_std_logic_vector(46, 8),
50238 => conv_std_logic_vector(47, 8),
50239 => conv_std_logic_vector(48, 8),
50240 => conv_std_logic_vector(49, 8),
50241 => conv_std_logic_vector(49, 8),
50242 => conv_std_logic_vector(50, 8),
50243 => conv_std_logic_vector(51, 8),
50244 => conv_std_logic_vector(52, 8),
50245 => conv_std_logic_vector(52, 8),
50246 => conv_std_logic_vector(53, 8),
50247 => conv_std_logic_vector(54, 8),
50248 => conv_std_logic_vector(55, 8),
50249 => conv_std_logic_vector(55, 8),
50250 => conv_std_logic_vector(56, 8),
50251 => conv_std_logic_vector(57, 8),
50252 => conv_std_logic_vector(58, 8),
50253 => conv_std_logic_vector(58, 8),
50254 => conv_std_logic_vector(59, 8),
50255 => conv_std_logic_vector(60, 8),
50256 => conv_std_logic_vector(61, 8),
50257 => conv_std_logic_vector(62, 8),
50258 => conv_std_logic_vector(62, 8),
50259 => conv_std_logic_vector(63, 8),
50260 => conv_std_logic_vector(64, 8),
50261 => conv_std_logic_vector(65, 8),
50262 => conv_std_logic_vector(65, 8),
50263 => conv_std_logic_vector(66, 8),
50264 => conv_std_logic_vector(67, 8),
50265 => conv_std_logic_vector(68, 8),
50266 => conv_std_logic_vector(68, 8),
50267 => conv_std_logic_vector(69, 8),
50268 => conv_std_logic_vector(70, 8),
50269 => conv_std_logic_vector(71, 8),
50270 => conv_std_logic_vector(71, 8),
50271 => conv_std_logic_vector(72, 8),
50272 => conv_std_logic_vector(73, 8),
50273 => conv_std_logic_vector(74, 8),
50274 => conv_std_logic_vector(75, 8),
50275 => conv_std_logic_vector(75, 8),
50276 => conv_std_logic_vector(76, 8),
50277 => conv_std_logic_vector(77, 8),
50278 => conv_std_logic_vector(78, 8),
50279 => conv_std_logic_vector(78, 8),
50280 => conv_std_logic_vector(79, 8),
50281 => conv_std_logic_vector(80, 8),
50282 => conv_std_logic_vector(81, 8),
50283 => conv_std_logic_vector(81, 8),
50284 => conv_std_logic_vector(82, 8),
50285 => conv_std_logic_vector(83, 8),
50286 => conv_std_logic_vector(84, 8),
50287 => conv_std_logic_vector(84, 8),
50288 => conv_std_logic_vector(85, 8),
50289 => conv_std_logic_vector(86, 8),
50290 => conv_std_logic_vector(87, 8),
50291 => conv_std_logic_vector(88, 8),
50292 => conv_std_logic_vector(88, 8),
50293 => conv_std_logic_vector(89, 8),
50294 => conv_std_logic_vector(90, 8),
50295 => conv_std_logic_vector(91, 8),
50296 => conv_std_logic_vector(91, 8),
50297 => conv_std_logic_vector(92, 8),
50298 => conv_std_logic_vector(93, 8),
50299 => conv_std_logic_vector(94, 8),
50300 => conv_std_logic_vector(94, 8),
50301 => conv_std_logic_vector(95, 8),
50302 => conv_std_logic_vector(96, 8),
50303 => conv_std_logic_vector(97, 8),
50304 => conv_std_logic_vector(98, 8),
50305 => conv_std_logic_vector(98, 8),
50306 => conv_std_logic_vector(99, 8),
50307 => conv_std_logic_vector(100, 8),
50308 => conv_std_logic_vector(101, 8),
50309 => conv_std_logic_vector(101, 8),
50310 => conv_std_logic_vector(102, 8),
50311 => conv_std_logic_vector(103, 8),
50312 => conv_std_logic_vector(104, 8),
50313 => conv_std_logic_vector(104, 8),
50314 => conv_std_logic_vector(105, 8),
50315 => conv_std_logic_vector(106, 8),
50316 => conv_std_logic_vector(107, 8),
50317 => conv_std_logic_vector(107, 8),
50318 => conv_std_logic_vector(108, 8),
50319 => conv_std_logic_vector(109, 8),
50320 => conv_std_logic_vector(110, 8),
50321 => conv_std_logic_vector(111, 8),
50322 => conv_std_logic_vector(111, 8),
50323 => conv_std_logic_vector(112, 8),
50324 => conv_std_logic_vector(113, 8),
50325 => conv_std_logic_vector(114, 8),
50326 => conv_std_logic_vector(114, 8),
50327 => conv_std_logic_vector(115, 8),
50328 => conv_std_logic_vector(116, 8),
50329 => conv_std_logic_vector(117, 8),
50330 => conv_std_logic_vector(117, 8),
50331 => conv_std_logic_vector(118, 8),
50332 => conv_std_logic_vector(119, 8),
50333 => conv_std_logic_vector(120, 8),
50334 => conv_std_logic_vector(120, 8),
50335 => conv_std_logic_vector(121, 8),
50336 => conv_std_logic_vector(122, 8),
50337 => conv_std_logic_vector(123, 8),
50338 => conv_std_logic_vector(124, 8),
50339 => conv_std_logic_vector(124, 8),
50340 => conv_std_logic_vector(125, 8),
50341 => conv_std_logic_vector(126, 8),
50342 => conv_std_logic_vector(127, 8),
50343 => conv_std_logic_vector(127, 8),
50344 => conv_std_logic_vector(128, 8),
50345 => conv_std_logic_vector(129, 8),
50346 => conv_std_logic_vector(130, 8),
50347 => conv_std_logic_vector(130, 8),
50348 => conv_std_logic_vector(131, 8),
50349 => conv_std_logic_vector(132, 8),
50350 => conv_std_logic_vector(133, 8),
50351 => conv_std_logic_vector(133, 8),
50352 => conv_std_logic_vector(134, 8),
50353 => conv_std_logic_vector(135, 8),
50354 => conv_std_logic_vector(136, 8),
50355 => conv_std_logic_vector(137, 8),
50356 => conv_std_logic_vector(137, 8),
50357 => conv_std_logic_vector(138, 8),
50358 => conv_std_logic_vector(139, 8),
50359 => conv_std_logic_vector(140, 8),
50360 => conv_std_logic_vector(140, 8),
50361 => conv_std_logic_vector(141, 8),
50362 => conv_std_logic_vector(142, 8),
50363 => conv_std_logic_vector(143, 8),
50364 => conv_std_logic_vector(143, 8),
50365 => conv_std_logic_vector(144, 8),
50366 => conv_std_logic_vector(145, 8),
50367 => conv_std_logic_vector(146, 8),
50368 => conv_std_logic_vector(147, 8),
50369 => conv_std_logic_vector(147, 8),
50370 => conv_std_logic_vector(148, 8),
50371 => conv_std_logic_vector(149, 8),
50372 => conv_std_logic_vector(150, 8),
50373 => conv_std_logic_vector(150, 8),
50374 => conv_std_logic_vector(151, 8),
50375 => conv_std_logic_vector(152, 8),
50376 => conv_std_logic_vector(153, 8),
50377 => conv_std_logic_vector(153, 8),
50378 => conv_std_logic_vector(154, 8),
50379 => conv_std_logic_vector(155, 8),
50380 => conv_std_logic_vector(156, 8),
50381 => conv_std_logic_vector(156, 8),
50382 => conv_std_logic_vector(157, 8),
50383 => conv_std_logic_vector(158, 8),
50384 => conv_std_logic_vector(159, 8),
50385 => conv_std_logic_vector(160, 8),
50386 => conv_std_logic_vector(160, 8),
50387 => conv_std_logic_vector(161, 8),
50388 => conv_std_logic_vector(162, 8),
50389 => conv_std_logic_vector(163, 8),
50390 => conv_std_logic_vector(163, 8),
50391 => conv_std_logic_vector(164, 8),
50392 => conv_std_logic_vector(165, 8),
50393 => conv_std_logic_vector(166, 8),
50394 => conv_std_logic_vector(166, 8),
50395 => conv_std_logic_vector(167, 8),
50396 => conv_std_logic_vector(168, 8),
50397 => conv_std_logic_vector(169, 8),
50398 => conv_std_logic_vector(169, 8),
50399 => conv_std_logic_vector(170, 8),
50400 => conv_std_logic_vector(171, 8),
50401 => conv_std_logic_vector(172, 8),
50402 => conv_std_logic_vector(173, 8),
50403 => conv_std_logic_vector(173, 8),
50404 => conv_std_logic_vector(174, 8),
50405 => conv_std_logic_vector(175, 8),
50406 => conv_std_logic_vector(176, 8),
50407 => conv_std_logic_vector(176, 8),
50408 => conv_std_logic_vector(177, 8),
50409 => conv_std_logic_vector(178, 8),
50410 => conv_std_logic_vector(179, 8),
50411 => conv_std_logic_vector(179, 8),
50412 => conv_std_logic_vector(180, 8),
50413 => conv_std_logic_vector(181, 8),
50414 => conv_std_logic_vector(182, 8),
50415 => conv_std_logic_vector(182, 8),
50416 => conv_std_logic_vector(183, 8),
50417 => conv_std_logic_vector(184, 8),
50418 => conv_std_logic_vector(185, 8),
50419 => conv_std_logic_vector(186, 8),
50420 => conv_std_logic_vector(186, 8),
50421 => conv_std_logic_vector(187, 8),
50422 => conv_std_logic_vector(188, 8),
50423 => conv_std_logic_vector(189, 8),
50424 => conv_std_logic_vector(189, 8),
50425 => conv_std_logic_vector(190, 8),
50426 => conv_std_logic_vector(191, 8),
50427 => conv_std_logic_vector(192, 8),
50428 => conv_std_logic_vector(192, 8),
50429 => conv_std_logic_vector(193, 8),
50430 => conv_std_logic_vector(194, 8),
50431 => conv_std_logic_vector(195, 8),
50432 => conv_std_logic_vector(0, 8),
50433 => conv_std_logic_vector(0, 8),
50434 => conv_std_logic_vector(1, 8),
50435 => conv_std_logic_vector(2, 8),
50436 => conv_std_logic_vector(3, 8),
50437 => conv_std_logic_vector(3, 8),
50438 => conv_std_logic_vector(4, 8),
50439 => conv_std_logic_vector(5, 8),
50440 => conv_std_logic_vector(6, 8),
50441 => conv_std_logic_vector(6, 8),
50442 => conv_std_logic_vector(7, 8),
50443 => conv_std_logic_vector(8, 8),
50444 => conv_std_logic_vector(9, 8),
50445 => conv_std_logic_vector(10, 8),
50446 => conv_std_logic_vector(10, 8),
50447 => conv_std_logic_vector(11, 8),
50448 => conv_std_logic_vector(12, 8),
50449 => conv_std_logic_vector(13, 8),
50450 => conv_std_logic_vector(13, 8),
50451 => conv_std_logic_vector(14, 8),
50452 => conv_std_logic_vector(15, 8),
50453 => conv_std_logic_vector(16, 8),
50454 => conv_std_logic_vector(16, 8),
50455 => conv_std_logic_vector(17, 8),
50456 => conv_std_logic_vector(18, 8),
50457 => conv_std_logic_vector(19, 8),
50458 => conv_std_logic_vector(20, 8),
50459 => conv_std_logic_vector(20, 8),
50460 => conv_std_logic_vector(21, 8),
50461 => conv_std_logic_vector(22, 8),
50462 => conv_std_logic_vector(23, 8),
50463 => conv_std_logic_vector(23, 8),
50464 => conv_std_logic_vector(24, 8),
50465 => conv_std_logic_vector(25, 8),
50466 => conv_std_logic_vector(26, 8),
50467 => conv_std_logic_vector(26, 8),
50468 => conv_std_logic_vector(27, 8),
50469 => conv_std_logic_vector(28, 8),
50470 => conv_std_logic_vector(29, 8),
50471 => conv_std_logic_vector(30, 8),
50472 => conv_std_logic_vector(30, 8),
50473 => conv_std_logic_vector(31, 8),
50474 => conv_std_logic_vector(32, 8),
50475 => conv_std_logic_vector(33, 8),
50476 => conv_std_logic_vector(33, 8),
50477 => conv_std_logic_vector(34, 8),
50478 => conv_std_logic_vector(35, 8),
50479 => conv_std_logic_vector(36, 8),
50480 => conv_std_logic_vector(36, 8),
50481 => conv_std_logic_vector(37, 8),
50482 => conv_std_logic_vector(38, 8),
50483 => conv_std_logic_vector(39, 8),
50484 => conv_std_logic_vector(40, 8),
50485 => conv_std_logic_vector(40, 8),
50486 => conv_std_logic_vector(41, 8),
50487 => conv_std_logic_vector(42, 8),
50488 => conv_std_logic_vector(43, 8),
50489 => conv_std_logic_vector(43, 8),
50490 => conv_std_logic_vector(44, 8),
50491 => conv_std_logic_vector(45, 8),
50492 => conv_std_logic_vector(46, 8),
50493 => conv_std_logic_vector(46, 8),
50494 => conv_std_logic_vector(47, 8),
50495 => conv_std_logic_vector(48, 8),
50496 => conv_std_logic_vector(49, 8),
50497 => conv_std_logic_vector(50, 8),
50498 => conv_std_logic_vector(50, 8),
50499 => conv_std_logic_vector(51, 8),
50500 => conv_std_logic_vector(52, 8),
50501 => conv_std_logic_vector(53, 8),
50502 => conv_std_logic_vector(53, 8),
50503 => conv_std_logic_vector(54, 8),
50504 => conv_std_logic_vector(55, 8),
50505 => conv_std_logic_vector(56, 8),
50506 => conv_std_logic_vector(56, 8),
50507 => conv_std_logic_vector(57, 8),
50508 => conv_std_logic_vector(58, 8),
50509 => conv_std_logic_vector(59, 8),
50510 => conv_std_logic_vector(60, 8),
50511 => conv_std_logic_vector(60, 8),
50512 => conv_std_logic_vector(61, 8),
50513 => conv_std_logic_vector(62, 8),
50514 => conv_std_logic_vector(63, 8),
50515 => conv_std_logic_vector(63, 8),
50516 => conv_std_logic_vector(64, 8),
50517 => conv_std_logic_vector(65, 8),
50518 => conv_std_logic_vector(66, 8),
50519 => conv_std_logic_vector(66, 8),
50520 => conv_std_logic_vector(67, 8),
50521 => conv_std_logic_vector(68, 8),
50522 => conv_std_logic_vector(69, 8),
50523 => conv_std_logic_vector(70, 8),
50524 => conv_std_logic_vector(70, 8),
50525 => conv_std_logic_vector(71, 8),
50526 => conv_std_logic_vector(72, 8),
50527 => conv_std_logic_vector(73, 8),
50528 => conv_std_logic_vector(73, 8),
50529 => conv_std_logic_vector(74, 8),
50530 => conv_std_logic_vector(75, 8),
50531 => conv_std_logic_vector(76, 8),
50532 => conv_std_logic_vector(76, 8),
50533 => conv_std_logic_vector(77, 8),
50534 => conv_std_logic_vector(78, 8),
50535 => conv_std_logic_vector(79, 8),
50536 => conv_std_logic_vector(80, 8),
50537 => conv_std_logic_vector(80, 8),
50538 => conv_std_logic_vector(81, 8),
50539 => conv_std_logic_vector(82, 8),
50540 => conv_std_logic_vector(83, 8),
50541 => conv_std_logic_vector(83, 8),
50542 => conv_std_logic_vector(84, 8),
50543 => conv_std_logic_vector(85, 8),
50544 => conv_std_logic_vector(86, 8),
50545 => conv_std_logic_vector(86, 8),
50546 => conv_std_logic_vector(87, 8),
50547 => conv_std_logic_vector(88, 8),
50548 => conv_std_logic_vector(89, 8),
50549 => conv_std_logic_vector(90, 8),
50550 => conv_std_logic_vector(90, 8),
50551 => conv_std_logic_vector(91, 8),
50552 => conv_std_logic_vector(92, 8),
50553 => conv_std_logic_vector(93, 8),
50554 => conv_std_logic_vector(93, 8),
50555 => conv_std_logic_vector(94, 8),
50556 => conv_std_logic_vector(95, 8),
50557 => conv_std_logic_vector(96, 8),
50558 => conv_std_logic_vector(96, 8),
50559 => conv_std_logic_vector(97, 8),
50560 => conv_std_logic_vector(98, 8),
50561 => conv_std_logic_vector(99, 8),
50562 => conv_std_logic_vector(100, 8),
50563 => conv_std_logic_vector(100, 8),
50564 => conv_std_logic_vector(101, 8),
50565 => conv_std_logic_vector(102, 8),
50566 => conv_std_logic_vector(103, 8),
50567 => conv_std_logic_vector(103, 8),
50568 => conv_std_logic_vector(104, 8),
50569 => conv_std_logic_vector(105, 8),
50570 => conv_std_logic_vector(106, 8),
50571 => conv_std_logic_vector(106, 8),
50572 => conv_std_logic_vector(107, 8),
50573 => conv_std_logic_vector(108, 8),
50574 => conv_std_logic_vector(109, 8),
50575 => conv_std_logic_vector(110, 8),
50576 => conv_std_logic_vector(110, 8),
50577 => conv_std_logic_vector(111, 8),
50578 => conv_std_logic_vector(112, 8),
50579 => conv_std_logic_vector(113, 8),
50580 => conv_std_logic_vector(113, 8),
50581 => conv_std_logic_vector(114, 8),
50582 => conv_std_logic_vector(115, 8),
50583 => conv_std_logic_vector(116, 8),
50584 => conv_std_logic_vector(116, 8),
50585 => conv_std_logic_vector(117, 8),
50586 => conv_std_logic_vector(118, 8),
50587 => conv_std_logic_vector(119, 8),
50588 => conv_std_logic_vector(120, 8),
50589 => conv_std_logic_vector(120, 8),
50590 => conv_std_logic_vector(121, 8),
50591 => conv_std_logic_vector(122, 8),
50592 => conv_std_logic_vector(123, 8),
50593 => conv_std_logic_vector(123, 8),
50594 => conv_std_logic_vector(124, 8),
50595 => conv_std_logic_vector(125, 8),
50596 => conv_std_logic_vector(126, 8),
50597 => conv_std_logic_vector(126, 8),
50598 => conv_std_logic_vector(127, 8),
50599 => conv_std_logic_vector(128, 8),
50600 => conv_std_logic_vector(129, 8),
50601 => conv_std_logic_vector(130, 8),
50602 => conv_std_logic_vector(130, 8),
50603 => conv_std_logic_vector(131, 8),
50604 => conv_std_logic_vector(132, 8),
50605 => conv_std_logic_vector(133, 8),
50606 => conv_std_logic_vector(133, 8),
50607 => conv_std_logic_vector(134, 8),
50608 => conv_std_logic_vector(135, 8),
50609 => conv_std_logic_vector(136, 8),
50610 => conv_std_logic_vector(136, 8),
50611 => conv_std_logic_vector(137, 8),
50612 => conv_std_logic_vector(138, 8),
50613 => conv_std_logic_vector(139, 8),
50614 => conv_std_logic_vector(140, 8),
50615 => conv_std_logic_vector(140, 8),
50616 => conv_std_logic_vector(141, 8),
50617 => conv_std_logic_vector(142, 8),
50618 => conv_std_logic_vector(143, 8),
50619 => conv_std_logic_vector(143, 8),
50620 => conv_std_logic_vector(144, 8),
50621 => conv_std_logic_vector(145, 8),
50622 => conv_std_logic_vector(146, 8),
50623 => conv_std_logic_vector(146, 8),
50624 => conv_std_logic_vector(147, 8),
50625 => conv_std_logic_vector(148, 8),
50626 => conv_std_logic_vector(149, 8),
50627 => conv_std_logic_vector(150, 8),
50628 => conv_std_logic_vector(150, 8),
50629 => conv_std_logic_vector(151, 8),
50630 => conv_std_logic_vector(152, 8),
50631 => conv_std_logic_vector(153, 8),
50632 => conv_std_logic_vector(153, 8),
50633 => conv_std_logic_vector(154, 8),
50634 => conv_std_logic_vector(155, 8),
50635 => conv_std_logic_vector(156, 8),
50636 => conv_std_logic_vector(156, 8),
50637 => conv_std_logic_vector(157, 8),
50638 => conv_std_logic_vector(158, 8),
50639 => conv_std_logic_vector(159, 8),
50640 => conv_std_logic_vector(160, 8),
50641 => conv_std_logic_vector(160, 8),
50642 => conv_std_logic_vector(161, 8),
50643 => conv_std_logic_vector(162, 8),
50644 => conv_std_logic_vector(163, 8),
50645 => conv_std_logic_vector(163, 8),
50646 => conv_std_logic_vector(164, 8),
50647 => conv_std_logic_vector(165, 8),
50648 => conv_std_logic_vector(166, 8),
50649 => conv_std_logic_vector(166, 8),
50650 => conv_std_logic_vector(167, 8),
50651 => conv_std_logic_vector(168, 8),
50652 => conv_std_logic_vector(169, 8),
50653 => conv_std_logic_vector(170, 8),
50654 => conv_std_logic_vector(170, 8),
50655 => conv_std_logic_vector(171, 8),
50656 => conv_std_logic_vector(172, 8),
50657 => conv_std_logic_vector(173, 8),
50658 => conv_std_logic_vector(173, 8),
50659 => conv_std_logic_vector(174, 8),
50660 => conv_std_logic_vector(175, 8),
50661 => conv_std_logic_vector(176, 8),
50662 => conv_std_logic_vector(176, 8),
50663 => conv_std_logic_vector(177, 8),
50664 => conv_std_logic_vector(178, 8),
50665 => conv_std_logic_vector(179, 8),
50666 => conv_std_logic_vector(180, 8),
50667 => conv_std_logic_vector(180, 8),
50668 => conv_std_logic_vector(181, 8),
50669 => conv_std_logic_vector(182, 8),
50670 => conv_std_logic_vector(183, 8),
50671 => conv_std_logic_vector(183, 8),
50672 => conv_std_logic_vector(184, 8),
50673 => conv_std_logic_vector(185, 8),
50674 => conv_std_logic_vector(186, 8),
50675 => conv_std_logic_vector(186, 8),
50676 => conv_std_logic_vector(187, 8),
50677 => conv_std_logic_vector(188, 8),
50678 => conv_std_logic_vector(189, 8),
50679 => conv_std_logic_vector(190, 8),
50680 => conv_std_logic_vector(190, 8),
50681 => conv_std_logic_vector(191, 8),
50682 => conv_std_logic_vector(192, 8),
50683 => conv_std_logic_vector(193, 8),
50684 => conv_std_logic_vector(193, 8),
50685 => conv_std_logic_vector(194, 8),
50686 => conv_std_logic_vector(195, 8),
50687 => conv_std_logic_vector(196, 8),
50688 => conv_std_logic_vector(0, 8),
50689 => conv_std_logic_vector(0, 8),
50690 => conv_std_logic_vector(1, 8),
50691 => conv_std_logic_vector(2, 8),
50692 => conv_std_logic_vector(3, 8),
50693 => conv_std_logic_vector(3, 8),
50694 => conv_std_logic_vector(4, 8),
50695 => conv_std_logic_vector(5, 8),
50696 => conv_std_logic_vector(6, 8),
50697 => conv_std_logic_vector(6, 8),
50698 => conv_std_logic_vector(7, 8),
50699 => conv_std_logic_vector(8, 8),
50700 => conv_std_logic_vector(9, 8),
50701 => conv_std_logic_vector(10, 8),
50702 => conv_std_logic_vector(10, 8),
50703 => conv_std_logic_vector(11, 8),
50704 => conv_std_logic_vector(12, 8),
50705 => conv_std_logic_vector(13, 8),
50706 => conv_std_logic_vector(13, 8),
50707 => conv_std_logic_vector(14, 8),
50708 => conv_std_logic_vector(15, 8),
50709 => conv_std_logic_vector(16, 8),
50710 => conv_std_logic_vector(17, 8),
50711 => conv_std_logic_vector(17, 8),
50712 => conv_std_logic_vector(18, 8),
50713 => conv_std_logic_vector(19, 8),
50714 => conv_std_logic_vector(20, 8),
50715 => conv_std_logic_vector(20, 8),
50716 => conv_std_logic_vector(21, 8),
50717 => conv_std_logic_vector(22, 8),
50718 => conv_std_logic_vector(23, 8),
50719 => conv_std_logic_vector(23, 8),
50720 => conv_std_logic_vector(24, 8),
50721 => conv_std_logic_vector(25, 8),
50722 => conv_std_logic_vector(26, 8),
50723 => conv_std_logic_vector(27, 8),
50724 => conv_std_logic_vector(27, 8),
50725 => conv_std_logic_vector(28, 8),
50726 => conv_std_logic_vector(29, 8),
50727 => conv_std_logic_vector(30, 8),
50728 => conv_std_logic_vector(30, 8),
50729 => conv_std_logic_vector(31, 8),
50730 => conv_std_logic_vector(32, 8),
50731 => conv_std_logic_vector(33, 8),
50732 => conv_std_logic_vector(34, 8),
50733 => conv_std_logic_vector(34, 8),
50734 => conv_std_logic_vector(35, 8),
50735 => conv_std_logic_vector(36, 8),
50736 => conv_std_logic_vector(37, 8),
50737 => conv_std_logic_vector(37, 8),
50738 => conv_std_logic_vector(38, 8),
50739 => conv_std_logic_vector(39, 8),
50740 => conv_std_logic_vector(40, 8),
50741 => conv_std_logic_vector(40, 8),
50742 => conv_std_logic_vector(41, 8),
50743 => conv_std_logic_vector(42, 8),
50744 => conv_std_logic_vector(43, 8),
50745 => conv_std_logic_vector(44, 8),
50746 => conv_std_logic_vector(44, 8),
50747 => conv_std_logic_vector(45, 8),
50748 => conv_std_logic_vector(46, 8),
50749 => conv_std_logic_vector(47, 8),
50750 => conv_std_logic_vector(47, 8),
50751 => conv_std_logic_vector(48, 8),
50752 => conv_std_logic_vector(49, 8),
50753 => conv_std_logic_vector(50, 8),
50754 => conv_std_logic_vector(51, 8),
50755 => conv_std_logic_vector(51, 8),
50756 => conv_std_logic_vector(52, 8),
50757 => conv_std_logic_vector(53, 8),
50758 => conv_std_logic_vector(54, 8),
50759 => conv_std_logic_vector(54, 8),
50760 => conv_std_logic_vector(55, 8),
50761 => conv_std_logic_vector(56, 8),
50762 => conv_std_logic_vector(57, 8),
50763 => conv_std_logic_vector(58, 8),
50764 => conv_std_logic_vector(58, 8),
50765 => conv_std_logic_vector(59, 8),
50766 => conv_std_logic_vector(60, 8),
50767 => conv_std_logic_vector(61, 8),
50768 => conv_std_logic_vector(61, 8),
50769 => conv_std_logic_vector(62, 8),
50770 => conv_std_logic_vector(63, 8),
50771 => conv_std_logic_vector(64, 8),
50772 => conv_std_logic_vector(64, 8),
50773 => conv_std_logic_vector(65, 8),
50774 => conv_std_logic_vector(66, 8),
50775 => conv_std_logic_vector(67, 8),
50776 => conv_std_logic_vector(68, 8),
50777 => conv_std_logic_vector(68, 8),
50778 => conv_std_logic_vector(69, 8),
50779 => conv_std_logic_vector(70, 8),
50780 => conv_std_logic_vector(71, 8),
50781 => conv_std_logic_vector(71, 8),
50782 => conv_std_logic_vector(72, 8),
50783 => conv_std_logic_vector(73, 8),
50784 => conv_std_logic_vector(74, 8),
50785 => conv_std_logic_vector(75, 8),
50786 => conv_std_logic_vector(75, 8),
50787 => conv_std_logic_vector(76, 8),
50788 => conv_std_logic_vector(77, 8),
50789 => conv_std_logic_vector(78, 8),
50790 => conv_std_logic_vector(78, 8),
50791 => conv_std_logic_vector(79, 8),
50792 => conv_std_logic_vector(80, 8),
50793 => conv_std_logic_vector(81, 8),
50794 => conv_std_logic_vector(81, 8),
50795 => conv_std_logic_vector(82, 8),
50796 => conv_std_logic_vector(83, 8),
50797 => conv_std_logic_vector(84, 8),
50798 => conv_std_logic_vector(85, 8),
50799 => conv_std_logic_vector(85, 8),
50800 => conv_std_logic_vector(86, 8),
50801 => conv_std_logic_vector(87, 8),
50802 => conv_std_logic_vector(88, 8),
50803 => conv_std_logic_vector(88, 8),
50804 => conv_std_logic_vector(89, 8),
50805 => conv_std_logic_vector(90, 8),
50806 => conv_std_logic_vector(91, 8),
50807 => conv_std_logic_vector(92, 8),
50808 => conv_std_logic_vector(92, 8),
50809 => conv_std_logic_vector(93, 8),
50810 => conv_std_logic_vector(94, 8),
50811 => conv_std_logic_vector(95, 8),
50812 => conv_std_logic_vector(95, 8),
50813 => conv_std_logic_vector(96, 8),
50814 => conv_std_logic_vector(97, 8),
50815 => conv_std_logic_vector(98, 8),
50816 => conv_std_logic_vector(99, 8),
50817 => conv_std_logic_vector(99, 8),
50818 => conv_std_logic_vector(100, 8),
50819 => conv_std_logic_vector(101, 8),
50820 => conv_std_logic_vector(102, 8),
50821 => conv_std_logic_vector(102, 8),
50822 => conv_std_logic_vector(103, 8),
50823 => conv_std_logic_vector(104, 8),
50824 => conv_std_logic_vector(105, 8),
50825 => conv_std_logic_vector(105, 8),
50826 => conv_std_logic_vector(106, 8),
50827 => conv_std_logic_vector(107, 8),
50828 => conv_std_logic_vector(108, 8),
50829 => conv_std_logic_vector(109, 8),
50830 => conv_std_logic_vector(109, 8),
50831 => conv_std_logic_vector(110, 8),
50832 => conv_std_logic_vector(111, 8),
50833 => conv_std_logic_vector(112, 8),
50834 => conv_std_logic_vector(112, 8),
50835 => conv_std_logic_vector(113, 8),
50836 => conv_std_logic_vector(114, 8),
50837 => conv_std_logic_vector(115, 8),
50838 => conv_std_logic_vector(116, 8),
50839 => conv_std_logic_vector(116, 8),
50840 => conv_std_logic_vector(117, 8),
50841 => conv_std_logic_vector(118, 8),
50842 => conv_std_logic_vector(119, 8),
50843 => conv_std_logic_vector(119, 8),
50844 => conv_std_logic_vector(120, 8),
50845 => conv_std_logic_vector(121, 8),
50846 => conv_std_logic_vector(122, 8),
50847 => conv_std_logic_vector(122, 8),
50848 => conv_std_logic_vector(123, 8),
50849 => conv_std_logic_vector(124, 8),
50850 => conv_std_logic_vector(125, 8),
50851 => conv_std_logic_vector(126, 8),
50852 => conv_std_logic_vector(126, 8),
50853 => conv_std_logic_vector(127, 8),
50854 => conv_std_logic_vector(128, 8),
50855 => conv_std_logic_vector(129, 8),
50856 => conv_std_logic_vector(129, 8),
50857 => conv_std_logic_vector(130, 8),
50858 => conv_std_logic_vector(131, 8),
50859 => conv_std_logic_vector(132, 8),
50860 => conv_std_logic_vector(133, 8),
50861 => conv_std_logic_vector(133, 8),
50862 => conv_std_logic_vector(134, 8),
50863 => conv_std_logic_vector(135, 8),
50864 => conv_std_logic_vector(136, 8),
50865 => conv_std_logic_vector(136, 8),
50866 => conv_std_logic_vector(137, 8),
50867 => conv_std_logic_vector(138, 8),
50868 => conv_std_logic_vector(139, 8),
50869 => conv_std_logic_vector(139, 8),
50870 => conv_std_logic_vector(140, 8),
50871 => conv_std_logic_vector(141, 8),
50872 => conv_std_logic_vector(142, 8),
50873 => conv_std_logic_vector(143, 8),
50874 => conv_std_logic_vector(143, 8),
50875 => conv_std_logic_vector(144, 8),
50876 => conv_std_logic_vector(145, 8),
50877 => conv_std_logic_vector(146, 8),
50878 => conv_std_logic_vector(146, 8),
50879 => conv_std_logic_vector(147, 8),
50880 => conv_std_logic_vector(148, 8),
50881 => conv_std_logic_vector(149, 8),
50882 => conv_std_logic_vector(150, 8),
50883 => conv_std_logic_vector(150, 8),
50884 => conv_std_logic_vector(151, 8),
50885 => conv_std_logic_vector(152, 8),
50886 => conv_std_logic_vector(153, 8),
50887 => conv_std_logic_vector(153, 8),
50888 => conv_std_logic_vector(154, 8),
50889 => conv_std_logic_vector(155, 8),
50890 => conv_std_logic_vector(156, 8),
50891 => conv_std_logic_vector(157, 8),
50892 => conv_std_logic_vector(157, 8),
50893 => conv_std_logic_vector(158, 8),
50894 => conv_std_logic_vector(159, 8),
50895 => conv_std_logic_vector(160, 8),
50896 => conv_std_logic_vector(160, 8),
50897 => conv_std_logic_vector(161, 8),
50898 => conv_std_logic_vector(162, 8),
50899 => conv_std_logic_vector(163, 8),
50900 => conv_std_logic_vector(163, 8),
50901 => conv_std_logic_vector(164, 8),
50902 => conv_std_logic_vector(165, 8),
50903 => conv_std_logic_vector(166, 8),
50904 => conv_std_logic_vector(167, 8),
50905 => conv_std_logic_vector(167, 8),
50906 => conv_std_logic_vector(168, 8),
50907 => conv_std_logic_vector(169, 8),
50908 => conv_std_logic_vector(170, 8),
50909 => conv_std_logic_vector(170, 8),
50910 => conv_std_logic_vector(171, 8),
50911 => conv_std_logic_vector(172, 8),
50912 => conv_std_logic_vector(173, 8),
50913 => conv_std_logic_vector(174, 8),
50914 => conv_std_logic_vector(174, 8),
50915 => conv_std_logic_vector(175, 8),
50916 => conv_std_logic_vector(176, 8),
50917 => conv_std_logic_vector(177, 8),
50918 => conv_std_logic_vector(177, 8),
50919 => conv_std_logic_vector(178, 8),
50920 => conv_std_logic_vector(179, 8),
50921 => conv_std_logic_vector(180, 8),
50922 => conv_std_logic_vector(180, 8),
50923 => conv_std_logic_vector(181, 8),
50924 => conv_std_logic_vector(182, 8),
50925 => conv_std_logic_vector(183, 8),
50926 => conv_std_logic_vector(184, 8),
50927 => conv_std_logic_vector(184, 8),
50928 => conv_std_logic_vector(185, 8),
50929 => conv_std_logic_vector(186, 8),
50930 => conv_std_logic_vector(187, 8),
50931 => conv_std_logic_vector(187, 8),
50932 => conv_std_logic_vector(188, 8),
50933 => conv_std_logic_vector(189, 8),
50934 => conv_std_logic_vector(190, 8),
50935 => conv_std_logic_vector(191, 8),
50936 => conv_std_logic_vector(191, 8),
50937 => conv_std_logic_vector(192, 8),
50938 => conv_std_logic_vector(193, 8),
50939 => conv_std_logic_vector(194, 8),
50940 => conv_std_logic_vector(194, 8),
50941 => conv_std_logic_vector(195, 8),
50942 => conv_std_logic_vector(196, 8),
50943 => conv_std_logic_vector(197, 8),
50944 => conv_std_logic_vector(0, 8),
50945 => conv_std_logic_vector(0, 8),
50946 => conv_std_logic_vector(1, 8),
50947 => conv_std_logic_vector(2, 8),
50948 => conv_std_logic_vector(3, 8),
50949 => conv_std_logic_vector(3, 8),
50950 => conv_std_logic_vector(4, 8),
50951 => conv_std_logic_vector(5, 8),
50952 => conv_std_logic_vector(6, 8),
50953 => conv_std_logic_vector(6, 8),
50954 => conv_std_logic_vector(7, 8),
50955 => conv_std_logic_vector(8, 8),
50956 => conv_std_logic_vector(9, 8),
50957 => conv_std_logic_vector(10, 8),
50958 => conv_std_logic_vector(10, 8),
50959 => conv_std_logic_vector(11, 8),
50960 => conv_std_logic_vector(12, 8),
50961 => conv_std_logic_vector(13, 8),
50962 => conv_std_logic_vector(13, 8),
50963 => conv_std_logic_vector(14, 8),
50964 => conv_std_logic_vector(15, 8),
50965 => conv_std_logic_vector(16, 8),
50966 => conv_std_logic_vector(17, 8),
50967 => conv_std_logic_vector(17, 8),
50968 => conv_std_logic_vector(18, 8),
50969 => conv_std_logic_vector(19, 8),
50970 => conv_std_logic_vector(20, 8),
50971 => conv_std_logic_vector(20, 8),
50972 => conv_std_logic_vector(21, 8),
50973 => conv_std_logic_vector(22, 8),
50974 => conv_std_logic_vector(23, 8),
50975 => conv_std_logic_vector(24, 8),
50976 => conv_std_logic_vector(24, 8),
50977 => conv_std_logic_vector(25, 8),
50978 => conv_std_logic_vector(26, 8),
50979 => conv_std_logic_vector(27, 8),
50980 => conv_std_logic_vector(27, 8),
50981 => conv_std_logic_vector(28, 8),
50982 => conv_std_logic_vector(29, 8),
50983 => conv_std_logic_vector(30, 8),
50984 => conv_std_logic_vector(31, 8),
50985 => conv_std_logic_vector(31, 8),
50986 => conv_std_logic_vector(32, 8),
50987 => conv_std_logic_vector(33, 8),
50988 => conv_std_logic_vector(34, 8),
50989 => conv_std_logic_vector(34, 8),
50990 => conv_std_logic_vector(35, 8),
50991 => conv_std_logic_vector(36, 8),
50992 => conv_std_logic_vector(37, 8),
50993 => conv_std_logic_vector(38, 8),
50994 => conv_std_logic_vector(38, 8),
50995 => conv_std_logic_vector(39, 8),
50996 => conv_std_logic_vector(40, 8),
50997 => conv_std_logic_vector(41, 8),
50998 => conv_std_logic_vector(41, 8),
50999 => conv_std_logic_vector(42, 8),
51000 => conv_std_logic_vector(43, 8),
51001 => conv_std_logic_vector(44, 8),
51002 => conv_std_logic_vector(45, 8),
51003 => conv_std_logic_vector(45, 8),
51004 => conv_std_logic_vector(46, 8),
51005 => conv_std_logic_vector(47, 8),
51006 => conv_std_logic_vector(48, 8),
51007 => conv_std_logic_vector(48, 8),
51008 => conv_std_logic_vector(49, 8),
51009 => conv_std_logic_vector(50, 8),
51010 => conv_std_logic_vector(51, 8),
51011 => conv_std_logic_vector(52, 8),
51012 => conv_std_logic_vector(52, 8),
51013 => conv_std_logic_vector(53, 8),
51014 => conv_std_logic_vector(54, 8),
51015 => conv_std_logic_vector(55, 8),
51016 => conv_std_logic_vector(55, 8),
51017 => conv_std_logic_vector(56, 8),
51018 => conv_std_logic_vector(57, 8),
51019 => conv_std_logic_vector(58, 8),
51020 => conv_std_logic_vector(59, 8),
51021 => conv_std_logic_vector(59, 8),
51022 => conv_std_logic_vector(60, 8),
51023 => conv_std_logic_vector(61, 8),
51024 => conv_std_logic_vector(62, 8),
51025 => conv_std_logic_vector(62, 8),
51026 => conv_std_logic_vector(63, 8),
51027 => conv_std_logic_vector(64, 8),
51028 => conv_std_logic_vector(65, 8),
51029 => conv_std_logic_vector(66, 8),
51030 => conv_std_logic_vector(66, 8),
51031 => conv_std_logic_vector(67, 8),
51032 => conv_std_logic_vector(68, 8),
51033 => conv_std_logic_vector(69, 8),
51034 => conv_std_logic_vector(69, 8),
51035 => conv_std_logic_vector(70, 8),
51036 => conv_std_logic_vector(71, 8),
51037 => conv_std_logic_vector(72, 8),
51038 => conv_std_logic_vector(73, 8),
51039 => conv_std_logic_vector(73, 8),
51040 => conv_std_logic_vector(74, 8),
51041 => conv_std_logic_vector(75, 8),
51042 => conv_std_logic_vector(76, 8),
51043 => conv_std_logic_vector(76, 8),
51044 => conv_std_logic_vector(77, 8),
51045 => conv_std_logic_vector(78, 8),
51046 => conv_std_logic_vector(79, 8),
51047 => conv_std_logic_vector(80, 8),
51048 => conv_std_logic_vector(80, 8),
51049 => conv_std_logic_vector(81, 8),
51050 => conv_std_logic_vector(82, 8),
51051 => conv_std_logic_vector(83, 8),
51052 => conv_std_logic_vector(83, 8),
51053 => conv_std_logic_vector(84, 8),
51054 => conv_std_logic_vector(85, 8),
51055 => conv_std_logic_vector(86, 8),
51056 => conv_std_logic_vector(87, 8),
51057 => conv_std_logic_vector(87, 8),
51058 => conv_std_logic_vector(88, 8),
51059 => conv_std_logic_vector(89, 8),
51060 => conv_std_logic_vector(90, 8),
51061 => conv_std_logic_vector(90, 8),
51062 => conv_std_logic_vector(91, 8),
51063 => conv_std_logic_vector(92, 8),
51064 => conv_std_logic_vector(93, 8),
51065 => conv_std_logic_vector(94, 8),
51066 => conv_std_logic_vector(94, 8),
51067 => conv_std_logic_vector(95, 8),
51068 => conv_std_logic_vector(96, 8),
51069 => conv_std_logic_vector(97, 8),
51070 => conv_std_logic_vector(97, 8),
51071 => conv_std_logic_vector(98, 8),
51072 => conv_std_logic_vector(99, 8),
51073 => conv_std_logic_vector(100, 8),
51074 => conv_std_logic_vector(101, 8),
51075 => conv_std_logic_vector(101, 8),
51076 => conv_std_logic_vector(102, 8),
51077 => conv_std_logic_vector(103, 8),
51078 => conv_std_logic_vector(104, 8),
51079 => conv_std_logic_vector(104, 8),
51080 => conv_std_logic_vector(105, 8),
51081 => conv_std_logic_vector(106, 8),
51082 => conv_std_logic_vector(107, 8),
51083 => conv_std_logic_vector(108, 8),
51084 => conv_std_logic_vector(108, 8),
51085 => conv_std_logic_vector(109, 8),
51086 => conv_std_logic_vector(110, 8),
51087 => conv_std_logic_vector(111, 8),
51088 => conv_std_logic_vector(111, 8),
51089 => conv_std_logic_vector(112, 8),
51090 => conv_std_logic_vector(113, 8),
51091 => conv_std_logic_vector(114, 8),
51092 => conv_std_logic_vector(115, 8),
51093 => conv_std_logic_vector(115, 8),
51094 => conv_std_logic_vector(116, 8),
51095 => conv_std_logic_vector(117, 8),
51096 => conv_std_logic_vector(118, 8),
51097 => conv_std_logic_vector(118, 8),
51098 => conv_std_logic_vector(119, 8),
51099 => conv_std_logic_vector(120, 8),
51100 => conv_std_logic_vector(121, 8),
51101 => conv_std_logic_vector(122, 8),
51102 => conv_std_logic_vector(122, 8),
51103 => conv_std_logic_vector(123, 8),
51104 => conv_std_logic_vector(124, 8),
51105 => conv_std_logic_vector(125, 8),
51106 => conv_std_logic_vector(125, 8),
51107 => conv_std_logic_vector(126, 8),
51108 => conv_std_logic_vector(127, 8),
51109 => conv_std_logic_vector(128, 8),
51110 => conv_std_logic_vector(129, 8),
51111 => conv_std_logic_vector(129, 8),
51112 => conv_std_logic_vector(130, 8),
51113 => conv_std_logic_vector(131, 8),
51114 => conv_std_logic_vector(132, 8),
51115 => conv_std_logic_vector(132, 8),
51116 => conv_std_logic_vector(133, 8),
51117 => conv_std_logic_vector(134, 8),
51118 => conv_std_logic_vector(135, 8),
51119 => conv_std_logic_vector(136, 8),
51120 => conv_std_logic_vector(136, 8),
51121 => conv_std_logic_vector(137, 8),
51122 => conv_std_logic_vector(138, 8),
51123 => conv_std_logic_vector(139, 8),
51124 => conv_std_logic_vector(139, 8),
51125 => conv_std_logic_vector(140, 8),
51126 => conv_std_logic_vector(141, 8),
51127 => conv_std_logic_vector(142, 8),
51128 => conv_std_logic_vector(143, 8),
51129 => conv_std_logic_vector(143, 8),
51130 => conv_std_logic_vector(144, 8),
51131 => conv_std_logic_vector(145, 8),
51132 => conv_std_logic_vector(146, 8),
51133 => conv_std_logic_vector(146, 8),
51134 => conv_std_logic_vector(147, 8),
51135 => conv_std_logic_vector(148, 8),
51136 => conv_std_logic_vector(149, 8),
51137 => conv_std_logic_vector(150, 8),
51138 => conv_std_logic_vector(150, 8),
51139 => conv_std_logic_vector(151, 8),
51140 => conv_std_logic_vector(152, 8),
51141 => conv_std_logic_vector(153, 8),
51142 => conv_std_logic_vector(153, 8),
51143 => conv_std_logic_vector(154, 8),
51144 => conv_std_logic_vector(155, 8),
51145 => conv_std_logic_vector(156, 8),
51146 => conv_std_logic_vector(157, 8),
51147 => conv_std_logic_vector(157, 8),
51148 => conv_std_logic_vector(158, 8),
51149 => conv_std_logic_vector(159, 8),
51150 => conv_std_logic_vector(160, 8),
51151 => conv_std_logic_vector(160, 8),
51152 => conv_std_logic_vector(161, 8),
51153 => conv_std_logic_vector(162, 8),
51154 => conv_std_logic_vector(163, 8),
51155 => conv_std_logic_vector(164, 8),
51156 => conv_std_logic_vector(164, 8),
51157 => conv_std_logic_vector(165, 8),
51158 => conv_std_logic_vector(166, 8),
51159 => conv_std_logic_vector(167, 8),
51160 => conv_std_logic_vector(167, 8),
51161 => conv_std_logic_vector(168, 8),
51162 => conv_std_logic_vector(169, 8),
51163 => conv_std_logic_vector(170, 8),
51164 => conv_std_logic_vector(171, 8),
51165 => conv_std_logic_vector(171, 8),
51166 => conv_std_logic_vector(172, 8),
51167 => conv_std_logic_vector(173, 8),
51168 => conv_std_logic_vector(174, 8),
51169 => conv_std_logic_vector(174, 8),
51170 => conv_std_logic_vector(175, 8),
51171 => conv_std_logic_vector(176, 8),
51172 => conv_std_logic_vector(177, 8),
51173 => conv_std_logic_vector(178, 8),
51174 => conv_std_logic_vector(178, 8),
51175 => conv_std_logic_vector(179, 8),
51176 => conv_std_logic_vector(180, 8),
51177 => conv_std_logic_vector(181, 8),
51178 => conv_std_logic_vector(181, 8),
51179 => conv_std_logic_vector(182, 8),
51180 => conv_std_logic_vector(183, 8),
51181 => conv_std_logic_vector(184, 8),
51182 => conv_std_logic_vector(185, 8),
51183 => conv_std_logic_vector(185, 8),
51184 => conv_std_logic_vector(186, 8),
51185 => conv_std_logic_vector(187, 8),
51186 => conv_std_logic_vector(188, 8),
51187 => conv_std_logic_vector(188, 8),
51188 => conv_std_logic_vector(189, 8),
51189 => conv_std_logic_vector(190, 8),
51190 => conv_std_logic_vector(191, 8),
51191 => conv_std_logic_vector(192, 8),
51192 => conv_std_logic_vector(192, 8),
51193 => conv_std_logic_vector(193, 8),
51194 => conv_std_logic_vector(194, 8),
51195 => conv_std_logic_vector(195, 8),
51196 => conv_std_logic_vector(195, 8),
51197 => conv_std_logic_vector(196, 8),
51198 => conv_std_logic_vector(197, 8),
51199 => conv_std_logic_vector(198, 8),
51200 => conv_std_logic_vector(0, 8),
51201 => conv_std_logic_vector(0, 8),
51202 => conv_std_logic_vector(1, 8),
51203 => conv_std_logic_vector(2, 8),
51204 => conv_std_logic_vector(3, 8),
51205 => conv_std_logic_vector(3, 8),
51206 => conv_std_logic_vector(4, 8),
51207 => conv_std_logic_vector(5, 8),
51208 => conv_std_logic_vector(6, 8),
51209 => conv_std_logic_vector(7, 8),
51210 => conv_std_logic_vector(7, 8),
51211 => conv_std_logic_vector(8, 8),
51212 => conv_std_logic_vector(9, 8),
51213 => conv_std_logic_vector(10, 8),
51214 => conv_std_logic_vector(10, 8),
51215 => conv_std_logic_vector(11, 8),
51216 => conv_std_logic_vector(12, 8),
51217 => conv_std_logic_vector(13, 8),
51218 => conv_std_logic_vector(14, 8),
51219 => conv_std_logic_vector(14, 8),
51220 => conv_std_logic_vector(15, 8),
51221 => conv_std_logic_vector(16, 8),
51222 => conv_std_logic_vector(17, 8),
51223 => conv_std_logic_vector(17, 8),
51224 => conv_std_logic_vector(18, 8),
51225 => conv_std_logic_vector(19, 8),
51226 => conv_std_logic_vector(20, 8),
51227 => conv_std_logic_vector(21, 8),
51228 => conv_std_logic_vector(21, 8),
51229 => conv_std_logic_vector(22, 8),
51230 => conv_std_logic_vector(23, 8),
51231 => conv_std_logic_vector(24, 8),
51232 => conv_std_logic_vector(25, 8),
51233 => conv_std_logic_vector(25, 8),
51234 => conv_std_logic_vector(26, 8),
51235 => conv_std_logic_vector(27, 8),
51236 => conv_std_logic_vector(28, 8),
51237 => conv_std_logic_vector(28, 8),
51238 => conv_std_logic_vector(29, 8),
51239 => conv_std_logic_vector(30, 8),
51240 => conv_std_logic_vector(31, 8),
51241 => conv_std_logic_vector(32, 8),
51242 => conv_std_logic_vector(32, 8),
51243 => conv_std_logic_vector(33, 8),
51244 => conv_std_logic_vector(34, 8),
51245 => conv_std_logic_vector(35, 8),
51246 => conv_std_logic_vector(35, 8),
51247 => conv_std_logic_vector(36, 8),
51248 => conv_std_logic_vector(37, 8),
51249 => conv_std_logic_vector(38, 8),
51250 => conv_std_logic_vector(39, 8),
51251 => conv_std_logic_vector(39, 8),
51252 => conv_std_logic_vector(40, 8),
51253 => conv_std_logic_vector(41, 8),
51254 => conv_std_logic_vector(42, 8),
51255 => conv_std_logic_vector(42, 8),
51256 => conv_std_logic_vector(43, 8),
51257 => conv_std_logic_vector(44, 8),
51258 => conv_std_logic_vector(45, 8),
51259 => conv_std_logic_vector(46, 8),
51260 => conv_std_logic_vector(46, 8),
51261 => conv_std_logic_vector(47, 8),
51262 => conv_std_logic_vector(48, 8),
51263 => conv_std_logic_vector(49, 8),
51264 => conv_std_logic_vector(50, 8),
51265 => conv_std_logic_vector(50, 8),
51266 => conv_std_logic_vector(51, 8),
51267 => conv_std_logic_vector(52, 8),
51268 => conv_std_logic_vector(53, 8),
51269 => conv_std_logic_vector(53, 8),
51270 => conv_std_logic_vector(54, 8),
51271 => conv_std_logic_vector(55, 8),
51272 => conv_std_logic_vector(56, 8),
51273 => conv_std_logic_vector(57, 8),
51274 => conv_std_logic_vector(57, 8),
51275 => conv_std_logic_vector(58, 8),
51276 => conv_std_logic_vector(59, 8),
51277 => conv_std_logic_vector(60, 8),
51278 => conv_std_logic_vector(60, 8),
51279 => conv_std_logic_vector(61, 8),
51280 => conv_std_logic_vector(62, 8),
51281 => conv_std_logic_vector(63, 8),
51282 => conv_std_logic_vector(64, 8),
51283 => conv_std_logic_vector(64, 8),
51284 => conv_std_logic_vector(65, 8),
51285 => conv_std_logic_vector(66, 8),
51286 => conv_std_logic_vector(67, 8),
51287 => conv_std_logic_vector(67, 8),
51288 => conv_std_logic_vector(68, 8),
51289 => conv_std_logic_vector(69, 8),
51290 => conv_std_logic_vector(70, 8),
51291 => conv_std_logic_vector(71, 8),
51292 => conv_std_logic_vector(71, 8),
51293 => conv_std_logic_vector(72, 8),
51294 => conv_std_logic_vector(73, 8),
51295 => conv_std_logic_vector(74, 8),
51296 => conv_std_logic_vector(75, 8),
51297 => conv_std_logic_vector(75, 8),
51298 => conv_std_logic_vector(76, 8),
51299 => conv_std_logic_vector(77, 8),
51300 => conv_std_logic_vector(78, 8),
51301 => conv_std_logic_vector(78, 8),
51302 => conv_std_logic_vector(79, 8),
51303 => conv_std_logic_vector(80, 8),
51304 => conv_std_logic_vector(81, 8),
51305 => conv_std_logic_vector(82, 8),
51306 => conv_std_logic_vector(82, 8),
51307 => conv_std_logic_vector(83, 8),
51308 => conv_std_logic_vector(84, 8),
51309 => conv_std_logic_vector(85, 8),
51310 => conv_std_logic_vector(85, 8),
51311 => conv_std_logic_vector(86, 8),
51312 => conv_std_logic_vector(87, 8),
51313 => conv_std_logic_vector(88, 8),
51314 => conv_std_logic_vector(89, 8),
51315 => conv_std_logic_vector(89, 8),
51316 => conv_std_logic_vector(90, 8),
51317 => conv_std_logic_vector(91, 8),
51318 => conv_std_logic_vector(92, 8),
51319 => conv_std_logic_vector(92, 8),
51320 => conv_std_logic_vector(93, 8),
51321 => conv_std_logic_vector(94, 8),
51322 => conv_std_logic_vector(95, 8),
51323 => conv_std_logic_vector(96, 8),
51324 => conv_std_logic_vector(96, 8),
51325 => conv_std_logic_vector(97, 8),
51326 => conv_std_logic_vector(98, 8),
51327 => conv_std_logic_vector(99, 8),
51328 => conv_std_logic_vector(100, 8),
51329 => conv_std_logic_vector(100, 8),
51330 => conv_std_logic_vector(101, 8),
51331 => conv_std_logic_vector(102, 8),
51332 => conv_std_logic_vector(103, 8),
51333 => conv_std_logic_vector(103, 8),
51334 => conv_std_logic_vector(104, 8),
51335 => conv_std_logic_vector(105, 8),
51336 => conv_std_logic_vector(106, 8),
51337 => conv_std_logic_vector(107, 8),
51338 => conv_std_logic_vector(107, 8),
51339 => conv_std_logic_vector(108, 8),
51340 => conv_std_logic_vector(109, 8),
51341 => conv_std_logic_vector(110, 8),
51342 => conv_std_logic_vector(110, 8),
51343 => conv_std_logic_vector(111, 8),
51344 => conv_std_logic_vector(112, 8),
51345 => conv_std_logic_vector(113, 8),
51346 => conv_std_logic_vector(114, 8),
51347 => conv_std_logic_vector(114, 8),
51348 => conv_std_logic_vector(115, 8),
51349 => conv_std_logic_vector(116, 8),
51350 => conv_std_logic_vector(117, 8),
51351 => conv_std_logic_vector(117, 8),
51352 => conv_std_logic_vector(118, 8),
51353 => conv_std_logic_vector(119, 8),
51354 => conv_std_logic_vector(120, 8),
51355 => conv_std_logic_vector(121, 8),
51356 => conv_std_logic_vector(121, 8),
51357 => conv_std_logic_vector(122, 8),
51358 => conv_std_logic_vector(123, 8),
51359 => conv_std_logic_vector(124, 8),
51360 => conv_std_logic_vector(125, 8),
51361 => conv_std_logic_vector(125, 8),
51362 => conv_std_logic_vector(126, 8),
51363 => conv_std_logic_vector(127, 8),
51364 => conv_std_logic_vector(128, 8),
51365 => conv_std_logic_vector(128, 8),
51366 => conv_std_logic_vector(129, 8),
51367 => conv_std_logic_vector(130, 8),
51368 => conv_std_logic_vector(131, 8),
51369 => conv_std_logic_vector(132, 8),
51370 => conv_std_logic_vector(132, 8),
51371 => conv_std_logic_vector(133, 8),
51372 => conv_std_logic_vector(134, 8),
51373 => conv_std_logic_vector(135, 8),
51374 => conv_std_logic_vector(135, 8),
51375 => conv_std_logic_vector(136, 8),
51376 => conv_std_logic_vector(137, 8),
51377 => conv_std_logic_vector(138, 8),
51378 => conv_std_logic_vector(139, 8),
51379 => conv_std_logic_vector(139, 8),
51380 => conv_std_logic_vector(140, 8),
51381 => conv_std_logic_vector(141, 8),
51382 => conv_std_logic_vector(142, 8),
51383 => conv_std_logic_vector(142, 8),
51384 => conv_std_logic_vector(143, 8),
51385 => conv_std_logic_vector(144, 8),
51386 => conv_std_logic_vector(145, 8),
51387 => conv_std_logic_vector(146, 8),
51388 => conv_std_logic_vector(146, 8),
51389 => conv_std_logic_vector(147, 8),
51390 => conv_std_logic_vector(148, 8),
51391 => conv_std_logic_vector(149, 8),
51392 => conv_std_logic_vector(150, 8),
51393 => conv_std_logic_vector(150, 8),
51394 => conv_std_logic_vector(151, 8),
51395 => conv_std_logic_vector(152, 8),
51396 => conv_std_logic_vector(153, 8),
51397 => conv_std_logic_vector(153, 8),
51398 => conv_std_logic_vector(154, 8),
51399 => conv_std_logic_vector(155, 8),
51400 => conv_std_logic_vector(156, 8),
51401 => conv_std_logic_vector(157, 8),
51402 => conv_std_logic_vector(157, 8),
51403 => conv_std_logic_vector(158, 8),
51404 => conv_std_logic_vector(159, 8),
51405 => conv_std_logic_vector(160, 8),
51406 => conv_std_logic_vector(160, 8),
51407 => conv_std_logic_vector(161, 8),
51408 => conv_std_logic_vector(162, 8),
51409 => conv_std_logic_vector(163, 8),
51410 => conv_std_logic_vector(164, 8),
51411 => conv_std_logic_vector(164, 8),
51412 => conv_std_logic_vector(165, 8),
51413 => conv_std_logic_vector(166, 8),
51414 => conv_std_logic_vector(167, 8),
51415 => conv_std_logic_vector(167, 8),
51416 => conv_std_logic_vector(168, 8),
51417 => conv_std_logic_vector(169, 8),
51418 => conv_std_logic_vector(170, 8),
51419 => conv_std_logic_vector(171, 8),
51420 => conv_std_logic_vector(171, 8),
51421 => conv_std_logic_vector(172, 8),
51422 => conv_std_logic_vector(173, 8),
51423 => conv_std_logic_vector(174, 8),
51424 => conv_std_logic_vector(175, 8),
51425 => conv_std_logic_vector(175, 8),
51426 => conv_std_logic_vector(176, 8),
51427 => conv_std_logic_vector(177, 8),
51428 => conv_std_logic_vector(178, 8),
51429 => conv_std_logic_vector(178, 8),
51430 => conv_std_logic_vector(179, 8),
51431 => conv_std_logic_vector(180, 8),
51432 => conv_std_logic_vector(181, 8),
51433 => conv_std_logic_vector(182, 8),
51434 => conv_std_logic_vector(182, 8),
51435 => conv_std_logic_vector(183, 8),
51436 => conv_std_logic_vector(184, 8),
51437 => conv_std_logic_vector(185, 8),
51438 => conv_std_logic_vector(185, 8),
51439 => conv_std_logic_vector(186, 8),
51440 => conv_std_logic_vector(187, 8),
51441 => conv_std_logic_vector(188, 8),
51442 => conv_std_logic_vector(189, 8),
51443 => conv_std_logic_vector(189, 8),
51444 => conv_std_logic_vector(190, 8),
51445 => conv_std_logic_vector(191, 8),
51446 => conv_std_logic_vector(192, 8),
51447 => conv_std_logic_vector(192, 8),
51448 => conv_std_logic_vector(193, 8),
51449 => conv_std_logic_vector(194, 8),
51450 => conv_std_logic_vector(195, 8),
51451 => conv_std_logic_vector(196, 8),
51452 => conv_std_logic_vector(196, 8),
51453 => conv_std_logic_vector(197, 8),
51454 => conv_std_logic_vector(198, 8),
51455 => conv_std_logic_vector(199, 8),
51456 => conv_std_logic_vector(0, 8),
51457 => conv_std_logic_vector(0, 8),
51458 => conv_std_logic_vector(1, 8),
51459 => conv_std_logic_vector(2, 8),
51460 => conv_std_logic_vector(3, 8),
51461 => conv_std_logic_vector(3, 8),
51462 => conv_std_logic_vector(4, 8),
51463 => conv_std_logic_vector(5, 8),
51464 => conv_std_logic_vector(6, 8),
51465 => conv_std_logic_vector(7, 8),
51466 => conv_std_logic_vector(7, 8),
51467 => conv_std_logic_vector(8, 8),
51468 => conv_std_logic_vector(9, 8),
51469 => conv_std_logic_vector(10, 8),
51470 => conv_std_logic_vector(10, 8),
51471 => conv_std_logic_vector(11, 8),
51472 => conv_std_logic_vector(12, 8),
51473 => conv_std_logic_vector(13, 8),
51474 => conv_std_logic_vector(14, 8),
51475 => conv_std_logic_vector(14, 8),
51476 => conv_std_logic_vector(15, 8),
51477 => conv_std_logic_vector(16, 8),
51478 => conv_std_logic_vector(17, 8),
51479 => conv_std_logic_vector(18, 8),
51480 => conv_std_logic_vector(18, 8),
51481 => conv_std_logic_vector(19, 8),
51482 => conv_std_logic_vector(20, 8),
51483 => conv_std_logic_vector(21, 8),
51484 => conv_std_logic_vector(21, 8),
51485 => conv_std_logic_vector(22, 8),
51486 => conv_std_logic_vector(23, 8),
51487 => conv_std_logic_vector(24, 8),
51488 => conv_std_logic_vector(25, 8),
51489 => conv_std_logic_vector(25, 8),
51490 => conv_std_logic_vector(26, 8),
51491 => conv_std_logic_vector(27, 8),
51492 => conv_std_logic_vector(28, 8),
51493 => conv_std_logic_vector(29, 8),
51494 => conv_std_logic_vector(29, 8),
51495 => conv_std_logic_vector(30, 8),
51496 => conv_std_logic_vector(31, 8),
51497 => conv_std_logic_vector(32, 8),
51498 => conv_std_logic_vector(32, 8),
51499 => conv_std_logic_vector(33, 8),
51500 => conv_std_logic_vector(34, 8),
51501 => conv_std_logic_vector(35, 8),
51502 => conv_std_logic_vector(36, 8),
51503 => conv_std_logic_vector(36, 8),
51504 => conv_std_logic_vector(37, 8),
51505 => conv_std_logic_vector(38, 8),
51506 => conv_std_logic_vector(39, 8),
51507 => conv_std_logic_vector(40, 8),
51508 => conv_std_logic_vector(40, 8),
51509 => conv_std_logic_vector(41, 8),
51510 => conv_std_logic_vector(42, 8),
51511 => conv_std_logic_vector(43, 8),
51512 => conv_std_logic_vector(43, 8),
51513 => conv_std_logic_vector(44, 8),
51514 => conv_std_logic_vector(45, 8),
51515 => conv_std_logic_vector(46, 8),
51516 => conv_std_logic_vector(47, 8),
51517 => conv_std_logic_vector(47, 8),
51518 => conv_std_logic_vector(48, 8),
51519 => conv_std_logic_vector(49, 8),
51520 => conv_std_logic_vector(50, 8),
51521 => conv_std_logic_vector(51, 8),
51522 => conv_std_logic_vector(51, 8),
51523 => conv_std_logic_vector(52, 8),
51524 => conv_std_logic_vector(53, 8),
51525 => conv_std_logic_vector(54, 8),
51526 => conv_std_logic_vector(54, 8),
51527 => conv_std_logic_vector(55, 8),
51528 => conv_std_logic_vector(56, 8),
51529 => conv_std_logic_vector(57, 8),
51530 => conv_std_logic_vector(58, 8),
51531 => conv_std_logic_vector(58, 8),
51532 => conv_std_logic_vector(59, 8),
51533 => conv_std_logic_vector(60, 8),
51534 => conv_std_logic_vector(61, 8),
51535 => conv_std_logic_vector(62, 8),
51536 => conv_std_logic_vector(62, 8),
51537 => conv_std_logic_vector(63, 8),
51538 => conv_std_logic_vector(64, 8),
51539 => conv_std_logic_vector(65, 8),
51540 => conv_std_logic_vector(65, 8),
51541 => conv_std_logic_vector(66, 8),
51542 => conv_std_logic_vector(67, 8),
51543 => conv_std_logic_vector(68, 8),
51544 => conv_std_logic_vector(69, 8),
51545 => conv_std_logic_vector(69, 8),
51546 => conv_std_logic_vector(70, 8),
51547 => conv_std_logic_vector(71, 8),
51548 => conv_std_logic_vector(72, 8),
51549 => conv_std_logic_vector(73, 8),
51550 => conv_std_logic_vector(73, 8),
51551 => conv_std_logic_vector(74, 8),
51552 => conv_std_logic_vector(75, 8),
51553 => conv_std_logic_vector(76, 8),
51554 => conv_std_logic_vector(76, 8),
51555 => conv_std_logic_vector(77, 8),
51556 => conv_std_logic_vector(78, 8),
51557 => conv_std_logic_vector(79, 8),
51558 => conv_std_logic_vector(80, 8),
51559 => conv_std_logic_vector(80, 8),
51560 => conv_std_logic_vector(81, 8),
51561 => conv_std_logic_vector(82, 8),
51562 => conv_std_logic_vector(83, 8),
51563 => conv_std_logic_vector(84, 8),
51564 => conv_std_logic_vector(84, 8),
51565 => conv_std_logic_vector(85, 8),
51566 => conv_std_logic_vector(86, 8),
51567 => conv_std_logic_vector(87, 8),
51568 => conv_std_logic_vector(87, 8),
51569 => conv_std_logic_vector(88, 8),
51570 => conv_std_logic_vector(89, 8),
51571 => conv_std_logic_vector(90, 8),
51572 => conv_std_logic_vector(91, 8),
51573 => conv_std_logic_vector(91, 8),
51574 => conv_std_logic_vector(92, 8),
51575 => conv_std_logic_vector(93, 8),
51576 => conv_std_logic_vector(94, 8),
51577 => conv_std_logic_vector(95, 8),
51578 => conv_std_logic_vector(95, 8),
51579 => conv_std_logic_vector(96, 8),
51580 => conv_std_logic_vector(97, 8),
51581 => conv_std_logic_vector(98, 8),
51582 => conv_std_logic_vector(98, 8),
51583 => conv_std_logic_vector(99, 8),
51584 => conv_std_logic_vector(100, 8),
51585 => conv_std_logic_vector(101, 8),
51586 => conv_std_logic_vector(102, 8),
51587 => conv_std_logic_vector(102, 8),
51588 => conv_std_logic_vector(103, 8),
51589 => conv_std_logic_vector(104, 8),
51590 => conv_std_logic_vector(105, 8),
51591 => conv_std_logic_vector(105, 8),
51592 => conv_std_logic_vector(106, 8),
51593 => conv_std_logic_vector(107, 8),
51594 => conv_std_logic_vector(108, 8),
51595 => conv_std_logic_vector(109, 8),
51596 => conv_std_logic_vector(109, 8),
51597 => conv_std_logic_vector(110, 8),
51598 => conv_std_logic_vector(111, 8),
51599 => conv_std_logic_vector(112, 8),
51600 => conv_std_logic_vector(113, 8),
51601 => conv_std_logic_vector(113, 8),
51602 => conv_std_logic_vector(114, 8),
51603 => conv_std_logic_vector(115, 8),
51604 => conv_std_logic_vector(116, 8),
51605 => conv_std_logic_vector(116, 8),
51606 => conv_std_logic_vector(117, 8),
51607 => conv_std_logic_vector(118, 8),
51608 => conv_std_logic_vector(119, 8),
51609 => conv_std_logic_vector(120, 8),
51610 => conv_std_logic_vector(120, 8),
51611 => conv_std_logic_vector(121, 8),
51612 => conv_std_logic_vector(122, 8),
51613 => conv_std_logic_vector(123, 8),
51614 => conv_std_logic_vector(124, 8),
51615 => conv_std_logic_vector(124, 8),
51616 => conv_std_logic_vector(125, 8),
51617 => conv_std_logic_vector(126, 8),
51618 => conv_std_logic_vector(127, 8),
51619 => conv_std_logic_vector(127, 8),
51620 => conv_std_logic_vector(128, 8),
51621 => conv_std_logic_vector(129, 8),
51622 => conv_std_logic_vector(130, 8),
51623 => conv_std_logic_vector(131, 8),
51624 => conv_std_logic_vector(131, 8),
51625 => conv_std_logic_vector(132, 8),
51626 => conv_std_logic_vector(133, 8),
51627 => conv_std_logic_vector(134, 8),
51628 => conv_std_logic_vector(135, 8),
51629 => conv_std_logic_vector(135, 8),
51630 => conv_std_logic_vector(136, 8),
51631 => conv_std_logic_vector(137, 8),
51632 => conv_std_logic_vector(138, 8),
51633 => conv_std_logic_vector(138, 8),
51634 => conv_std_logic_vector(139, 8),
51635 => conv_std_logic_vector(140, 8),
51636 => conv_std_logic_vector(141, 8),
51637 => conv_std_logic_vector(142, 8),
51638 => conv_std_logic_vector(142, 8),
51639 => conv_std_logic_vector(143, 8),
51640 => conv_std_logic_vector(144, 8),
51641 => conv_std_logic_vector(145, 8),
51642 => conv_std_logic_vector(146, 8),
51643 => conv_std_logic_vector(146, 8),
51644 => conv_std_logic_vector(147, 8),
51645 => conv_std_logic_vector(148, 8),
51646 => conv_std_logic_vector(149, 8),
51647 => conv_std_logic_vector(149, 8),
51648 => conv_std_logic_vector(150, 8),
51649 => conv_std_logic_vector(151, 8),
51650 => conv_std_logic_vector(152, 8),
51651 => conv_std_logic_vector(153, 8),
51652 => conv_std_logic_vector(153, 8),
51653 => conv_std_logic_vector(154, 8),
51654 => conv_std_logic_vector(155, 8),
51655 => conv_std_logic_vector(156, 8),
51656 => conv_std_logic_vector(157, 8),
51657 => conv_std_logic_vector(157, 8),
51658 => conv_std_logic_vector(158, 8),
51659 => conv_std_logic_vector(159, 8),
51660 => conv_std_logic_vector(160, 8),
51661 => conv_std_logic_vector(160, 8),
51662 => conv_std_logic_vector(161, 8),
51663 => conv_std_logic_vector(162, 8),
51664 => conv_std_logic_vector(163, 8),
51665 => conv_std_logic_vector(164, 8),
51666 => conv_std_logic_vector(164, 8),
51667 => conv_std_logic_vector(165, 8),
51668 => conv_std_logic_vector(166, 8),
51669 => conv_std_logic_vector(167, 8),
51670 => conv_std_logic_vector(168, 8),
51671 => conv_std_logic_vector(168, 8),
51672 => conv_std_logic_vector(169, 8),
51673 => conv_std_logic_vector(170, 8),
51674 => conv_std_logic_vector(171, 8),
51675 => conv_std_logic_vector(171, 8),
51676 => conv_std_logic_vector(172, 8),
51677 => conv_std_logic_vector(173, 8),
51678 => conv_std_logic_vector(174, 8),
51679 => conv_std_logic_vector(175, 8),
51680 => conv_std_logic_vector(175, 8),
51681 => conv_std_logic_vector(176, 8),
51682 => conv_std_logic_vector(177, 8),
51683 => conv_std_logic_vector(178, 8),
51684 => conv_std_logic_vector(179, 8),
51685 => conv_std_logic_vector(179, 8),
51686 => conv_std_logic_vector(180, 8),
51687 => conv_std_logic_vector(181, 8),
51688 => conv_std_logic_vector(182, 8),
51689 => conv_std_logic_vector(182, 8),
51690 => conv_std_logic_vector(183, 8),
51691 => conv_std_logic_vector(184, 8),
51692 => conv_std_logic_vector(185, 8),
51693 => conv_std_logic_vector(186, 8),
51694 => conv_std_logic_vector(186, 8),
51695 => conv_std_logic_vector(187, 8),
51696 => conv_std_logic_vector(188, 8),
51697 => conv_std_logic_vector(189, 8),
51698 => conv_std_logic_vector(190, 8),
51699 => conv_std_logic_vector(190, 8),
51700 => conv_std_logic_vector(191, 8),
51701 => conv_std_logic_vector(192, 8),
51702 => conv_std_logic_vector(193, 8),
51703 => conv_std_logic_vector(193, 8),
51704 => conv_std_logic_vector(194, 8),
51705 => conv_std_logic_vector(195, 8),
51706 => conv_std_logic_vector(196, 8),
51707 => conv_std_logic_vector(197, 8),
51708 => conv_std_logic_vector(197, 8),
51709 => conv_std_logic_vector(198, 8),
51710 => conv_std_logic_vector(199, 8),
51711 => conv_std_logic_vector(200, 8),
51712 => conv_std_logic_vector(0, 8),
51713 => conv_std_logic_vector(0, 8),
51714 => conv_std_logic_vector(1, 8),
51715 => conv_std_logic_vector(2, 8),
51716 => conv_std_logic_vector(3, 8),
51717 => conv_std_logic_vector(3, 8),
51718 => conv_std_logic_vector(4, 8),
51719 => conv_std_logic_vector(5, 8),
51720 => conv_std_logic_vector(6, 8),
51721 => conv_std_logic_vector(7, 8),
51722 => conv_std_logic_vector(7, 8),
51723 => conv_std_logic_vector(8, 8),
51724 => conv_std_logic_vector(9, 8),
51725 => conv_std_logic_vector(10, 8),
51726 => conv_std_logic_vector(11, 8),
51727 => conv_std_logic_vector(11, 8),
51728 => conv_std_logic_vector(12, 8),
51729 => conv_std_logic_vector(13, 8),
51730 => conv_std_logic_vector(14, 8),
51731 => conv_std_logic_vector(14, 8),
51732 => conv_std_logic_vector(15, 8),
51733 => conv_std_logic_vector(16, 8),
51734 => conv_std_logic_vector(17, 8),
51735 => conv_std_logic_vector(18, 8),
51736 => conv_std_logic_vector(18, 8),
51737 => conv_std_logic_vector(19, 8),
51738 => conv_std_logic_vector(20, 8),
51739 => conv_std_logic_vector(21, 8),
51740 => conv_std_logic_vector(22, 8),
51741 => conv_std_logic_vector(22, 8),
51742 => conv_std_logic_vector(23, 8),
51743 => conv_std_logic_vector(24, 8),
51744 => conv_std_logic_vector(25, 8),
51745 => conv_std_logic_vector(26, 8),
51746 => conv_std_logic_vector(26, 8),
51747 => conv_std_logic_vector(27, 8),
51748 => conv_std_logic_vector(28, 8),
51749 => conv_std_logic_vector(29, 8),
51750 => conv_std_logic_vector(29, 8),
51751 => conv_std_logic_vector(30, 8),
51752 => conv_std_logic_vector(31, 8),
51753 => conv_std_logic_vector(32, 8),
51754 => conv_std_logic_vector(33, 8),
51755 => conv_std_logic_vector(33, 8),
51756 => conv_std_logic_vector(34, 8),
51757 => conv_std_logic_vector(35, 8),
51758 => conv_std_logic_vector(36, 8),
51759 => conv_std_logic_vector(37, 8),
51760 => conv_std_logic_vector(37, 8),
51761 => conv_std_logic_vector(38, 8),
51762 => conv_std_logic_vector(39, 8),
51763 => conv_std_logic_vector(40, 8),
51764 => conv_std_logic_vector(41, 8),
51765 => conv_std_logic_vector(41, 8),
51766 => conv_std_logic_vector(42, 8),
51767 => conv_std_logic_vector(43, 8),
51768 => conv_std_logic_vector(44, 8),
51769 => conv_std_logic_vector(44, 8),
51770 => conv_std_logic_vector(45, 8),
51771 => conv_std_logic_vector(46, 8),
51772 => conv_std_logic_vector(47, 8),
51773 => conv_std_logic_vector(48, 8),
51774 => conv_std_logic_vector(48, 8),
51775 => conv_std_logic_vector(49, 8),
51776 => conv_std_logic_vector(50, 8),
51777 => conv_std_logic_vector(51, 8),
51778 => conv_std_logic_vector(52, 8),
51779 => conv_std_logic_vector(52, 8),
51780 => conv_std_logic_vector(53, 8),
51781 => conv_std_logic_vector(54, 8),
51782 => conv_std_logic_vector(55, 8),
51783 => conv_std_logic_vector(56, 8),
51784 => conv_std_logic_vector(56, 8),
51785 => conv_std_logic_vector(57, 8),
51786 => conv_std_logic_vector(58, 8),
51787 => conv_std_logic_vector(59, 8),
51788 => conv_std_logic_vector(59, 8),
51789 => conv_std_logic_vector(60, 8),
51790 => conv_std_logic_vector(61, 8),
51791 => conv_std_logic_vector(62, 8),
51792 => conv_std_logic_vector(63, 8),
51793 => conv_std_logic_vector(63, 8),
51794 => conv_std_logic_vector(64, 8),
51795 => conv_std_logic_vector(65, 8),
51796 => conv_std_logic_vector(66, 8),
51797 => conv_std_logic_vector(67, 8),
51798 => conv_std_logic_vector(67, 8),
51799 => conv_std_logic_vector(68, 8),
51800 => conv_std_logic_vector(69, 8),
51801 => conv_std_logic_vector(70, 8),
51802 => conv_std_logic_vector(71, 8),
51803 => conv_std_logic_vector(71, 8),
51804 => conv_std_logic_vector(72, 8),
51805 => conv_std_logic_vector(73, 8),
51806 => conv_std_logic_vector(74, 8),
51807 => conv_std_logic_vector(74, 8),
51808 => conv_std_logic_vector(75, 8),
51809 => conv_std_logic_vector(76, 8),
51810 => conv_std_logic_vector(77, 8),
51811 => conv_std_logic_vector(78, 8),
51812 => conv_std_logic_vector(78, 8),
51813 => conv_std_logic_vector(79, 8),
51814 => conv_std_logic_vector(80, 8),
51815 => conv_std_logic_vector(81, 8),
51816 => conv_std_logic_vector(82, 8),
51817 => conv_std_logic_vector(82, 8),
51818 => conv_std_logic_vector(83, 8),
51819 => conv_std_logic_vector(84, 8),
51820 => conv_std_logic_vector(85, 8),
51821 => conv_std_logic_vector(86, 8),
51822 => conv_std_logic_vector(86, 8),
51823 => conv_std_logic_vector(87, 8),
51824 => conv_std_logic_vector(88, 8),
51825 => conv_std_logic_vector(89, 8),
51826 => conv_std_logic_vector(89, 8),
51827 => conv_std_logic_vector(90, 8),
51828 => conv_std_logic_vector(91, 8),
51829 => conv_std_logic_vector(92, 8),
51830 => conv_std_logic_vector(93, 8),
51831 => conv_std_logic_vector(93, 8),
51832 => conv_std_logic_vector(94, 8),
51833 => conv_std_logic_vector(95, 8),
51834 => conv_std_logic_vector(96, 8),
51835 => conv_std_logic_vector(97, 8),
51836 => conv_std_logic_vector(97, 8),
51837 => conv_std_logic_vector(98, 8),
51838 => conv_std_logic_vector(99, 8),
51839 => conv_std_logic_vector(100, 8),
51840 => conv_std_logic_vector(101, 8),
51841 => conv_std_logic_vector(101, 8),
51842 => conv_std_logic_vector(102, 8),
51843 => conv_std_logic_vector(103, 8),
51844 => conv_std_logic_vector(104, 8),
51845 => conv_std_logic_vector(104, 8),
51846 => conv_std_logic_vector(105, 8),
51847 => conv_std_logic_vector(106, 8),
51848 => conv_std_logic_vector(107, 8),
51849 => conv_std_logic_vector(108, 8),
51850 => conv_std_logic_vector(108, 8),
51851 => conv_std_logic_vector(109, 8),
51852 => conv_std_logic_vector(110, 8),
51853 => conv_std_logic_vector(111, 8),
51854 => conv_std_logic_vector(112, 8),
51855 => conv_std_logic_vector(112, 8),
51856 => conv_std_logic_vector(113, 8),
51857 => conv_std_logic_vector(114, 8),
51858 => conv_std_logic_vector(115, 8),
51859 => conv_std_logic_vector(115, 8),
51860 => conv_std_logic_vector(116, 8),
51861 => conv_std_logic_vector(117, 8),
51862 => conv_std_logic_vector(118, 8),
51863 => conv_std_logic_vector(119, 8),
51864 => conv_std_logic_vector(119, 8),
51865 => conv_std_logic_vector(120, 8),
51866 => conv_std_logic_vector(121, 8),
51867 => conv_std_logic_vector(122, 8),
51868 => conv_std_logic_vector(123, 8),
51869 => conv_std_logic_vector(123, 8),
51870 => conv_std_logic_vector(124, 8),
51871 => conv_std_logic_vector(125, 8),
51872 => conv_std_logic_vector(126, 8),
51873 => conv_std_logic_vector(127, 8),
51874 => conv_std_logic_vector(127, 8),
51875 => conv_std_logic_vector(128, 8),
51876 => conv_std_logic_vector(129, 8),
51877 => conv_std_logic_vector(130, 8),
51878 => conv_std_logic_vector(130, 8),
51879 => conv_std_logic_vector(131, 8),
51880 => conv_std_logic_vector(132, 8),
51881 => conv_std_logic_vector(133, 8),
51882 => conv_std_logic_vector(134, 8),
51883 => conv_std_logic_vector(134, 8),
51884 => conv_std_logic_vector(135, 8),
51885 => conv_std_logic_vector(136, 8),
51886 => conv_std_logic_vector(137, 8),
51887 => conv_std_logic_vector(138, 8),
51888 => conv_std_logic_vector(138, 8),
51889 => conv_std_logic_vector(139, 8),
51890 => conv_std_logic_vector(140, 8),
51891 => conv_std_logic_vector(141, 8),
51892 => conv_std_logic_vector(142, 8),
51893 => conv_std_logic_vector(142, 8),
51894 => conv_std_logic_vector(143, 8),
51895 => conv_std_logic_vector(144, 8),
51896 => conv_std_logic_vector(145, 8),
51897 => conv_std_logic_vector(145, 8),
51898 => conv_std_logic_vector(146, 8),
51899 => conv_std_logic_vector(147, 8),
51900 => conv_std_logic_vector(148, 8),
51901 => conv_std_logic_vector(149, 8),
51902 => conv_std_logic_vector(149, 8),
51903 => conv_std_logic_vector(150, 8),
51904 => conv_std_logic_vector(151, 8),
51905 => conv_std_logic_vector(152, 8),
51906 => conv_std_logic_vector(153, 8),
51907 => conv_std_logic_vector(153, 8),
51908 => conv_std_logic_vector(154, 8),
51909 => conv_std_logic_vector(155, 8),
51910 => conv_std_logic_vector(156, 8),
51911 => conv_std_logic_vector(157, 8),
51912 => conv_std_logic_vector(157, 8),
51913 => conv_std_logic_vector(158, 8),
51914 => conv_std_logic_vector(159, 8),
51915 => conv_std_logic_vector(160, 8),
51916 => conv_std_logic_vector(160, 8),
51917 => conv_std_logic_vector(161, 8),
51918 => conv_std_logic_vector(162, 8),
51919 => conv_std_logic_vector(163, 8),
51920 => conv_std_logic_vector(164, 8),
51921 => conv_std_logic_vector(164, 8),
51922 => conv_std_logic_vector(165, 8),
51923 => conv_std_logic_vector(166, 8),
51924 => conv_std_logic_vector(167, 8),
51925 => conv_std_logic_vector(168, 8),
51926 => conv_std_logic_vector(168, 8),
51927 => conv_std_logic_vector(169, 8),
51928 => conv_std_logic_vector(170, 8),
51929 => conv_std_logic_vector(171, 8),
51930 => conv_std_logic_vector(172, 8),
51931 => conv_std_logic_vector(172, 8),
51932 => conv_std_logic_vector(173, 8),
51933 => conv_std_logic_vector(174, 8),
51934 => conv_std_logic_vector(175, 8),
51935 => conv_std_logic_vector(175, 8),
51936 => conv_std_logic_vector(176, 8),
51937 => conv_std_logic_vector(177, 8),
51938 => conv_std_logic_vector(178, 8),
51939 => conv_std_logic_vector(179, 8),
51940 => conv_std_logic_vector(179, 8),
51941 => conv_std_logic_vector(180, 8),
51942 => conv_std_logic_vector(181, 8),
51943 => conv_std_logic_vector(182, 8),
51944 => conv_std_logic_vector(183, 8),
51945 => conv_std_logic_vector(183, 8),
51946 => conv_std_logic_vector(184, 8),
51947 => conv_std_logic_vector(185, 8),
51948 => conv_std_logic_vector(186, 8),
51949 => conv_std_logic_vector(187, 8),
51950 => conv_std_logic_vector(187, 8),
51951 => conv_std_logic_vector(188, 8),
51952 => conv_std_logic_vector(189, 8),
51953 => conv_std_logic_vector(190, 8),
51954 => conv_std_logic_vector(190, 8),
51955 => conv_std_logic_vector(191, 8),
51956 => conv_std_logic_vector(192, 8),
51957 => conv_std_logic_vector(193, 8),
51958 => conv_std_logic_vector(194, 8),
51959 => conv_std_logic_vector(194, 8),
51960 => conv_std_logic_vector(195, 8),
51961 => conv_std_logic_vector(196, 8),
51962 => conv_std_logic_vector(197, 8),
51963 => conv_std_logic_vector(198, 8),
51964 => conv_std_logic_vector(198, 8),
51965 => conv_std_logic_vector(199, 8),
51966 => conv_std_logic_vector(200, 8),
51967 => conv_std_logic_vector(201, 8),
51968 => conv_std_logic_vector(0, 8),
51969 => conv_std_logic_vector(0, 8),
51970 => conv_std_logic_vector(1, 8),
51971 => conv_std_logic_vector(2, 8),
51972 => conv_std_logic_vector(3, 8),
51973 => conv_std_logic_vector(3, 8),
51974 => conv_std_logic_vector(4, 8),
51975 => conv_std_logic_vector(5, 8),
51976 => conv_std_logic_vector(6, 8),
51977 => conv_std_logic_vector(7, 8),
51978 => conv_std_logic_vector(7, 8),
51979 => conv_std_logic_vector(8, 8),
51980 => conv_std_logic_vector(9, 8),
51981 => conv_std_logic_vector(10, 8),
51982 => conv_std_logic_vector(11, 8),
51983 => conv_std_logic_vector(11, 8),
51984 => conv_std_logic_vector(12, 8),
51985 => conv_std_logic_vector(13, 8),
51986 => conv_std_logic_vector(14, 8),
51987 => conv_std_logic_vector(15, 8),
51988 => conv_std_logic_vector(15, 8),
51989 => conv_std_logic_vector(16, 8),
51990 => conv_std_logic_vector(17, 8),
51991 => conv_std_logic_vector(18, 8),
51992 => conv_std_logic_vector(19, 8),
51993 => conv_std_logic_vector(19, 8),
51994 => conv_std_logic_vector(20, 8),
51995 => conv_std_logic_vector(21, 8),
51996 => conv_std_logic_vector(22, 8),
51997 => conv_std_logic_vector(22, 8),
51998 => conv_std_logic_vector(23, 8),
51999 => conv_std_logic_vector(24, 8),
52000 => conv_std_logic_vector(25, 8),
52001 => conv_std_logic_vector(26, 8),
52002 => conv_std_logic_vector(26, 8),
52003 => conv_std_logic_vector(27, 8),
52004 => conv_std_logic_vector(28, 8),
52005 => conv_std_logic_vector(29, 8),
52006 => conv_std_logic_vector(30, 8),
52007 => conv_std_logic_vector(30, 8),
52008 => conv_std_logic_vector(31, 8),
52009 => conv_std_logic_vector(32, 8),
52010 => conv_std_logic_vector(33, 8),
52011 => conv_std_logic_vector(34, 8),
52012 => conv_std_logic_vector(34, 8),
52013 => conv_std_logic_vector(35, 8),
52014 => conv_std_logic_vector(36, 8),
52015 => conv_std_logic_vector(37, 8),
52016 => conv_std_logic_vector(38, 8),
52017 => conv_std_logic_vector(38, 8),
52018 => conv_std_logic_vector(39, 8),
52019 => conv_std_logic_vector(40, 8),
52020 => conv_std_logic_vector(41, 8),
52021 => conv_std_logic_vector(42, 8),
52022 => conv_std_logic_vector(42, 8),
52023 => conv_std_logic_vector(43, 8),
52024 => conv_std_logic_vector(44, 8),
52025 => conv_std_logic_vector(45, 8),
52026 => conv_std_logic_vector(45, 8),
52027 => conv_std_logic_vector(46, 8),
52028 => conv_std_logic_vector(47, 8),
52029 => conv_std_logic_vector(48, 8),
52030 => conv_std_logic_vector(49, 8),
52031 => conv_std_logic_vector(49, 8),
52032 => conv_std_logic_vector(50, 8),
52033 => conv_std_logic_vector(51, 8),
52034 => conv_std_logic_vector(52, 8),
52035 => conv_std_logic_vector(53, 8),
52036 => conv_std_logic_vector(53, 8),
52037 => conv_std_logic_vector(54, 8),
52038 => conv_std_logic_vector(55, 8),
52039 => conv_std_logic_vector(56, 8),
52040 => conv_std_logic_vector(57, 8),
52041 => conv_std_logic_vector(57, 8),
52042 => conv_std_logic_vector(58, 8),
52043 => conv_std_logic_vector(59, 8),
52044 => conv_std_logic_vector(60, 8),
52045 => conv_std_logic_vector(61, 8),
52046 => conv_std_logic_vector(61, 8),
52047 => conv_std_logic_vector(62, 8),
52048 => conv_std_logic_vector(63, 8),
52049 => conv_std_logic_vector(64, 8),
52050 => conv_std_logic_vector(65, 8),
52051 => conv_std_logic_vector(65, 8),
52052 => conv_std_logic_vector(66, 8),
52053 => conv_std_logic_vector(67, 8),
52054 => conv_std_logic_vector(68, 8),
52055 => conv_std_logic_vector(68, 8),
52056 => conv_std_logic_vector(69, 8),
52057 => conv_std_logic_vector(70, 8),
52058 => conv_std_logic_vector(71, 8),
52059 => conv_std_logic_vector(72, 8),
52060 => conv_std_logic_vector(72, 8),
52061 => conv_std_logic_vector(73, 8),
52062 => conv_std_logic_vector(74, 8),
52063 => conv_std_logic_vector(75, 8),
52064 => conv_std_logic_vector(76, 8),
52065 => conv_std_logic_vector(76, 8),
52066 => conv_std_logic_vector(77, 8),
52067 => conv_std_logic_vector(78, 8),
52068 => conv_std_logic_vector(79, 8),
52069 => conv_std_logic_vector(80, 8),
52070 => conv_std_logic_vector(80, 8),
52071 => conv_std_logic_vector(81, 8),
52072 => conv_std_logic_vector(82, 8),
52073 => conv_std_logic_vector(83, 8),
52074 => conv_std_logic_vector(84, 8),
52075 => conv_std_logic_vector(84, 8),
52076 => conv_std_logic_vector(85, 8),
52077 => conv_std_logic_vector(86, 8),
52078 => conv_std_logic_vector(87, 8),
52079 => conv_std_logic_vector(88, 8),
52080 => conv_std_logic_vector(88, 8),
52081 => conv_std_logic_vector(89, 8),
52082 => conv_std_logic_vector(90, 8),
52083 => conv_std_logic_vector(91, 8),
52084 => conv_std_logic_vector(91, 8),
52085 => conv_std_logic_vector(92, 8),
52086 => conv_std_logic_vector(93, 8),
52087 => conv_std_logic_vector(94, 8),
52088 => conv_std_logic_vector(95, 8),
52089 => conv_std_logic_vector(95, 8),
52090 => conv_std_logic_vector(96, 8),
52091 => conv_std_logic_vector(97, 8),
52092 => conv_std_logic_vector(98, 8),
52093 => conv_std_logic_vector(99, 8),
52094 => conv_std_logic_vector(99, 8),
52095 => conv_std_logic_vector(100, 8),
52096 => conv_std_logic_vector(101, 8),
52097 => conv_std_logic_vector(102, 8),
52098 => conv_std_logic_vector(103, 8),
52099 => conv_std_logic_vector(103, 8),
52100 => conv_std_logic_vector(104, 8),
52101 => conv_std_logic_vector(105, 8),
52102 => conv_std_logic_vector(106, 8),
52103 => conv_std_logic_vector(107, 8),
52104 => conv_std_logic_vector(107, 8),
52105 => conv_std_logic_vector(108, 8),
52106 => conv_std_logic_vector(109, 8),
52107 => conv_std_logic_vector(110, 8),
52108 => conv_std_logic_vector(111, 8),
52109 => conv_std_logic_vector(111, 8),
52110 => conv_std_logic_vector(112, 8),
52111 => conv_std_logic_vector(113, 8),
52112 => conv_std_logic_vector(114, 8),
52113 => conv_std_logic_vector(114, 8),
52114 => conv_std_logic_vector(115, 8),
52115 => conv_std_logic_vector(116, 8),
52116 => conv_std_logic_vector(117, 8),
52117 => conv_std_logic_vector(118, 8),
52118 => conv_std_logic_vector(118, 8),
52119 => conv_std_logic_vector(119, 8),
52120 => conv_std_logic_vector(120, 8),
52121 => conv_std_logic_vector(121, 8),
52122 => conv_std_logic_vector(122, 8),
52123 => conv_std_logic_vector(122, 8),
52124 => conv_std_logic_vector(123, 8),
52125 => conv_std_logic_vector(124, 8),
52126 => conv_std_logic_vector(125, 8),
52127 => conv_std_logic_vector(126, 8),
52128 => conv_std_logic_vector(126, 8),
52129 => conv_std_logic_vector(127, 8),
52130 => conv_std_logic_vector(128, 8),
52131 => conv_std_logic_vector(129, 8),
52132 => conv_std_logic_vector(130, 8),
52133 => conv_std_logic_vector(130, 8),
52134 => conv_std_logic_vector(131, 8),
52135 => conv_std_logic_vector(132, 8),
52136 => conv_std_logic_vector(133, 8),
52137 => conv_std_logic_vector(134, 8),
52138 => conv_std_logic_vector(134, 8),
52139 => conv_std_logic_vector(135, 8),
52140 => conv_std_logic_vector(136, 8),
52141 => conv_std_logic_vector(137, 8),
52142 => conv_std_logic_vector(137, 8),
52143 => conv_std_logic_vector(138, 8),
52144 => conv_std_logic_vector(139, 8),
52145 => conv_std_logic_vector(140, 8),
52146 => conv_std_logic_vector(141, 8),
52147 => conv_std_logic_vector(141, 8),
52148 => conv_std_logic_vector(142, 8),
52149 => conv_std_logic_vector(143, 8),
52150 => conv_std_logic_vector(144, 8),
52151 => conv_std_logic_vector(145, 8),
52152 => conv_std_logic_vector(145, 8),
52153 => conv_std_logic_vector(146, 8),
52154 => conv_std_logic_vector(147, 8),
52155 => conv_std_logic_vector(148, 8),
52156 => conv_std_logic_vector(149, 8),
52157 => conv_std_logic_vector(149, 8),
52158 => conv_std_logic_vector(150, 8),
52159 => conv_std_logic_vector(151, 8),
52160 => conv_std_logic_vector(152, 8),
52161 => conv_std_logic_vector(153, 8),
52162 => conv_std_logic_vector(153, 8),
52163 => conv_std_logic_vector(154, 8),
52164 => conv_std_logic_vector(155, 8),
52165 => conv_std_logic_vector(156, 8),
52166 => conv_std_logic_vector(157, 8),
52167 => conv_std_logic_vector(157, 8),
52168 => conv_std_logic_vector(158, 8),
52169 => conv_std_logic_vector(159, 8),
52170 => conv_std_logic_vector(160, 8),
52171 => conv_std_logic_vector(160, 8),
52172 => conv_std_logic_vector(161, 8),
52173 => conv_std_logic_vector(162, 8),
52174 => conv_std_logic_vector(163, 8),
52175 => conv_std_logic_vector(164, 8),
52176 => conv_std_logic_vector(164, 8),
52177 => conv_std_logic_vector(165, 8),
52178 => conv_std_logic_vector(166, 8),
52179 => conv_std_logic_vector(167, 8),
52180 => conv_std_logic_vector(168, 8),
52181 => conv_std_logic_vector(168, 8),
52182 => conv_std_logic_vector(169, 8),
52183 => conv_std_logic_vector(170, 8),
52184 => conv_std_logic_vector(171, 8),
52185 => conv_std_logic_vector(172, 8),
52186 => conv_std_logic_vector(172, 8),
52187 => conv_std_logic_vector(173, 8),
52188 => conv_std_logic_vector(174, 8),
52189 => conv_std_logic_vector(175, 8),
52190 => conv_std_logic_vector(176, 8),
52191 => conv_std_logic_vector(176, 8),
52192 => conv_std_logic_vector(177, 8),
52193 => conv_std_logic_vector(178, 8),
52194 => conv_std_logic_vector(179, 8),
52195 => conv_std_logic_vector(180, 8),
52196 => conv_std_logic_vector(180, 8),
52197 => conv_std_logic_vector(181, 8),
52198 => conv_std_logic_vector(182, 8),
52199 => conv_std_logic_vector(183, 8),
52200 => conv_std_logic_vector(183, 8),
52201 => conv_std_logic_vector(184, 8),
52202 => conv_std_logic_vector(185, 8),
52203 => conv_std_logic_vector(186, 8),
52204 => conv_std_logic_vector(187, 8),
52205 => conv_std_logic_vector(187, 8),
52206 => conv_std_logic_vector(188, 8),
52207 => conv_std_logic_vector(189, 8),
52208 => conv_std_logic_vector(190, 8),
52209 => conv_std_logic_vector(191, 8),
52210 => conv_std_logic_vector(191, 8),
52211 => conv_std_logic_vector(192, 8),
52212 => conv_std_logic_vector(193, 8),
52213 => conv_std_logic_vector(194, 8),
52214 => conv_std_logic_vector(195, 8),
52215 => conv_std_logic_vector(195, 8),
52216 => conv_std_logic_vector(196, 8),
52217 => conv_std_logic_vector(197, 8),
52218 => conv_std_logic_vector(198, 8),
52219 => conv_std_logic_vector(199, 8),
52220 => conv_std_logic_vector(199, 8),
52221 => conv_std_logic_vector(200, 8),
52222 => conv_std_logic_vector(201, 8),
52223 => conv_std_logic_vector(202, 8),
52224 => conv_std_logic_vector(0, 8),
52225 => conv_std_logic_vector(0, 8),
52226 => conv_std_logic_vector(1, 8),
52227 => conv_std_logic_vector(2, 8),
52228 => conv_std_logic_vector(3, 8),
52229 => conv_std_logic_vector(3, 8),
52230 => conv_std_logic_vector(4, 8),
52231 => conv_std_logic_vector(5, 8),
52232 => conv_std_logic_vector(6, 8),
52233 => conv_std_logic_vector(7, 8),
52234 => conv_std_logic_vector(7, 8),
52235 => conv_std_logic_vector(8, 8),
52236 => conv_std_logic_vector(9, 8),
52237 => conv_std_logic_vector(10, 8),
52238 => conv_std_logic_vector(11, 8),
52239 => conv_std_logic_vector(11, 8),
52240 => conv_std_logic_vector(12, 8),
52241 => conv_std_logic_vector(13, 8),
52242 => conv_std_logic_vector(14, 8),
52243 => conv_std_logic_vector(15, 8),
52244 => conv_std_logic_vector(15, 8),
52245 => conv_std_logic_vector(16, 8),
52246 => conv_std_logic_vector(17, 8),
52247 => conv_std_logic_vector(18, 8),
52248 => conv_std_logic_vector(19, 8),
52249 => conv_std_logic_vector(19, 8),
52250 => conv_std_logic_vector(20, 8),
52251 => conv_std_logic_vector(21, 8),
52252 => conv_std_logic_vector(22, 8),
52253 => conv_std_logic_vector(23, 8),
52254 => conv_std_logic_vector(23, 8),
52255 => conv_std_logic_vector(24, 8),
52256 => conv_std_logic_vector(25, 8),
52257 => conv_std_logic_vector(26, 8),
52258 => conv_std_logic_vector(27, 8),
52259 => conv_std_logic_vector(27, 8),
52260 => conv_std_logic_vector(28, 8),
52261 => conv_std_logic_vector(29, 8),
52262 => conv_std_logic_vector(30, 8),
52263 => conv_std_logic_vector(31, 8),
52264 => conv_std_logic_vector(31, 8),
52265 => conv_std_logic_vector(32, 8),
52266 => conv_std_logic_vector(33, 8),
52267 => conv_std_logic_vector(34, 8),
52268 => conv_std_logic_vector(35, 8),
52269 => conv_std_logic_vector(35, 8),
52270 => conv_std_logic_vector(36, 8),
52271 => conv_std_logic_vector(37, 8),
52272 => conv_std_logic_vector(38, 8),
52273 => conv_std_logic_vector(39, 8),
52274 => conv_std_logic_vector(39, 8),
52275 => conv_std_logic_vector(40, 8),
52276 => conv_std_logic_vector(41, 8),
52277 => conv_std_logic_vector(42, 8),
52278 => conv_std_logic_vector(43, 8),
52279 => conv_std_logic_vector(43, 8),
52280 => conv_std_logic_vector(44, 8),
52281 => conv_std_logic_vector(45, 8),
52282 => conv_std_logic_vector(46, 8),
52283 => conv_std_logic_vector(47, 8),
52284 => conv_std_logic_vector(47, 8),
52285 => conv_std_logic_vector(48, 8),
52286 => conv_std_logic_vector(49, 8),
52287 => conv_std_logic_vector(50, 8),
52288 => conv_std_logic_vector(51, 8),
52289 => conv_std_logic_vector(51, 8),
52290 => conv_std_logic_vector(52, 8),
52291 => conv_std_logic_vector(53, 8),
52292 => conv_std_logic_vector(54, 8),
52293 => conv_std_logic_vector(54, 8),
52294 => conv_std_logic_vector(55, 8),
52295 => conv_std_logic_vector(56, 8),
52296 => conv_std_logic_vector(57, 8),
52297 => conv_std_logic_vector(58, 8),
52298 => conv_std_logic_vector(58, 8),
52299 => conv_std_logic_vector(59, 8),
52300 => conv_std_logic_vector(60, 8),
52301 => conv_std_logic_vector(61, 8),
52302 => conv_std_logic_vector(62, 8),
52303 => conv_std_logic_vector(62, 8),
52304 => conv_std_logic_vector(63, 8),
52305 => conv_std_logic_vector(64, 8),
52306 => conv_std_logic_vector(65, 8),
52307 => conv_std_logic_vector(66, 8),
52308 => conv_std_logic_vector(66, 8),
52309 => conv_std_logic_vector(67, 8),
52310 => conv_std_logic_vector(68, 8),
52311 => conv_std_logic_vector(69, 8),
52312 => conv_std_logic_vector(70, 8),
52313 => conv_std_logic_vector(70, 8),
52314 => conv_std_logic_vector(71, 8),
52315 => conv_std_logic_vector(72, 8),
52316 => conv_std_logic_vector(73, 8),
52317 => conv_std_logic_vector(74, 8),
52318 => conv_std_logic_vector(74, 8),
52319 => conv_std_logic_vector(75, 8),
52320 => conv_std_logic_vector(76, 8),
52321 => conv_std_logic_vector(77, 8),
52322 => conv_std_logic_vector(78, 8),
52323 => conv_std_logic_vector(78, 8),
52324 => conv_std_logic_vector(79, 8),
52325 => conv_std_logic_vector(80, 8),
52326 => conv_std_logic_vector(81, 8),
52327 => conv_std_logic_vector(82, 8),
52328 => conv_std_logic_vector(82, 8),
52329 => conv_std_logic_vector(83, 8),
52330 => conv_std_logic_vector(84, 8),
52331 => conv_std_logic_vector(85, 8),
52332 => conv_std_logic_vector(86, 8),
52333 => conv_std_logic_vector(86, 8),
52334 => conv_std_logic_vector(87, 8),
52335 => conv_std_logic_vector(88, 8),
52336 => conv_std_logic_vector(89, 8),
52337 => conv_std_logic_vector(90, 8),
52338 => conv_std_logic_vector(90, 8),
52339 => conv_std_logic_vector(91, 8),
52340 => conv_std_logic_vector(92, 8),
52341 => conv_std_logic_vector(93, 8),
52342 => conv_std_logic_vector(94, 8),
52343 => conv_std_logic_vector(94, 8),
52344 => conv_std_logic_vector(95, 8),
52345 => conv_std_logic_vector(96, 8),
52346 => conv_std_logic_vector(97, 8),
52347 => conv_std_logic_vector(98, 8),
52348 => conv_std_logic_vector(98, 8),
52349 => conv_std_logic_vector(99, 8),
52350 => conv_std_logic_vector(100, 8),
52351 => conv_std_logic_vector(101, 8),
52352 => conv_std_logic_vector(102, 8),
52353 => conv_std_logic_vector(102, 8),
52354 => conv_std_logic_vector(103, 8),
52355 => conv_std_logic_vector(104, 8),
52356 => conv_std_logic_vector(105, 8),
52357 => conv_std_logic_vector(105, 8),
52358 => conv_std_logic_vector(106, 8),
52359 => conv_std_logic_vector(107, 8),
52360 => conv_std_logic_vector(108, 8),
52361 => conv_std_logic_vector(109, 8),
52362 => conv_std_logic_vector(109, 8),
52363 => conv_std_logic_vector(110, 8),
52364 => conv_std_logic_vector(111, 8),
52365 => conv_std_logic_vector(112, 8),
52366 => conv_std_logic_vector(113, 8),
52367 => conv_std_logic_vector(113, 8),
52368 => conv_std_logic_vector(114, 8),
52369 => conv_std_logic_vector(115, 8),
52370 => conv_std_logic_vector(116, 8),
52371 => conv_std_logic_vector(117, 8),
52372 => conv_std_logic_vector(117, 8),
52373 => conv_std_logic_vector(118, 8),
52374 => conv_std_logic_vector(119, 8),
52375 => conv_std_logic_vector(120, 8),
52376 => conv_std_logic_vector(121, 8),
52377 => conv_std_logic_vector(121, 8),
52378 => conv_std_logic_vector(122, 8),
52379 => conv_std_logic_vector(123, 8),
52380 => conv_std_logic_vector(124, 8),
52381 => conv_std_logic_vector(125, 8),
52382 => conv_std_logic_vector(125, 8),
52383 => conv_std_logic_vector(126, 8),
52384 => conv_std_logic_vector(127, 8),
52385 => conv_std_logic_vector(128, 8),
52386 => conv_std_logic_vector(129, 8),
52387 => conv_std_logic_vector(129, 8),
52388 => conv_std_logic_vector(130, 8),
52389 => conv_std_logic_vector(131, 8),
52390 => conv_std_logic_vector(132, 8),
52391 => conv_std_logic_vector(133, 8),
52392 => conv_std_logic_vector(133, 8),
52393 => conv_std_logic_vector(134, 8),
52394 => conv_std_logic_vector(135, 8),
52395 => conv_std_logic_vector(136, 8),
52396 => conv_std_logic_vector(137, 8),
52397 => conv_std_logic_vector(137, 8),
52398 => conv_std_logic_vector(138, 8),
52399 => conv_std_logic_vector(139, 8),
52400 => conv_std_logic_vector(140, 8),
52401 => conv_std_logic_vector(141, 8),
52402 => conv_std_logic_vector(141, 8),
52403 => conv_std_logic_vector(142, 8),
52404 => conv_std_logic_vector(143, 8),
52405 => conv_std_logic_vector(144, 8),
52406 => conv_std_logic_vector(145, 8),
52407 => conv_std_logic_vector(145, 8),
52408 => conv_std_logic_vector(146, 8),
52409 => conv_std_logic_vector(147, 8),
52410 => conv_std_logic_vector(148, 8),
52411 => conv_std_logic_vector(149, 8),
52412 => conv_std_logic_vector(149, 8),
52413 => conv_std_logic_vector(150, 8),
52414 => conv_std_logic_vector(151, 8),
52415 => conv_std_logic_vector(152, 8),
52416 => conv_std_logic_vector(153, 8),
52417 => conv_std_logic_vector(153, 8),
52418 => conv_std_logic_vector(154, 8),
52419 => conv_std_logic_vector(155, 8),
52420 => conv_std_logic_vector(156, 8),
52421 => conv_std_logic_vector(156, 8),
52422 => conv_std_logic_vector(157, 8),
52423 => conv_std_logic_vector(158, 8),
52424 => conv_std_logic_vector(159, 8),
52425 => conv_std_logic_vector(160, 8),
52426 => conv_std_logic_vector(160, 8),
52427 => conv_std_logic_vector(161, 8),
52428 => conv_std_logic_vector(162, 8),
52429 => conv_std_logic_vector(163, 8),
52430 => conv_std_logic_vector(164, 8),
52431 => conv_std_logic_vector(164, 8),
52432 => conv_std_logic_vector(165, 8),
52433 => conv_std_logic_vector(166, 8),
52434 => conv_std_logic_vector(167, 8),
52435 => conv_std_logic_vector(168, 8),
52436 => conv_std_logic_vector(168, 8),
52437 => conv_std_logic_vector(169, 8),
52438 => conv_std_logic_vector(170, 8),
52439 => conv_std_logic_vector(171, 8),
52440 => conv_std_logic_vector(172, 8),
52441 => conv_std_logic_vector(172, 8),
52442 => conv_std_logic_vector(173, 8),
52443 => conv_std_logic_vector(174, 8),
52444 => conv_std_logic_vector(175, 8),
52445 => conv_std_logic_vector(176, 8),
52446 => conv_std_logic_vector(176, 8),
52447 => conv_std_logic_vector(177, 8),
52448 => conv_std_logic_vector(178, 8),
52449 => conv_std_logic_vector(179, 8),
52450 => conv_std_logic_vector(180, 8),
52451 => conv_std_logic_vector(180, 8),
52452 => conv_std_logic_vector(181, 8),
52453 => conv_std_logic_vector(182, 8),
52454 => conv_std_logic_vector(183, 8),
52455 => conv_std_logic_vector(184, 8),
52456 => conv_std_logic_vector(184, 8),
52457 => conv_std_logic_vector(185, 8),
52458 => conv_std_logic_vector(186, 8),
52459 => conv_std_logic_vector(187, 8),
52460 => conv_std_logic_vector(188, 8),
52461 => conv_std_logic_vector(188, 8),
52462 => conv_std_logic_vector(189, 8),
52463 => conv_std_logic_vector(190, 8),
52464 => conv_std_logic_vector(191, 8),
52465 => conv_std_logic_vector(192, 8),
52466 => conv_std_logic_vector(192, 8),
52467 => conv_std_logic_vector(193, 8),
52468 => conv_std_logic_vector(194, 8),
52469 => conv_std_logic_vector(195, 8),
52470 => conv_std_logic_vector(196, 8),
52471 => conv_std_logic_vector(196, 8),
52472 => conv_std_logic_vector(197, 8),
52473 => conv_std_logic_vector(198, 8),
52474 => conv_std_logic_vector(199, 8),
52475 => conv_std_logic_vector(200, 8),
52476 => conv_std_logic_vector(200, 8),
52477 => conv_std_logic_vector(201, 8),
52478 => conv_std_logic_vector(202, 8),
52479 => conv_std_logic_vector(203, 8),
52480 => conv_std_logic_vector(0, 8),
52481 => conv_std_logic_vector(0, 8),
52482 => conv_std_logic_vector(1, 8),
52483 => conv_std_logic_vector(2, 8),
52484 => conv_std_logic_vector(3, 8),
52485 => conv_std_logic_vector(4, 8),
52486 => conv_std_logic_vector(4, 8),
52487 => conv_std_logic_vector(5, 8),
52488 => conv_std_logic_vector(6, 8),
52489 => conv_std_logic_vector(7, 8),
52490 => conv_std_logic_vector(8, 8),
52491 => conv_std_logic_vector(8, 8),
52492 => conv_std_logic_vector(9, 8),
52493 => conv_std_logic_vector(10, 8),
52494 => conv_std_logic_vector(11, 8),
52495 => conv_std_logic_vector(12, 8),
52496 => conv_std_logic_vector(12, 8),
52497 => conv_std_logic_vector(13, 8),
52498 => conv_std_logic_vector(14, 8),
52499 => conv_std_logic_vector(15, 8),
52500 => conv_std_logic_vector(16, 8),
52501 => conv_std_logic_vector(16, 8),
52502 => conv_std_logic_vector(17, 8),
52503 => conv_std_logic_vector(18, 8),
52504 => conv_std_logic_vector(19, 8),
52505 => conv_std_logic_vector(20, 8),
52506 => conv_std_logic_vector(20, 8),
52507 => conv_std_logic_vector(21, 8),
52508 => conv_std_logic_vector(22, 8),
52509 => conv_std_logic_vector(23, 8),
52510 => conv_std_logic_vector(24, 8),
52511 => conv_std_logic_vector(24, 8),
52512 => conv_std_logic_vector(25, 8),
52513 => conv_std_logic_vector(26, 8),
52514 => conv_std_logic_vector(27, 8),
52515 => conv_std_logic_vector(28, 8),
52516 => conv_std_logic_vector(28, 8),
52517 => conv_std_logic_vector(29, 8),
52518 => conv_std_logic_vector(30, 8),
52519 => conv_std_logic_vector(31, 8),
52520 => conv_std_logic_vector(32, 8),
52521 => conv_std_logic_vector(32, 8),
52522 => conv_std_logic_vector(33, 8),
52523 => conv_std_logic_vector(34, 8),
52524 => conv_std_logic_vector(35, 8),
52525 => conv_std_logic_vector(36, 8),
52526 => conv_std_logic_vector(36, 8),
52527 => conv_std_logic_vector(37, 8),
52528 => conv_std_logic_vector(38, 8),
52529 => conv_std_logic_vector(39, 8),
52530 => conv_std_logic_vector(40, 8),
52531 => conv_std_logic_vector(40, 8),
52532 => conv_std_logic_vector(41, 8),
52533 => conv_std_logic_vector(42, 8),
52534 => conv_std_logic_vector(43, 8),
52535 => conv_std_logic_vector(44, 8),
52536 => conv_std_logic_vector(44, 8),
52537 => conv_std_logic_vector(45, 8),
52538 => conv_std_logic_vector(46, 8),
52539 => conv_std_logic_vector(47, 8),
52540 => conv_std_logic_vector(48, 8),
52541 => conv_std_logic_vector(48, 8),
52542 => conv_std_logic_vector(49, 8),
52543 => conv_std_logic_vector(50, 8),
52544 => conv_std_logic_vector(51, 8),
52545 => conv_std_logic_vector(52, 8),
52546 => conv_std_logic_vector(52, 8),
52547 => conv_std_logic_vector(53, 8),
52548 => conv_std_logic_vector(54, 8),
52549 => conv_std_logic_vector(55, 8),
52550 => conv_std_logic_vector(56, 8),
52551 => conv_std_logic_vector(56, 8),
52552 => conv_std_logic_vector(57, 8),
52553 => conv_std_logic_vector(58, 8),
52554 => conv_std_logic_vector(59, 8),
52555 => conv_std_logic_vector(60, 8),
52556 => conv_std_logic_vector(60, 8),
52557 => conv_std_logic_vector(61, 8),
52558 => conv_std_logic_vector(62, 8),
52559 => conv_std_logic_vector(63, 8),
52560 => conv_std_logic_vector(64, 8),
52561 => conv_std_logic_vector(64, 8),
52562 => conv_std_logic_vector(65, 8),
52563 => conv_std_logic_vector(66, 8),
52564 => conv_std_logic_vector(67, 8),
52565 => conv_std_logic_vector(68, 8),
52566 => conv_std_logic_vector(68, 8),
52567 => conv_std_logic_vector(69, 8),
52568 => conv_std_logic_vector(70, 8),
52569 => conv_std_logic_vector(71, 8),
52570 => conv_std_logic_vector(72, 8),
52571 => conv_std_logic_vector(72, 8),
52572 => conv_std_logic_vector(73, 8),
52573 => conv_std_logic_vector(74, 8),
52574 => conv_std_logic_vector(75, 8),
52575 => conv_std_logic_vector(76, 8),
52576 => conv_std_logic_vector(76, 8),
52577 => conv_std_logic_vector(77, 8),
52578 => conv_std_logic_vector(78, 8),
52579 => conv_std_logic_vector(79, 8),
52580 => conv_std_logic_vector(80, 8),
52581 => conv_std_logic_vector(80, 8),
52582 => conv_std_logic_vector(81, 8),
52583 => conv_std_logic_vector(82, 8),
52584 => conv_std_logic_vector(83, 8),
52585 => conv_std_logic_vector(84, 8),
52586 => conv_std_logic_vector(84, 8),
52587 => conv_std_logic_vector(85, 8),
52588 => conv_std_logic_vector(86, 8),
52589 => conv_std_logic_vector(87, 8),
52590 => conv_std_logic_vector(88, 8),
52591 => conv_std_logic_vector(88, 8),
52592 => conv_std_logic_vector(89, 8),
52593 => conv_std_logic_vector(90, 8),
52594 => conv_std_logic_vector(91, 8),
52595 => conv_std_logic_vector(92, 8),
52596 => conv_std_logic_vector(92, 8),
52597 => conv_std_logic_vector(93, 8),
52598 => conv_std_logic_vector(94, 8),
52599 => conv_std_logic_vector(95, 8),
52600 => conv_std_logic_vector(96, 8),
52601 => conv_std_logic_vector(96, 8),
52602 => conv_std_logic_vector(97, 8),
52603 => conv_std_logic_vector(98, 8),
52604 => conv_std_logic_vector(99, 8),
52605 => conv_std_logic_vector(100, 8),
52606 => conv_std_logic_vector(100, 8),
52607 => conv_std_logic_vector(101, 8),
52608 => conv_std_logic_vector(102, 8),
52609 => conv_std_logic_vector(103, 8),
52610 => conv_std_logic_vector(104, 8),
52611 => conv_std_logic_vector(104, 8),
52612 => conv_std_logic_vector(105, 8),
52613 => conv_std_logic_vector(106, 8),
52614 => conv_std_logic_vector(107, 8),
52615 => conv_std_logic_vector(108, 8),
52616 => conv_std_logic_vector(108, 8),
52617 => conv_std_logic_vector(109, 8),
52618 => conv_std_logic_vector(110, 8),
52619 => conv_std_logic_vector(111, 8),
52620 => conv_std_logic_vector(112, 8),
52621 => conv_std_logic_vector(112, 8),
52622 => conv_std_logic_vector(113, 8),
52623 => conv_std_logic_vector(114, 8),
52624 => conv_std_logic_vector(115, 8),
52625 => conv_std_logic_vector(116, 8),
52626 => conv_std_logic_vector(116, 8),
52627 => conv_std_logic_vector(117, 8),
52628 => conv_std_logic_vector(118, 8),
52629 => conv_std_logic_vector(119, 8),
52630 => conv_std_logic_vector(120, 8),
52631 => conv_std_logic_vector(120, 8),
52632 => conv_std_logic_vector(121, 8),
52633 => conv_std_logic_vector(122, 8),
52634 => conv_std_logic_vector(123, 8),
52635 => conv_std_logic_vector(124, 8),
52636 => conv_std_logic_vector(124, 8),
52637 => conv_std_logic_vector(125, 8),
52638 => conv_std_logic_vector(126, 8),
52639 => conv_std_logic_vector(127, 8),
52640 => conv_std_logic_vector(128, 8),
52641 => conv_std_logic_vector(128, 8),
52642 => conv_std_logic_vector(129, 8),
52643 => conv_std_logic_vector(130, 8),
52644 => conv_std_logic_vector(131, 8),
52645 => conv_std_logic_vector(132, 8),
52646 => conv_std_logic_vector(132, 8),
52647 => conv_std_logic_vector(133, 8),
52648 => conv_std_logic_vector(134, 8),
52649 => conv_std_logic_vector(135, 8),
52650 => conv_std_logic_vector(136, 8),
52651 => conv_std_logic_vector(136, 8),
52652 => conv_std_logic_vector(137, 8),
52653 => conv_std_logic_vector(138, 8),
52654 => conv_std_logic_vector(139, 8),
52655 => conv_std_logic_vector(140, 8),
52656 => conv_std_logic_vector(140, 8),
52657 => conv_std_logic_vector(141, 8),
52658 => conv_std_logic_vector(142, 8),
52659 => conv_std_logic_vector(143, 8),
52660 => conv_std_logic_vector(144, 8),
52661 => conv_std_logic_vector(144, 8),
52662 => conv_std_logic_vector(145, 8),
52663 => conv_std_logic_vector(146, 8),
52664 => conv_std_logic_vector(147, 8),
52665 => conv_std_logic_vector(148, 8),
52666 => conv_std_logic_vector(148, 8),
52667 => conv_std_logic_vector(149, 8),
52668 => conv_std_logic_vector(150, 8),
52669 => conv_std_logic_vector(151, 8),
52670 => conv_std_logic_vector(152, 8),
52671 => conv_std_logic_vector(152, 8),
52672 => conv_std_logic_vector(153, 8),
52673 => conv_std_logic_vector(154, 8),
52674 => conv_std_logic_vector(155, 8),
52675 => conv_std_logic_vector(156, 8),
52676 => conv_std_logic_vector(156, 8),
52677 => conv_std_logic_vector(157, 8),
52678 => conv_std_logic_vector(158, 8),
52679 => conv_std_logic_vector(159, 8),
52680 => conv_std_logic_vector(160, 8),
52681 => conv_std_logic_vector(160, 8),
52682 => conv_std_logic_vector(161, 8),
52683 => conv_std_logic_vector(162, 8),
52684 => conv_std_logic_vector(163, 8),
52685 => conv_std_logic_vector(164, 8),
52686 => conv_std_logic_vector(164, 8),
52687 => conv_std_logic_vector(165, 8),
52688 => conv_std_logic_vector(166, 8),
52689 => conv_std_logic_vector(167, 8),
52690 => conv_std_logic_vector(168, 8),
52691 => conv_std_logic_vector(168, 8),
52692 => conv_std_logic_vector(169, 8),
52693 => conv_std_logic_vector(170, 8),
52694 => conv_std_logic_vector(171, 8),
52695 => conv_std_logic_vector(172, 8),
52696 => conv_std_logic_vector(172, 8),
52697 => conv_std_logic_vector(173, 8),
52698 => conv_std_logic_vector(174, 8),
52699 => conv_std_logic_vector(175, 8),
52700 => conv_std_logic_vector(176, 8),
52701 => conv_std_logic_vector(176, 8),
52702 => conv_std_logic_vector(177, 8),
52703 => conv_std_logic_vector(178, 8),
52704 => conv_std_logic_vector(179, 8),
52705 => conv_std_logic_vector(180, 8),
52706 => conv_std_logic_vector(180, 8),
52707 => conv_std_logic_vector(181, 8),
52708 => conv_std_logic_vector(182, 8),
52709 => conv_std_logic_vector(183, 8),
52710 => conv_std_logic_vector(184, 8),
52711 => conv_std_logic_vector(184, 8),
52712 => conv_std_logic_vector(185, 8),
52713 => conv_std_logic_vector(186, 8),
52714 => conv_std_logic_vector(187, 8),
52715 => conv_std_logic_vector(188, 8),
52716 => conv_std_logic_vector(188, 8),
52717 => conv_std_logic_vector(189, 8),
52718 => conv_std_logic_vector(190, 8),
52719 => conv_std_logic_vector(191, 8),
52720 => conv_std_logic_vector(192, 8),
52721 => conv_std_logic_vector(192, 8),
52722 => conv_std_logic_vector(193, 8),
52723 => conv_std_logic_vector(194, 8),
52724 => conv_std_logic_vector(195, 8),
52725 => conv_std_logic_vector(196, 8),
52726 => conv_std_logic_vector(196, 8),
52727 => conv_std_logic_vector(197, 8),
52728 => conv_std_logic_vector(198, 8),
52729 => conv_std_logic_vector(199, 8),
52730 => conv_std_logic_vector(200, 8),
52731 => conv_std_logic_vector(200, 8),
52732 => conv_std_logic_vector(201, 8),
52733 => conv_std_logic_vector(202, 8),
52734 => conv_std_logic_vector(203, 8),
52735 => conv_std_logic_vector(204, 8),
52736 => conv_std_logic_vector(0, 8),
52737 => conv_std_logic_vector(0, 8),
52738 => conv_std_logic_vector(1, 8),
52739 => conv_std_logic_vector(2, 8),
52740 => conv_std_logic_vector(3, 8),
52741 => conv_std_logic_vector(4, 8),
52742 => conv_std_logic_vector(4, 8),
52743 => conv_std_logic_vector(5, 8),
52744 => conv_std_logic_vector(6, 8),
52745 => conv_std_logic_vector(7, 8),
52746 => conv_std_logic_vector(8, 8),
52747 => conv_std_logic_vector(8, 8),
52748 => conv_std_logic_vector(9, 8),
52749 => conv_std_logic_vector(10, 8),
52750 => conv_std_logic_vector(11, 8),
52751 => conv_std_logic_vector(12, 8),
52752 => conv_std_logic_vector(12, 8),
52753 => conv_std_logic_vector(13, 8),
52754 => conv_std_logic_vector(14, 8),
52755 => conv_std_logic_vector(15, 8),
52756 => conv_std_logic_vector(16, 8),
52757 => conv_std_logic_vector(16, 8),
52758 => conv_std_logic_vector(17, 8),
52759 => conv_std_logic_vector(18, 8),
52760 => conv_std_logic_vector(19, 8),
52761 => conv_std_logic_vector(20, 8),
52762 => conv_std_logic_vector(20, 8),
52763 => conv_std_logic_vector(21, 8),
52764 => conv_std_logic_vector(22, 8),
52765 => conv_std_logic_vector(23, 8),
52766 => conv_std_logic_vector(24, 8),
52767 => conv_std_logic_vector(24, 8),
52768 => conv_std_logic_vector(25, 8),
52769 => conv_std_logic_vector(26, 8),
52770 => conv_std_logic_vector(27, 8),
52771 => conv_std_logic_vector(28, 8),
52772 => conv_std_logic_vector(28, 8),
52773 => conv_std_logic_vector(29, 8),
52774 => conv_std_logic_vector(30, 8),
52775 => conv_std_logic_vector(31, 8),
52776 => conv_std_logic_vector(32, 8),
52777 => conv_std_logic_vector(32, 8),
52778 => conv_std_logic_vector(33, 8),
52779 => conv_std_logic_vector(34, 8),
52780 => conv_std_logic_vector(35, 8),
52781 => conv_std_logic_vector(36, 8),
52782 => conv_std_logic_vector(37, 8),
52783 => conv_std_logic_vector(37, 8),
52784 => conv_std_logic_vector(38, 8),
52785 => conv_std_logic_vector(39, 8),
52786 => conv_std_logic_vector(40, 8),
52787 => conv_std_logic_vector(41, 8),
52788 => conv_std_logic_vector(41, 8),
52789 => conv_std_logic_vector(42, 8),
52790 => conv_std_logic_vector(43, 8),
52791 => conv_std_logic_vector(44, 8),
52792 => conv_std_logic_vector(45, 8),
52793 => conv_std_logic_vector(45, 8),
52794 => conv_std_logic_vector(46, 8),
52795 => conv_std_logic_vector(47, 8),
52796 => conv_std_logic_vector(48, 8),
52797 => conv_std_logic_vector(49, 8),
52798 => conv_std_logic_vector(49, 8),
52799 => conv_std_logic_vector(50, 8),
52800 => conv_std_logic_vector(51, 8),
52801 => conv_std_logic_vector(52, 8),
52802 => conv_std_logic_vector(53, 8),
52803 => conv_std_logic_vector(53, 8),
52804 => conv_std_logic_vector(54, 8),
52805 => conv_std_logic_vector(55, 8),
52806 => conv_std_logic_vector(56, 8),
52807 => conv_std_logic_vector(57, 8),
52808 => conv_std_logic_vector(57, 8),
52809 => conv_std_logic_vector(58, 8),
52810 => conv_std_logic_vector(59, 8),
52811 => conv_std_logic_vector(60, 8),
52812 => conv_std_logic_vector(61, 8),
52813 => conv_std_logic_vector(61, 8),
52814 => conv_std_logic_vector(62, 8),
52815 => conv_std_logic_vector(63, 8),
52816 => conv_std_logic_vector(64, 8),
52817 => conv_std_logic_vector(65, 8),
52818 => conv_std_logic_vector(65, 8),
52819 => conv_std_logic_vector(66, 8),
52820 => conv_std_logic_vector(67, 8),
52821 => conv_std_logic_vector(68, 8),
52822 => conv_std_logic_vector(69, 8),
52823 => conv_std_logic_vector(70, 8),
52824 => conv_std_logic_vector(70, 8),
52825 => conv_std_logic_vector(71, 8),
52826 => conv_std_logic_vector(72, 8),
52827 => conv_std_logic_vector(73, 8),
52828 => conv_std_logic_vector(74, 8),
52829 => conv_std_logic_vector(74, 8),
52830 => conv_std_logic_vector(75, 8),
52831 => conv_std_logic_vector(76, 8),
52832 => conv_std_logic_vector(77, 8),
52833 => conv_std_logic_vector(78, 8),
52834 => conv_std_logic_vector(78, 8),
52835 => conv_std_logic_vector(79, 8),
52836 => conv_std_logic_vector(80, 8),
52837 => conv_std_logic_vector(81, 8),
52838 => conv_std_logic_vector(82, 8),
52839 => conv_std_logic_vector(82, 8),
52840 => conv_std_logic_vector(83, 8),
52841 => conv_std_logic_vector(84, 8),
52842 => conv_std_logic_vector(85, 8),
52843 => conv_std_logic_vector(86, 8),
52844 => conv_std_logic_vector(86, 8),
52845 => conv_std_logic_vector(87, 8),
52846 => conv_std_logic_vector(88, 8),
52847 => conv_std_logic_vector(89, 8),
52848 => conv_std_logic_vector(90, 8),
52849 => conv_std_logic_vector(90, 8),
52850 => conv_std_logic_vector(91, 8),
52851 => conv_std_logic_vector(92, 8),
52852 => conv_std_logic_vector(93, 8),
52853 => conv_std_logic_vector(94, 8),
52854 => conv_std_logic_vector(94, 8),
52855 => conv_std_logic_vector(95, 8),
52856 => conv_std_logic_vector(96, 8),
52857 => conv_std_logic_vector(97, 8),
52858 => conv_std_logic_vector(98, 8),
52859 => conv_std_logic_vector(98, 8),
52860 => conv_std_logic_vector(99, 8),
52861 => conv_std_logic_vector(100, 8),
52862 => conv_std_logic_vector(101, 8),
52863 => conv_std_logic_vector(102, 8),
52864 => conv_std_logic_vector(103, 8),
52865 => conv_std_logic_vector(103, 8),
52866 => conv_std_logic_vector(104, 8),
52867 => conv_std_logic_vector(105, 8),
52868 => conv_std_logic_vector(106, 8),
52869 => conv_std_logic_vector(107, 8),
52870 => conv_std_logic_vector(107, 8),
52871 => conv_std_logic_vector(108, 8),
52872 => conv_std_logic_vector(109, 8),
52873 => conv_std_logic_vector(110, 8),
52874 => conv_std_logic_vector(111, 8),
52875 => conv_std_logic_vector(111, 8),
52876 => conv_std_logic_vector(112, 8),
52877 => conv_std_logic_vector(113, 8),
52878 => conv_std_logic_vector(114, 8),
52879 => conv_std_logic_vector(115, 8),
52880 => conv_std_logic_vector(115, 8),
52881 => conv_std_logic_vector(116, 8),
52882 => conv_std_logic_vector(117, 8),
52883 => conv_std_logic_vector(118, 8),
52884 => conv_std_logic_vector(119, 8),
52885 => conv_std_logic_vector(119, 8),
52886 => conv_std_logic_vector(120, 8),
52887 => conv_std_logic_vector(121, 8),
52888 => conv_std_logic_vector(122, 8),
52889 => conv_std_logic_vector(123, 8),
52890 => conv_std_logic_vector(123, 8),
52891 => conv_std_logic_vector(124, 8),
52892 => conv_std_logic_vector(125, 8),
52893 => conv_std_logic_vector(126, 8),
52894 => conv_std_logic_vector(127, 8),
52895 => conv_std_logic_vector(127, 8),
52896 => conv_std_logic_vector(128, 8),
52897 => conv_std_logic_vector(129, 8),
52898 => conv_std_logic_vector(130, 8),
52899 => conv_std_logic_vector(131, 8),
52900 => conv_std_logic_vector(131, 8),
52901 => conv_std_logic_vector(132, 8),
52902 => conv_std_logic_vector(133, 8),
52903 => conv_std_logic_vector(134, 8),
52904 => conv_std_logic_vector(135, 8),
52905 => conv_std_logic_vector(135, 8),
52906 => conv_std_logic_vector(136, 8),
52907 => conv_std_logic_vector(137, 8),
52908 => conv_std_logic_vector(138, 8),
52909 => conv_std_logic_vector(139, 8),
52910 => conv_std_logic_vector(140, 8),
52911 => conv_std_logic_vector(140, 8),
52912 => conv_std_logic_vector(141, 8),
52913 => conv_std_logic_vector(142, 8),
52914 => conv_std_logic_vector(143, 8),
52915 => conv_std_logic_vector(144, 8),
52916 => conv_std_logic_vector(144, 8),
52917 => conv_std_logic_vector(145, 8),
52918 => conv_std_logic_vector(146, 8),
52919 => conv_std_logic_vector(147, 8),
52920 => conv_std_logic_vector(148, 8),
52921 => conv_std_logic_vector(148, 8),
52922 => conv_std_logic_vector(149, 8),
52923 => conv_std_logic_vector(150, 8),
52924 => conv_std_logic_vector(151, 8),
52925 => conv_std_logic_vector(152, 8),
52926 => conv_std_logic_vector(152, 8),
52927 => conv_std_logic_vector(153, 8),
52928 => conv_std_logic_vector(154, 8),
52929 => conv_std_logic_vector(155, 8),
52930 => conv_std_logic_vector(156, 8),
52931 => conv_std_logic_vector(156, 8),
52932 => conv_std_logic_vector(157, 8),
52933 => conv_std_logic_vector(158, 8),
52934 => conv_std_logic_vector(159, 8),
52935 => conv_std_logic_vector(160, 8),
52936 => conv_std_logic_vector(160, 8),
52937 => conv_std_logic_vector(161, 8),
52938 => conv_std_logic_vector(162, 8),
52939 => conv_std_logic_vector(163, 8),
52940 => conv_std_logic_vector(164, 8),
52941 => conv_std_logic_vector(164, 8),
52942 => conv_std_logic_vector(165, 8),
52943 => conv_std_logic_vector(166, 8),
52944 => conv_std_logic_vector(167, 8),
52945 => conv_std_logic_vector(168, 8),
52946 => conv_std_logic_vector(168, 8),
52947 => conv_std_logic_vector(169, 8),
52948 => conv_std_logic_vector(170, 8),
52949 => conv_std_logic_vector(171, 8),
52950 => conv_std_logic_vector(172, 8),
52951 => conv_std_logic_vector(173, 8),
52952 => conv_std_logic_vector(173, 8),
52953 => conv_std_logic_vector(174, 8),
52954 => conv_std_logic_vector(175, 8),
52955 => conv_std_logic_vector(176, 8),
52956 => conv_std_logic_vector(177, 8),
52957 => conv_std_logic_vector(177, 8),
52958 => conv_std_logic_vector(178, 8),
52959 => conv_std_logic_vector(179, 8),
52960 => conv_std_logic_vector(180, 8),
52961 => conv_std_logic_vector(181, 8),
52962 => conv_std_logic_vector(181, 8),
52963 => conv_std_logic_vector(182, 8),
52964 => conv_std_logic_vector(183, 8),
52965 => conv_std_logic_vector(184, 8),
52966 => conv_std_logic_vector(185, 8),
52967 => conv_std_logic_vector(185, 8),
52968 => conv_std_logic_vector(186, 8),
52969 => conv_std_logic_vector(187, 8),
52970 => conv_std_logic_vector(188, 8),
52971 => conv_std_logic_vector(189, 8),
52972 => conv_std_logic_vector(189, 8),
52973 => conv_std_logic_vector(190, 8),
52974 => conv_std_logic_vector(191, 8),
52975 => conv_std_logic_vector(192, 8),
52976 => conv_std_logic_vector(193, 8),
52977 => conv_std_logic_vector(193, 8),
52978 => conv_std_logic_vector(194, 8),
52979 => conv_std_logic_vector(195, 8),
52980 => conv_std_logic_vector(196, 8),
52981 => conv_std_logic_vector(197, 8),
52982 => conv_std_logic_vector(197, 8),
52983 => conv_std_logic_vector(198, 8),
52984 => conv_std_logic_vector(199, 8),
52985 => conv_std_logic_vector(200, 8),
52986 => conv_std_logic_vector(201, 8),
52987 => conv_std_logic_vector(201, 8),
52988 => conv_std_logic_vector(202, 8),
52989 => conv_std_logic_vector(203, 8),
52990 => conv_std_logic_vector(204, 8),
52991 => conv_std_logic_vector(205, 8),
52992 => conv_std_logic_vector(0, 8),
52993 => conv_std_logic_vector(0, 8),
52994 => conv_std_logic_vector(1, 8),
52995 => conv_std_logic_vector(2, 8),
52996 => conv_std_logic_vector(3, 8),
52997 => conv_std_logic_vector(4, 8),
52998 => conv_std_logic_vector(4, 8),
52999 => conv_std_logic_vector(5, 8),
53000 => conv_std_logic_vector(6, 8),
53001 => conv_std_logic_vector(7, 8),
53002 => conv_std_logic_vector(8, 8),
53003 => conv_std_logic_vector(8, 8),
53004 => conv_std_logic_vector(9, 8),
53005 => conv_std_logic_vector(10, 8),
53006 => conv_std_logic_vector(11, 8),
53007 => conv_std_logic_vector(12, 8),
53008 => conv_std_logic_vector(12, 8),
53009 => conv_std_logic_vector(13, 8),
53010 => conv_std_logic_vector(14, 8),
53011 => conv_std_logic_vector(15, 8),
53012 => conv_std_logic_vector(16, 8),
53013 => conv_std_logic_vector(16, 8),
53014 => conv_std_logic_vector(17, 8),
53015 => conv_std_logic_vector(18, 8),
53016 => conv_std_logic_vector(19, 8),
53017 => conv_std_logic_vector(20, 8),
53018 => conv_std_logic_vector(21, 8),
53019 => conv_std_logic_vector(21, 8),
53020 => conv_std_logic_vector(22, 8),
53021 => conv_std_logic_vector(23, 8),
53022 => conv_std_logic_vector(24, 8),
53023 => conv_std_logic_vector(25, 8),
53024 => conv_std_logic_vector(25, 8),
53025 => conv_std_logic_vector(26, 8),
53026 => conv_std_logic_vector(27, 8),
53027 => conv_std_logic_vector(28, 8),
53028 => conv_std_logic_vector(29, 8),
53029 => conv_std_logic_vector(29, 8),
53030 => conv_std_logic_vector(30, 8),
53031 => conv_std_logic_vector(31, 8),
53032 => conv_std_logic_vector(32, 8),
53033 => conv_std_logic_vector(33, 8),
53034 => conv_std_logic_vector(33, 8),
53035 => conv_std_logic_vector(34, 8),
53036 => conv_std_logic_vector(35, 8),
53037 => conv_std_logic_vector(36, 8),
53038 => conv_std_logic_vector(37, 8),
53039 => conv_std_logic_vector(38, 8),
53040 => conv_std_logic_vector(38, 8),
53041 => conv_std_logic_vector(39, 8),
53042 => conv_std_logic_vector(40, 8),
53043 => conv_std_logic_vector(41, 8),
53044 => conv_std_logic_vector(42, 8),
53045 => conv_std_logic_vector(42, 8),
53046 => conv_std_logic_vector(43, 8),
53047 => conv_std_logic_vector(44, 8),
53048 => conv_std_logic_vector(45, 8),
53049 => conv_std_logic_vector(46, 8),
53050 => conv_std_logic_vector(46, 8),
53051 => conv_std_logic_vector(47, 8),
53052 => conv_std_logic_vector(48, 8),
53053 => conv_std_logic_vector(49, 8),
53054 => conv_std_logic_vector(50, 8),
53055 => conv_std_logic_vector(50, 8),
53056 => conv_std_logic_vector(51, 8),
53057 => conv_std_logic_vector(52, 8),
53058 => conv_std_logic_vector(53, 8),
53059 => conv_std_logic_vector(54, 8),
53060 => conv_std_logic_vector(54, 8),
53061 => conv_std_logic_vector(55, 8),
53062 => conv_std_logic_vector(56, 8),
53063 => conv_std_logic_vector(57, 8),
53064 => conv_std_logic_vector(58, 8),
53065 => conv_std_logic_vector(59, 8),
53066 => conv_std_logic_vector(59, 8),
53067 => conv_std_logic_vector(60, 8),
53068 => conv_std_logic_vector(61, 8),
53069 => conv_std_logic_vector(62, 8),
53070 => conv_std_logic_vector(63, 8),
53071 => conv_std_logic_vector(63, 8),
53072 => conv_std_logic_vector(64, 8),
53073 => conv_std_logic_vector(65, 8),
53074 => conv_std_logic_vector(66, 8),
53075 => conv_std_logic_vector(67, 8),
53076 => conv_std_logic_vector(67, 8),
53077 => conv_std_logic_vector(68, 8),
53078 => conv_std_logic_vector(69, 8),
53079 => conv_std_logic_vector(70, 8),
53080 => conv_std_logic_vector(71, 8),
53081 => conv_std_logic_vector(71, 8),
53082 => conv_std_logic_vector(72, 8),
53083 => conv_std_logic_vector(73, 8),
53084 => conv_std_logic_vector(74, 8),
53085 => conv_std_logic_vector(75, 8),
53086 => conv_std_logic_vector(76, 8),
53087 => conv_std_logic_vector(76, 8),
53088 => conv_std_logic_vector(77, 8),
53089 => conv_std_logic_vector(78, 8),
53090 => conv_std_logic_vector(79, 8),
53091 => conv_std_logic_vector(80, 8),
53092 => conv_std_logic_vector(80, 8),
53093 => conv_std_logic_vector(81, 8),
53094 => conv_std_logic_vector(82, 8),
53095 => conv_std_logic_vector(83, 8),
53096 => conv_std_logic_vector(84, 8),
53097 => conv_std_logic_vector(84, 8),
53098 => conv_std_logic_vector(85, 8),
53099 => conv_std_logic_vector(86, 8),
53100 => conv_std_logic_vector(87, 8),
53101 => conv_std_logic_vector(88, 8),
53102 => conv_std_logic_vector(88, 8),
53103 => conv_std_logic_vector(89, 8),
53104 => conv_std_logic_vector(90, 8),
53105 => conv_std_logic_vector(91, 8),
53106 => conv_std_logic_vector(92, 8),
53107 => conv_std_logic_vector(92, 8),
53108 => conv_std_logic_vector(93, 8),
53109 => conv_std_logic_vector(94, 8),
53110 => conv_std_logic_vector(95, 8),
53111 => conv_std_logic_vector(96, 8),
53112 => conv_std_logic_vector(97, 8),
53113 => conv_std_logic_vector(97, 8),
53114 => conv_std_logic_vector(98, 8),
53115 => conv_std_logic_vector(99, 8),
53116 => conv_std_logic_vector(100, 8),
53117 => conv_std_logic_vector(101, 8),
53118 => conv_std_logic_vector(101, 8),
53119 => conv_std_logic_vector(102, 8),
53120 => conv_std_logic_vector(103, 8),
53121 => conv_std_logic_vector(104, 8),
53122 => conv_std_logic_vector(105, 8),
53123 => conv_std_logic_vector(105, 8),
53124 => conv_std_logic_vector(106, 8),
53125 => conv_std_logic_vector(107, 8),
53126 => conv_std_logic_vector(108, 8),
53127 => conv_std_logic_vector(109, 8),
53128 => conv_std_logic_vector(109, 8),
53129 => conv_std_logic_vector(110, 8),
53130 => conv_std_logic_vector(111, 8),
53131 => conv_std_logic_vector(112, 8),
53132 => conv_std_logic_vector(113, 8),
53133 => conv_std_logic_vector(114, 8),
53134 => conv_std_logic_vector(114, 8),
53135 => conv_std_logic_vector(115, 8),
53136 => conv_std_logic_vector(116, 8),
53137 => conv_std_logic_vector(117, 8),
53138 => conv_std_logic_vector(118, 8),
53139 => conv_std_logic_vector(118, 8),
53140 => conv_std_logic_vector(119, 8),
53141 => conv_std_logic_vector(120, 8),
53142 => conv_std_logic_vector(121, 8),
53143 => conv_std_logic_vector(122, 8),
53144 => conv_std_logic_vector(122, 8),
53145 => conv_std_logic_vector(123, 8),
53146 => conv_std_logic_vector(124, 8),
53147 => conv_std_logic_vector(125, 8),
53148 => conv_std_logic_vector(126, 8),
53149 => conv_std_logic_vector(126, 8),
53150 => conv_std_logic_vector(127, 8),
53151 => conv_std_logic_vector(128, 8),
53152 => conv_std_logic_vector(129, 8),
53153 => conv_std_logic_vector(130, 8),
53154 => conv_std_logic_vector(130, 8),
53155 => conv_std_logic_vector(131, 8),
53156 => conv_std_logic_vector(132, 8),
53157 => conv_std_logic_vector(133, 8),
53158 => conv_std_logic_vector(134, 8),
53159 => conv_std_logic_vector(135, 8),
53160 => conv_std_logic_vector(135, 8),
53161 => conv_std_logic_vector(136, 8),
53162 => conv_std_logic_vector(137, 8),
53163 => conv_std_logic_vector(138, 8),
53164 => conv_std_logic_vector(139, 8),
53165 => conv_std_logic_vector(139, 8),
53166 => conv_std_logic_vector(140, 8),
53167 => conv_std_logic_vector(141, 8),
53168 => conv_std_logic_vector(142, 8),
53169 => conv_std_logic_vector(143, 8),
53170 => conv_std_logic_vector(143, 8),
53171 => conv_std_logic_vector(144, 8),
53172 => conv_std_logic_vector(145, 8),
53173 => conv_std_logic_vector(146, 8),
53174 => conv_std_logic_vector(147, 8),
53175 => conv_std_logic_vector(147, 8),
53176 => conv_std_logic_vector(148, 8),
53177 => conv_std_logic_vector(149, 8),
53178 => conv_std_logic_vector(150, 8),
53179 => conv_std_logic_vector(151, 8),
53180 => conv_std_logic_vector(152, 8),
53181 => conv_std_logic_vector(152, 8),
53182 => conv_std_logic_vector(153, 8),
53183 => conv_std_logic_vector(154, 8),
53184 => conv_std_logic_vector(155, 8),
53185 => conv_std_logic_vector(156, 8),
53186 => conv_std_logic_vector(156, 8),
53187 => conv_std_logic_vector(157, 8),
53188 => conv_std_logic_vector(158, 8),
53189 => conv_std_logic_vector(159, 8),
53190 => conv_std_logic_vector(160, 8),
53191 => conv_std_logic_vector(160, 8),
53192 => conv_std_logic_vector(161, 8),
53193 => conv_std_logic_vector(162, 8),
53194 => conv_std_logic_vector(163, 8),
53195 => conv_std_logic_vector(164, 8),
53196 => conv_std_logic_vector(164, 8),
53197 => conv_std_logic_vector(165, 8),
53198 => conv_std_logic_vector(166, 8),
53199 => conv_std_logic_vector(167, 8),
53200 => conv_std_logic_vector(168, 8),
53201 => conv_std_logic_vector(168, 8),
53202 => conv_std_logic_vector(169, 8),
53203 => conv_std_logic_vector(170, 8),
53204 => conv_std_logic_vector(171, 8),
53205 => conv_std_logic_vector(172, 8),
53206 => conv_std_logic_vector(173, 8),
53207 => conv_std_logic_vector(173, 8),
53208 => conv_std_logic_vector(174, 8),
53209 => conv_std_logic_vector(175, 8),
53210 => conv_std_logic_vector(176, 8),
53211 => conv_std_logic_vector(177, 8),
53212 => conv_std_logic_vector(177, 8),
53213 => conv_std_logic_vector(178, 8),
53214 => conv_std_logic_vector(179, 8),
53215 => conv_std_logic_vector(180, 8),
53216 => conv_std_logic_vector(181, 8),
53217 => conv_std_logic_vector(181, 8),
53218 => conv_std_logic_vector(182, 8),
53219 => conv_std_logic_vector(183, 8),
53220 => conv_std_logic_vector(184, 8),
53221 => conv_std_logic_vector(185, 8),
53222 => conv_std_logic_vector(185, 8),
53223 => conv_std_logic_vector(186, 8),
53224 => conv_std_logic_vector(187, 8),
53225 => conv_std_logic_vector(188, 8),
53226 => conv_std_logic_vector(189, 8),
53227 => conv_std_logic_vector(190, 8),
53228 => conv_std_logic_vector(190, 8),
53229 => conv_std_logic_vector(191, 8),
53230 => conv_std_logic_vector(192, 8),
53231 => conv_std_logic_vector(193, 8),
53232 => conv_std_logic_vector(194, 8),
53233 => conv_std_logic_vector(194, 8),
53234 => conv_std_logic_vector(195, 8),
53235 => conv_std_logic_vector(196, 8),
53236 => conv_std_logic_vector(197, 8),
53237 => conv_std_logic_vector(198, 8),
53238 => conv_std_logic_vector(198, 8),
53239 => conv_std_logic_vector(199, 8),
53240 => conv_std_logic_vector(200, 8),
53241 => conv_std_logic_vector(201, 8),
53242 => conv_std_logic_vector(202, 8),
53243 => conv_std_logic_vector(202, 8),
53244 => conv_std_logic_vector(203, 8),
53245 => conv_std_logic_vector(204, 8),
53246 => conv_std_logic_vector(205, 8),
53247 => conv_std_logic_vector(206, 8),
53248 => conv_std_logic_vector(0, 8),
53249 => conv_std_logic_vector(0, 8),
53250 => conv_std_logic_vector(1, 8),
53251 => conv_std_logic_vector(2, 8),
53252 => conv_std_logic_vector(3, 8),
53253 => conv_std_logic_vector(4, 8),
53254 => conv_std_logic_vector(4, 8),
53255 => conv_std_logic_vector(5, 8),
53256 => conv_std_logic_vector(6, 8),
53257 => conv_std_logic_vector(7, 8),
53258 => conv_std_logic_vector(8, 8),
53259 => conv_std_logic_vector(8, 8),
53260 => conv_std_logic_vector(9, 8),
53261 => conv_std_logic_vector(10, 8),
53262 => conv_std_logic_vector(11, 8),
53263 => conv_std_logic_vector(12, 8),
53264 => conv_std_logic_vector(13, 8),
53265 => conv_std_logic_vector(13, 8),
53266 => conv_std_logic_vector(14, 8),
53267 => conv_std_logic_vector(15, 8),
53268 => conv_std_logic_vector(16, 8),
53269 => conv_std_logic_vector(17, 8),
53270 => conv_std_logic_vector(17, 8),
53271 => conv_std_logic_vector(18, 8),
53272 => conv_std_logic_vector(19, 8),
53273 => conv_std_logic_vector(20, 8),
53274 => conv_std_logic_vector(21, 8),
53275 => conv_std_logic_vector(21, 8),
53276 => conv_std_logic_vector(22, 8),
53277 => conv_std_logic_vector(23, 8),
53278 => conv_std_logic_vector(24, 8),
53279 => conv_std_logic_vector(25, 8),
53280 => conv_std_logic_vector(26, 8),
53281 => conv_std_logic_vector(26, 8),
53282 => conv_std_logic_vector(27, 8),
53283 => conv_std_logic_vector(28, 8),
53284 => conv_std_logic_vector(29, 8),
53285 => conv_std_logic_vector(30, 8),
53286 => conv_std_logic_vector(30, 8),
53287 => conv_std_logic_vector(31, 8),
53288 => conv_std_logic_vector(32, 8),
53289 => conv_std_logic_vector(33, 8),
53290 => conv_std_logic_vector(34, 8),
53291 => conv_std_logic_vector(34, 8),
53292 => conv_std_logic_vector(35, 8),
53293 => conv_std_logic_vector(36, 8),
53294 => conv_std_logic_vector(37, 8),
53295 => conv_std_logic_vector(38, 8),
53296 => conv_std_logic_vector(39, 8),
53297 => conv_std_logic_vector(39, 8),
53298 => conv_std_logic_vector(40, 8),
53299 => conv_std_logic_vector(41, 8),
53300 => conv_std_logic_vector(42, 8),
53301 => conv_std_logic_vector(43, 8),
53302 => conv_std_logic_vector(43, 8),
53303 => conv_std_logic_vector(44, 8),
53304 => conv_std_logic_vector(45, 8),
53305 => conv_std_logic_vector(46, 8),
53306 => conv_std_logic_vector(47, 8),
53307 => conv_std_logic_vector(47, 8),
53308 => conv_std_logic_vector(48, 8),
53309 => conv_std_logic_vector(49, 8),
53310 => conv_std_logic_vector(50, 8),
53311 => conv_std_logic_vector(51, 8),
53312 => conv_std_logic_vector(52, 8),
53313 => conv_std_logic_vector(52, 8),
53314 => conv_std_logic_vector(53, 8),
53315 => conv_std_logic_vector(54, 8),
53316 => conv_std_logic_vector(55, 8),
53317 => conv_std_logic_vector(56, 8),
53318 => conv_std_logic_vector(56, 8),
53319 => conv_std_logic_vector(57, 8),
53320 => conv_std_logic_vector(58, 8),
53321 => conv_std_logic_vector(59, 8),
53322 => conv_std_logic_vector(60, 8),
53323 => conv_std_logic_vector(60, 8),
53324 => conv_std_logic_vector(61, 8),
53325 => conv_std_logic_vector(62, 8),
53326 => conv_std_logic_vector(63, 8),
53327 => conv_std_logic_vector(64, 8),
53328 => conv_std_logic_vector(65, 8),
53329 => conv_std_logic_vector(65, 8),
53330 => conv_std_logic_vector(66, 8),
53331 => conv_std_logic_vector(67, 8),
53332 => conv_std_logic_vector(68, 8),
53333 => conv_std_logic_vector(69, 8),
53334 => conv_std_logic_vector(69, 8),
53335 => conv_std_logic_vector(70, 8),
53336 => conv_std_logic_vector(71, 8),
53337 => conv_std_logic_vector(72, 8),
53338 => conv_std_logic_vector(73, 8),
53339 => conv_std_logic_vector(73, 8),
53340 => conv_std_logic_vector(74, 8),
53341 => conv_std_logic_vector(75, 8),
53342 => conv_std_logic_vector(76, 8),
53343 => conv_std_logic_vector(77, 8),
53344 => conv_std_logic_vector(78, 8),
53345 => conv_std_logic_vector(78, 8),
53346 => conv_std_logic_vector(79, 8),
53347 => conv_std_logic_vector(80, 8),
53348 => conv_std_logic_vector(81, 8),
53349 => conv_std_logic_vector(82, 8),
53350 => conv_std_logic_vector(82, 8),
53351 => conv_std_logic_vector(83, 8),
53352 => conv_std_logic_vector(84, 8),
53353 => conv_std_logic_vector(85, 8),
53354 => conv_std_logic_vector(86, 8),
53355 => conv_std_logic_vector(86, 8),
53356 => conv_std_logic_vector(87, 8),
53357 => conv_std_logic_vector(88, 8),
53358 => conv_std_logic_vector(89, 8),
53359 => conv_std_logic_vector(90, 8),
53360 => conv_std_logic_vector(91, 8),
53361 => conv_std_logic_vector(91, 8),
53362 => conv_std_logic_vector(92, 8),
53363 => conv_std_logic_vector(93, 8),
53364 => conv_std_logic_vector(94, 8),
53365 => conv_std_logic_vector(95, 8),
53366 => conv_std_logic_vector(95, 8),
53367 => conv_std_logic_vector(96, 8),
53368 => conv_std_logic_vector(97, 8),
53369 => conv_std_logic_vector(98, 8),
53370 => conv_std_logic_vector(99, 8),
53371 => conv_std_logic_vector(99, 8),
53372 => conv_std_logic_vector(100, 8),
53373 => conv_std_logic_vector(101, 8),
53374 => conv_std_logic_vector(102, 8),
53375 => conv_std_logic_vector(103, 8),
53376 => conv_std_logic_vector(104, 8),
53377 => conv_std_logic_vector(104, 8),
53378 => conv_std_logic_vector(105, 8),
53379 => conv_std_logic_vector(106, 8),
53380 => conv_std_logic_vector(107, 8),
53381 => conv_std_logic_vector(108, 8),
53382 => conv_std_logic_vector(108, 8),
53383 => conv_std_logic_vector(109, 8),
53384 => conv_std_logic_vector(110, 8),
53385 => conv_std_logic_vector(111, 8),
53386 => conv_std_logic_vector(112, 8),
53387 => conv_std_logic_vector(112, 8),
53388 => conv_std_logic_vector(113, 8),
53389 => conv_std_logic_vector(114, 8),
53390 => conv_std_logic_vector(115, 8),
53391 => conv_std_logic_vector(116, 8),
53392 => conv_std_logic_vector(117, 8),
53393 => conv_std_logic_vector(117, 8),
53394 => conv_std_logic_vector(118, 8),
53395 => conv_std_logic_vector(119, 8),
53396 => conv_std_logic_vector(120, 8),
53397 => conv_std_logic_vector(121, 8),
53398 => conv_std_logic_vector(121, 8),
53399 => conv_std_logic_vector(122, 8),
53400 => conv_std_logic_vector(123, 8),
53401 => conv_std_logic_vector(124, 8),
53402 => conv_std_logic_vector(125, 8),
53403 => conv_std_logic_vector(125, 8),
53404 => conv_std_logic_vector(126, 8),
53405 => conv_std_logic_vector(127, 8),
53406 => conv_std_logic_vector(128, 8),
53407 => conv_std_logic_vector(129, 8),
53408 => conv_std_logic_vector(130, 8),
53409 => conv_std_logic_vector(130, 8),
53410 => conv_std_logic_vector(131, 8),
53411 => conv_std_logic_vector(132, 8),
53412 => conv_std_logic_vector(133, 8),
53413 => conv_std_logic_vector(134, 8),
53414 => conv_std_logic_vector(134, 8),
53415 => conv_std_logic_vector(135, 8),
53416 => conv_std_logic_vector(136, 8),
53417 => conv_std_logic_vector(137, 8),
53418 => conv_std_logic_vector(138, 8),
53419 => conv_std_logic_vector(138, 8),
53420 => conv_std_logic_vector(139, 8),
53421 => conv_std_logic_vector(140, 8),
53422 => conv_std_logic_vector(141, 8),
53423 => conv_std_logic_vector(142, 8),
53424 => conv_std_logic_vector(143, 8),
53425 => conv_std_logic_vector(143, 8),
53426 => conv_std_logic_vector(144, 8),
53427 => conv_std_logic_vector(145, 8),
53428 => conv_std_logic_vector(146, 8),
53429 => conv_std_logic_vector(147, 8),
53430 => conv_std_logic_vector(147, 8),
53431 => conv_std_logic_vector(148, 8),
53432 => conv_std_logic_vector(149, 8),
53433 => conv_std_logic_vector(150, 8),
53434 => conv_std_logic_vector(151, 8),
53435 => conv_std_logic_vector(151, 8),
53436 => conv_std_logic_vector(152, 8),
53437 => conv_std_logic_vector(153, 8),
53438 => conv_std_logic_vector(154, 8),
53439 => conv_std_logic_vector(155, 8),
53440 => conv_std_logic_vector(156, 8),
53441 => conv_std_logic_vector(156, 8),
53442 => conv_std_logic_vector(157, 8),
53443 => conv_std_logic_vector(158, 8),
53444 => conv_std_logic_vector(159, 8),
53445 => conv_std_logic_vector(160, 8),
53446 => conv_std_logic_vector(160, 8),
53447 => conv_std_logic_vector(161, 8),
53448 => conv_std_logic_vector(162, 8),
53449 => conv_std_logic_vector(163, 8),
53450 => conv_std_logic_vector(164, 8),
53451 => conv_std_logic_vector(164, 8),
53452 => conv_std_logic_vector(165, 8),
53453 => conv_std_logic_vector(166, 8),
53454 => conv_std_logic_vector(167, 8),
53455 => conv_std_logic_vector(168, 8),
53456 => conv_std_logic_vector(169, 8),
53457 => conv_std_logic_vector(169, 8),
53458 => conv_std_logic_vector(170, 8),
53459 => conv_std_logic_vector(171, 8),
53460 => conv_std_logic_vector(172, 8),
53461 => conv_std_logic_vector(173, 8),
53462 => conv_std_logic_vector(173, 8),
53463 => conv_std_logic_vector(174, 8),
53464 => conv_std_logic_vector(175, 8),
53465 => conv_std_logic_vector(176, 8),
53466 => conv_std_logic_vector(177, 8),
53467 => conv_std_logic_vector(177, 8),
53468 => conv_std_logic_vector(178, 8),
53469 => conv_std_logic_vector(179, 8),
53470 => conv_std_logic_vector(180, 8),
53471 => conv_std_logic_vector(181, 8),
53472 => conv_std_logic_vector(182, 8),
53473 => conv_std_logic_vector(182, 8),
53474 => conv_std_logic_vector(183, 8),
53475 => conv_std_logic_vector(184, 8),
53476 => conv_std_logic_vector(185, 8),
53477 => conv_std_logic_vector(186, 8),
53478 => conv_std_logic_vector(186, 8),
53479 => conv_std_logic_vector(187, 8),
53480 => conv_std_logic_vector(188, 8),
53481 => conv_std_logic_vector(189, 8),
53482 => conv_std_logic_vector(190, 8),
53483 => conv_std_logic_vector(190, 8),
53484 => conv_std_logic_vector(191, 8),
53485 => conv_std_logic_vector(192, 8),
53486 => conv_std_logic_vector(193, 8),
53487 => conv_std_logic_vector(194, 8),
53488 => conv_std_logic_vector(195, 8),
53489 => conv_std_logic_vector(195, 8),
53490 => conv_std_logic_vector(196, 8),
53491 => conv_std_logic_vector(197, 8),
53492 => conv_std_logic_vector(198, 8),
53493 => conv_std_logic_vector(199, 8),
53494 => conv_std_logic_vector(199, 8),
53495 => conv_std_logic_vector(200, 8),
53496 => conv_std_logic_vector(201, 8),
53497 => conv_std_logic_vector(202, 8),
53498 => conv_std_logic_vector(203, 8),
53499 => conv_std_logic_vector(203, 8),
53500 => conv_std_logic_vector(204, 8),
53501 => conv_std_logic_vector(205, 8),
53502 => conv_std_logic_vector(206, 8),
53503 => conv_std_logic_vector(207, 8),
53504 => conv_std_logic_vector(0, 8),
53505 => conv_std_logic_vector(0, 8),
53506 => conv_std_logic_vector(1, 8),
53507 => conv_std_logic_vector(2, 8),
53508 => conv_std_logic_vector(3, 8),
53509 => conv_std_logic_vector(4, 8),
53510 => conv_std_logic_vector(4, 8),
53511 => conv_std_logic_vector(5, 8),
53512 => conv_std_logic_vector(6, 8),
53513 => conv_std_logic_vector(7, 8),
53514 => conv_std_logic_vector(8, 8),
53515 => conv_std_logic_vector(8, 8),
53516 => conv_std_logic_vector(9, 8),
53517 => conv_std_logic_vector(10, 8),
53518 => conv_std_logic_vector(11, 8),
53519 => conv_std_logic_vector(12, 8),
53520 => conv_std_logic_vector(13, 8),
53521 => conv_std_logic_vector(13, 8),
53522 => conv_std_logic_vector(14, 8),
53523 => conv_std_logic_vector(15, 8),
53524 => conv_std_logic_vector(16, 8),
53525 => conv_std_logic_vector(17, 8),
53526 => conv_std_logic_vector(17, 8),
53527 => conv_std_logic_vector(18, 8),
53528 => conv_std_logic_vector(19, 8),
53529 => conv_std_logic_vector(20, 8),
53530 => conv_std_logic_vector(21, 8),
53531 => conv_std_logic_vector(22, 8),
53532 => conv_std_logic_vector(22, 8),
53533 => conv_std_logic_vector(23, 8),
53534 => conv_std_logic_vector(24, 8),
53535 => conv_std_logic_vector(25, 8),
53536 => conv_std_logic_vector(26, 8),
53537 => conv_std_logic_vector(26, 8),
53538 => conv_std_logic_vector(27, 8),
53539 => conv_std_logic_vector(28, 8),
53540 => conv_std_logic_vector(29, 8),
53541 => conv_std_logic_vector(30, 8),
53542 => conv_std_logic_vector(31, 8),
53543 => conv_std_logic_vector(31, 8),
53544 => conv_std_logic_vector(32, 8),
53545 => conv_std_logic_vector(33, 8),
53546 => conv_std_logic_vector(34, 8),
53547 => conv_std_logic_vector(35, 8),
53548 => conv_std_logic_vector(35, 8),
53549 => conv_std_logic_vector(36, 8),
53550 => conv_std_logic_vector(37, 8),
53551 => conv_std_logic_vector(38, 8),
53552 => conv_std_logic_vector(39, 8),
53553 => conv_std_logic_vector(40, 8),
53554 => conv_std_logic_vector(40, 8),
53555 => conv_std_logic_vector(41, 8),
53556 => conv_std_logic_vector(42, 8),
53557 => conv_std_logic_vector(43, 8),
53558 => conv_std_logic_vector(44, 8),
53559 => conv_std_logic_vector(44, 8),
53560 => conv_std_logic_vector(45, 8),
53561 => conv_std_logic_vector(46, 8),
53562 => conv_std_logic_vector(47, 8),
53563 => conv_std_logic_vector(48, 8),
53564 => conv_std_logic_vector(48, 8),
53565 => conv_std_logic_vector(49, 8),
53566 => conv_std_logic_vector(50, 8),
53567 => conv_std_logic_vector(51, 8),
53568 => conv_std_logic_vector(52, 8),
53569 => conv_std_logic_vector(53, 8),
53570 => conv_std_logic_vector(53, 8),
53571 => conv_std_logic_vector(54, 8),
53572 => conv_std_logic_vector(55, 8),
53573 => conv_std_logic_vector(56, 8),
53574 => conv_std_logic_vector(57, 8),
53575 => conv_std_logic_vector(57, 8),
53576 => conv_std_logic_vector(58, 8),
53577 => conv_std_logic_vector(59, 8),
53578 => conv_std_logic_vector(60, 8),
53579 => conv_std_logic_vector(61, 8),
53580 => conv_std_logic_vector(62, 8),
53581 => conv_std_logic_vector(62, 8),
53582 => conv_std_logic_vector(63, 8),
53583 => conv_std_logic_vector(64, 8),
53584 => conv_std_logic_vector(65, 8),
53585 => conv_std_logic_vector(66, 8),
53586 => conv_std_logic_vector(66, 8),
53587 => conv_std_logic_vector(67, 8),
53588 => conv_std_logic_vector(68, 8),
53589 => conv_std_logic_vector(69, 8),
53590 => conv_std_logic_vector(70, 8),
53591 => conv_std_logic_vector(71, 8),
53592 => conv_std_logic_vector(71, 8),
53593 => conv_std_logic_vector(72, 8),
53594 => conv_std_logic_vector(73, 8),
53595 => conv_std_logic_vector(74, 8),
53596 => conv_std_logic_vector(75, 8),
53597 => conv_std_logic_vector(75, 8),
53598 => conv_std_logic_vector(76, 8),
53599 => conv_std_logic_vector(77, 8),
53600 => conv_std_logic_vector(78, 8),
53601 => conv_std_logic_vector(79, 8),
53602 => conv_std_logic_vector(80, 8),
53603 => conv_std_logic_vector(80, 8),
53604 => conv_std_logic_vector(81, 8),
53605 => conv_std_logic_vector(82, 8),
53606 => conv_std_logic_vector(83, 8),
53607 => conv_std_logic_vector(84, 8),
53608 => conv_std_logic_vector(84, 8),
53609 => conv_std_logic_vector(85, 8),
53610 => conv_std_logic_vector(86, 8),
53611 => conv_std_logic_vector(87, 8),
53612 => conv_std_logic_vector(88, 8),
53613 => conv_std_logic_vector(88, 8),
53614 => conv_std_logic_vector(89, 8),
53615 => conv_std_logic_vector(90, 8),
53616 => conv_std_logic_vector(91, 8),
53617 => conv_std_logic_vector(92, 8),
53618 => conv_std_logic_vector(93, 8),
53619 => conv_std_logic_vector(93, 8),
53620 => conv_std_logic_vector(94, 8),
53621 => conv_std_logic_vector(95, 8),
53622 => conv_std_logic_vector(96, 8),
53623 => conv_std_logic_vector(97, 8),
53624 => conv_std_logic_vector(97, 8),
53625 => conv_std_logic_vector(98, 8),
53626 => conv_std_logic_vector(99, 8),
53627 => conv_std_logic_vector(100, 8),
53628 => conv_std_logic_vector(101, 8),
53629 => conv_std_logic_vector(102, 8),
53630 => conv_std_logic_vector(102, 8),
53631 => conv_std_logic_vector(103, 8),
53632 => conv_std_logic_vector(104, 8),
53633 => conv_std_logic_vector(105, 8),
53634 => conv_std_logic_vector(106, 8),
53635 => conv_std_logic_vector(106, 8),
53636 => conv_std_logic_vector(107, 8),
53637 => conv_std_logic_vector(108, 8),
53638 => conv_std_logic_vector(109, 8),
53639 => conv_std_logic_vector(110, 8),
53640 => conv_std_logic_vector(111, 8),
53641 => conv_std_logic_vector(111, 8),
53642 => conv_std_logic_vector(112, 8),
53643 => conv_std_logic_vector(113, 8),
53644 => conv_std_logic_vector(114, 8),
53645 => conv_std_logic_vector(115, 8),
53646 => conv_std_logic_vector(115, 8),
53647 => conv_std_logic_vector(116, 8),
53648 => conv_std_logic_vector(117, 8),
53649 => conv_std_logic_vector(118, 8),
53650 => conv_std_logic_vector(119, 8),
53651 => conv_std_logic_vector(120, 8),
53652 => conv_std_logic_vector(120, 8),
53653 => conv_std_logic_vector(121, 8),
53654 => conv_std_logic_vector(122, 8),
53655 => conv_std_logic_vector(123, 8),
53656 => conv_std_logic_vector(124, 8),
53657 => conv_std_logic_vector(124, 8),
53658 => conv_std_logic_vector(125, 8),
53659 => conv_std_logic_vector(126, 8),
53660 => conv_std_logic_vector(127, 8),
53661 => conv_std_logic_vector(128, 8),
53662 => conv_std_logic_vector(128, 8),
53663 => conv_std_logic_vector(129, 8),
53664 => conv_std_logic_vector(130, 8),
53665 => conv_std_logic_vector(131, 8),
53666 => conv_std_logic_vector(132, 8),
53667 => conv_std_logic_vector(133, 8),
53668 => conv_std_logic_vector(133, 8),
53669 => conv_std_logic_vector(134, 8),
53670 => conv_std_logic_vector(135, 8),
53671 => conv_std_logic_vector(136, 8),
53672 => conv_std_logic_vector(137, 8),
53673 => conv_std_logic_vector(137, 8),
53674 => conv_std_logic_vector(138, 8),
53675 => conv_std_logic_vector(139, 8),
53676 => conv_std_logic_vector(140, 8),
53677 => conv_std_logic_vector(141, 8),
53678 => conv_std_logic_vector(142, 8),
53679 => conv_std_logic_vector(142, 8),
53680 => conv_std_logic_vector(143, 8),
53681 => conv_std_logic_vector(144, 8),
53682 => conv_std_logic_vector(145, 8),
53683 => conv_std_logic_vector(146, 8),
53684 => conv_std_logic_vector(146, 8),
53685 => conv_std_logic_vector(147, 8),
53686 => conv_std_logic_vector(148, 8),
53687 => conv_std_logic_vector(149, 8),
53688 => conv_std_logic_vector(150, 8),
53689 => conv_std_logic_vector(151, 8),
53690 => conv_std_logic_vector(151, 8),
53691 => conv_std_logic_vector(152, 8),
53692 => conv_std_logic_vector(153, 8),
53693 => conv_std_logic_vector(154, 8),
53694 => conv_std_logic_vector(155, 8),
53695 => conv_std_logic_vector(155, 8),
53696 => conv_std_logic_vector(156, 8),
53697 => conv_std_logic_vector(157, 8),
53698 => conv_std_logic_vector(158, 8),
53699 => conv_std_logic_vector(159, 8),
53700 => conv_std_logic_vector(160, 8),
53701 => conv_std_logic_vector(160, 8),
53702 => conv_std_logic_vector(161, 8),
53703 => conv_std_logic_vector(162, 8),
53704 => conv_std_logic_vector(163, 8),
53705 => conv_std_logic_vector(164, 8),
53706 => conv_std_logic_vector(164, 8),
53707 => conv_std_logic_vector(165, 8),
53708 => conv_std_logic_vector(166, 8),
53709 => conv_std_logic_vector(167, 8),
53710 => conv_std_logic_vector(168, 8),
53711 => conv_std_logic_vector(168, 8),
53712 => conv_std_logic_vector(169, 8),
53713 => conv_std_logic_vector(170, 8),
53714 => conv_std_logic_vector(171, 8),
53715 => conv_std_logic_vector(172, 8),
53716 => conv_std_logic_vector(173, 8),
53717 => conv_std_logic_vector(173, 8),
53718 => conv_std_logic_vector(174, 8),
53719 => conv_std_logic_vector(175, 8),
53720 => conv_std_logic_vector(176, 8),
53721 => conv_std_logic_vector(177, 8),
53722 => conv_std_logic_vector(177, 8),
53723 => conv_std_logic_vector(178, 8),
53724 => conv_std_logic_vector(179, 8),
53725 => conv_std_logic_vector(180, 8),
53726 => conv_std_logic_vector(181, 8),
53727 => conv_std_logic_vector(182, 8),
53728 => conv_std_logic_vector(182, 8),
53729 => conv_std_logic_vector(183, 8),
53730 => conv_std_logic_vector(184, 8),
53731 => conv_std_logic_vector(185, 8),
53732 => conv_std_logic_vector(186, 8),
53733 => conv_std_logic_vector(186, 8),
53734 => conv_std_logic_vector(187, 8),
53735 => conv_std_logic_vector(188, 8),
53736 => conv_std_logic_vector(189, 8),
53737 => conv_std_logic_vector(190, 8),
53738 => conv_std_logic_vector(191, 8),
53739 => conv_std_logic_vector(191, 8),
53740 => conv_std_logic_vector(192, 8),
53741 => conv_std_logic_vector(193, 8),
53742 => conv_std_logic_vector(194, 8),
53743 => conv_std_logic_vector(195, 8),
53744 => conv_std_logic_vector(195, 8),
53745 => conv_std_logic_vector(196, 8),
53746 => conv_std_logic_vector(197, 8),
53747 => conv_std_logic_vector(198, 8),
53748 => conv_std_logic_vector(199, 8),
53749 => conv_std_logic_vector(200, 8),
53750 => conv_std_logic_vector(200, 8),
53751 => conv_std_logic_vector(201, 8),
53752 => conv_std_logic_vector(202, 8),
53753 => conv_std_logic_vector(203, 8),
53754 => conv_std_logic_vector(204, 8),
53755 => conv_std_logic_vector(204, 8),
53756 => conv_std_logic_vector(205, 8),
53757 => conv_std_logic_vector(206, 8),
53758 => conv_std_logic_vector(207, 8),
53759 => conv_std_logic_vector(208, 8),
53760 => conv_std_logic_vector(0, 8),
53761 => conv_std_logic_vector(0, 8),
53762 => conv_std_logic_vector(1, 8),
53763 => conv_std_logic_vector(2, 8),
53764 => conv_std_logic_vector(3, 8),
53765 => conv_std_logic_vector(4, 8),
53766 => conv_std_logic_vector(4, 8),
53767 => conv_std_logic_vector(5, 8),
53768 => conv_std_logic_vector(6, 8),
53769 => conv_std_logic_vector(7, 8),
53770 => conv_std_logic_vector(8, 8),
53771 => conv_std_logic_vector(9, 8),
53772 => conv_std_logic_vector(9, 8),
53773 => conv_std_logic_vector(10, 8),
53774 => conv_std_logic_vector(11, 8),
53775 => conv_std_logic_vector(12, 8),
53776 => conv_std_logic_vector(13, 8),
53777 => conv_std_logic_vector(13, 8),
53778 => conv_std_logic_vector(14, 8),
53779 => conv_std_logic_vector(15, 8),
53780 => conv_std_logic_vector(16, 8),
53781 => conv_std_logic_vector(17, 8),
53782 => conv_std_logic_vector(18, 8),
53783 => conv_std_logic_vector(18, 8),
53784 => conv_std_logic_vector(19, 8),
53785 => conv_std_logic_vector(20, 8),
53786 => conv_std_logic_vector(21, 8),
53787 => conv_std_logic_vector(22, 8),
53788 => conv_std_logic_vector(22, 8),
53789 => conv_std_logic_vector(23, 8),
53790 => conv_std_logic_vector(24, 8),
53791 => conv_std_logic_vector(25, 8),
53792 => conv_std_logic_vector(26, 8),
53793 => conv_std_logic_vector(27, 8),
53794 => conv_std_logic_vector(27, 8),
53795 => conv_std_logic_vector(28, 8),
53796 => conv_std_logic_vector(29, 8),
53797 => conv_std_logic_vector(30, 8),
53798 => conv_std_logic_vector(31, 8),
53799 => conv_std_logic_vector(31, 8),
53800 => conv_std_logic_vector(32, 8),
53801 => conv_std_logic_vector(33, 8),
53802 => conv_std_logic_vector(34, 8),
53803 => conv_std_logic_vector(35, 8),
53804 => conv_std_logic_vector(36, 8),
53805 => conv_std_logic_vector(36, 8),
53806 => conv_std_logic_vector(37, 8),
53807 => conv_std_logic_vector(38, 8),
53808 => conv_std_logic_vector(39, 8),
53809 => conv_std_logic_vector(40, 8),
53810 => conv_std_logic_vector(41, 8),
53811 => conv_std_logic_vector(41, 8),
53812 => conv_std_logic_vector(42, 8),
53813 => conv_std_logic_vector(43, 8),
53814 => conv_std_logic_vector(44, 8),
53815 => conv_std_logic_vector(45, 8),
53816 => conv_std_logic_vector(45, 8),
53817 => conv_std_logic_vector(46, 8),
53818 => conv_std_logic_vector(47, 8),
53819 => conv_std_logic_vector(48, 8),
53820 => conv_std_logic_vector(49, 8),
53821 => conv_std_logic_vector(50, 8),
53822 => conv_std_logic_vector(50, 8),
53823 => conv_std_logic_vector(51, 8),
53824 => conv_std_logic_vector(52, 8),
53825 => conv_std_logic_vector(53, 8),
53826 => conv_std_logic_vector(54, 8),
53827 => conv_std_logic_vector(54, 8),
53828 => conv_std_logic_vector(55, 8),
53829 => conv_std_logic_vector(56, 8),
53830 => conv_std_logic_vector(57, 8),
53831 => conv_std_logic_vector(58, 8),
53832 => conv_std_logic_vector(59, 8),
53833 => conv_std_logic_vector(59, 8),
53834 => conv_std_logic_vector(60, 8),
53835 => conv_std_logic_vector(61, 8),
53836 => conv_std_logic_vector(62, 8),
53837 => conv_std_logic_vector(63, 8),
53838 => conv_std_logic_vector(63, 8),
53839 => conv_std_logic_vector(64, 8),
53840 => conv_std_logic_vector(65, 8),
53841 => conv_std_logic_vector(66, 8),
53842 => conv_std_logic_vector(67, 8),
53843 => conv_std_logic_vector(68, 8),
53844 => conv_std_logic_vector(68, 8),
53845 => conv_std_logic_vector(69, 8),
53846 => conv_std_logic_vector(70, 8),
53847 => conv_std_logic_vector(71, 8),
53848 => conv_std_logic_vector(72, 8),
53849 => conv_std_logic_vector(73, 8),
53850 => conv_std_logic_vector(73, 8),
53851 => conv_std_logic_vector(74, 8),
53852 => conv_std_logic_vector(75, 8),
53853 => conv_std_logic_vector(76, 8),
53854 => conv_std_logic_vector(77, 8),
53855 => conv_std_logic_vector(77, 8),
53856 => conv_std_logic_vector(78, 8),
53857 => conv_std_logic_vector(79, 8),
53858 => conv_std_logic_vector(80, 8),
53859 => conv_std_logic_vector(81, 8),
53860 => conv_std_logic_vector(82, 8),
53861 => conv_std_logic_vector(82, 8),
53862 => conv_std_logic_vector(83, 8),
53863 => conv_std_logic_vector(84, 8),
53864 => conv_std_logic_vector(85, 8),
53865 => conv_std_logic_vector(86, 8),
53866 => conv_std_logic_vector(86, 8),
53867 => conv_std_logic_vector(87, 8),
53868 => conv_std_logic_vector(88, 8),
53869 => conv_std_logic_vector(89, 8),
53870 => conv_std_logic_vector(90, 8),
53871 => conv_std_logic_vector(91, 8),
53872 => conv_std_logic_vector(91, 8),
53873 => conv_std_logic_vector(92, 8),
53874 => conv_std_logic_vector(93, 8),
53875 => conv_std_logic_vector(94, 8),
53876 => conv_std_logic_vector(95, 8),
53877 => conv_std_logic_vector(95, 8),
53878 => conv_std_logic_vector(96, 8),
53879 => conv_std_logic_vector(97, 8),
53880 => conv_std_logic_vector(98, 8),
53881 => conv_std_logic_vector(99, 8),
53882 => conv_std_logic_vector(100, 8),
53883 => conv_std_logic_vector(100, 8),
53884 => conv_std_logic_vector(101, 8),
53885 => conv_std_logic_vector(102, 8),
53886 => conv_std_logic_vector(103, 8),
53887 => conv_std_logic_vector(104, 8),
53888 => conv_std_logic_vector(105, 8),
53889 => conv_std_logic_vector(105, 8),
53890 => conv_std_logic_vector(106, 8),
53891 => conv_std_logic_vector(107, 8),
53892 => conv_std_logic_vector(108, 8),
53893 => conv_std_logic_vector(109, 8),
53894 => conv_std_logic_vector(109, 8),
53895 => conv_std_logic_vector(110, 8),
53896 => conv_std_logic_vector(111, 8),
53897 => conv_std_logic_vector(112, 8),
53898 => conv_std_logic_vector(113, 8),
53899 => conv_std_logic_vector(114, 8),
53900 => conv_std_logic_vector(114, 8),
53901 => conv_std_logic_vector(115, 8),
53902 => conv_std_logic_vector(116, 8),
53903 => conv_std_logic_vector(117, 8),
53904 => conv_std_logic_vector(118, 8),
53905 => conv_std_logic_vector(118, 8),
53906 => conv_std_logic_vector(119, 8),
53907 => conv_std_logic_vector(120, 8),
53908 => conv_std_logic_vector(121, 8),
53909 => conv_std_logic_vector(122, 8),
53910 => conv_std_logic_vector(123, 8),
53911 => conv_std_logic_vector(123, 8),
53912 => conv_std_logic_vector(124, 8),
53913 => conv_std_logic_vector(125, 8),
53914 => conv_std_logic_vector(126, 8),
53915 => conv_std_logic_vector(127, 8),
53916 => conv_std_logic_vector(127, 8),
53917 => conv_std_logic_vector(128, 8),
53918 => conv_std_logic_vector(129, 8),
53919 => conv_std_logic_vector(130, 8),
53920 => conv_std_logic_vector(131, 8),
53921 => conv_std_logic_vector(132, 8),
53922 => conv_std_logic_vector(132, 8),
53923 => conv_std_logic_vector(133, 8),
53924 => conv_std_logic_vector(134, 8),
53925 => conv_std_logic_vector(135, 8),
53926 => conv_std_logic_vector(136, 8),
53927 => conv_std_logic_vector(136, 8),
53928 => conv_std_logic_vector(137, 8),
53929 => conv_std_logic_vector(138, 8),
53930 => conv_std_logic_vector(139, 8),
53931 => conv_std_logic_vector(140, 8),
53932 => conv_std_logic_vector(141, 8),
53933 => conv_std_logic_vector(141, 8),
53934 => conv_std_logic_vector(142, 8),
53935 => conv_std_logic_vector(143, 8),
53936 => conv_std_logic_vector(144, 8),
53937 => conv_std_logic_vector(145, 8),
53938 => conv_std_logic_vector(146, 8),
53939 => conv_std_logic_vector(146, 8),
53940 => conv_std_logic_vector(147, 8),
53941 => conv_std_logic_vector(148, 8),
53942 => conv_std_logic_vector(149, 8),
53943 => conv_std_logic_vector(150, 8),
53944 => conv_std_logic_vector(150, 8),
53945 => conv_std_logic_vector(151, 8),
53946 => conv_std_logic_vector(152, 8),
53947 => conv_std_logic_vector(153, 8),
53948 => conv_std_logic_vector(154, 8),
53949 => conv_std_logic_vector(155, 8),
53950 => conv_std_logic_vector(155, 8),
53951 => conv_std_logic_vector(156, 8),
53952 => conv_std_logic_vector(157, 8),
53953 => conv_std_logic_vector(158, 8),
53954 => conv_std_logic_vector(159, 8),
53955 => conv_std_logic_vector(159, 8),
53956 => conv_std_logic_vector(160, 8),
53957 => conv_std_logic_vector(161, 8),
53958 => conv_std_logic_vector(162, 8),
53959 => conv_std_logic_vector(163, 8),
53960 => conv_std_logic_vector(164, 8),
53961 => conv_std_logic_vector(164, 8),
53962 => conv_std_logic_vector(165, 8),
53963 => conv_std_logic_vector(166, 8),
53964 => conv_std_logic_vector(167, 8),
53965 => conv_std_logic_vector(168, 8),
53966 => conv_std_logic_vector(168, 8),
53967 => conv_std_logic_vector(169, 8),
53968 => conv_std_logic_vector(170, 8),
53969 => conv_std_logic_vector(171, 8),
53970 => conv_std_logic_vector(172, 8),
53971 => conv_std_logic_vector(173, 8),
53972 => conv_std_logic_vector(173, 8),
53973 => conv_std_logic_vector(174, 8),
53974 => conv_std_logic_vector(175, 8),
53975 => conv_std_logic_vector(176, 8),
53976 => conv_std_logic_vector(177, 8),
53977 => conv_std_logic_vector(178, 8),
53978 => conv_std_logic_vector(178, 8),
53979 => conv_std_logic_vector(179, 8),
53980 => conv_std_logic_vector(180, 8),
53981 => conv_std_logic_vector(181, 8),
53982 => conv_std_logic_vector(182, 8),
53983 => conv_std_logic_vector(182, 8),
53984 => conv_std_logic_vector(183, 8),
53985 => conv_std_logic_vector(184, 8),
53986 => conv_std_logic_vector(185, 8),
53987 => conv_std_logic_vector(186, 8),
53988 => conv_std_logic_vector(187, 8),
53989 => conv_std_logic_vector(187, 8),
53990 => conv_std_logic_vector(188, 8),
53991 => conv_std_logic_vector(189, 8),
53992 => conv_std_logic_vector(190, 8),
53993 => conv_std_logic_vector(191, 8),
53994 => conv_std_logic_vector(191, 8),
53995 => conv_std_logic_vector(192, 8),
53996 => conv_std_logic_vector(193, 8),
53997 => conv_std_logic_vector(194, 8),
53998 => conv_std_logic_vector(195, 8),
53999 => conv_std_logic_vector(196, 8),
54000 => conv_std_logic_vector(196, 8),
54001 => conv_std_logic_vector(197, 8),
54002 => conv_std_logic_vector(198, 8),
54003 => conv_std_logic_vector(199, 8),
54004 => conv_std_logic_vector(200, 8),
54005 => conv_std_logic_vector(200, 8),
54006 => conv_std_logic_vector(201, 8),
54007 => conv_std_logic_vector(202, 8),
54008 => conv_std_logic_vector(203, 8),
54009 => conv_std_logic_vector(204, 8),
54010 => conv_std_logic_vector(205, 8),
54011 => conv_std_logic_vector(205, 8),
54012 => conv_std_logic_vector(206, 8),
54013 => conv_std_logic_vector(207, 8),
54014 => conv_std_logic_vector(208, 8),
54015 => conv_std_logic_vector(209, 8),
54016 => conv_std_logic_vector(0, 8),
54017 => conv_std_logic_vector(0, 8),
54018 => conv_std_logic_vector(1, 8),
54019 => conv_std_logic_vector(2, 8),
54020 => conv_std_logic_vector(3, 8),
54021 => conv_std_logic_vector(4, 8),
54022 => conv_std_logic_vector(4, 8),
54023 => conv_std_logic_vector(5, 8),
54024 => conv_std_logic_vector(6, 8),
54025 => conv_std_logic_vector(7, 8),
54026 => conv_std_logic_vector(8, 8),
54027 => conv_std_logic_vector(9, 8),
54028 => conv_std_logic_vector(9, 8),
54029 => conv_std_logic_vector(10, 8),
54030 => conv_std_logic_vector(11, 8),
54031 => conv_std_logic_vector(12, 8),
54032 => conv_std_logic_vector(13, 8),
54033 => conv_std_logic_vector(14, 8),
54034 => conv_std_logic_vector(14, 8),
54035 => conv_std_logic_vector(15, 8),
54036 => conv_std_logic_vector(16, 8),
54037 => conv_std_logic_vector(17, 8),
54038 => conv_std_logic_vector(18, 8),
54039 => conv_std_logic_vector(18, 8),
54040 => conv_std_logic_vector(19, 8),
54041 => conv_std_logic_vector(20, 8),
54042 => conv_std_logic_vector(21, 8),
54043 => conv_std_logic_vector(22, 8),
54044 => conv_std_logic_vector(23, 8),
54045 => conv_std_logic_vector(23, 8),
54046 => conv_std_logic_vector(24, 8),
54047 => conv_std_logic_vector(25, 8),
54048 => conv_std_logic_vector(26, 8),
54049 => conv_std_logic_vector(27, 8),
54050 => conv_std_logic_vector(28, 8),
54051 => conv_std_logic_vector(28, 8),
54052 => conv_std_logic_vector(29, 8),
54053 => conv_std_logic_vector(30, 8),
54054 => conv_std_logic_vector(31, 8),
54055 => conv_std_logic_vector(32, 8),
54056 => conv_std_logic_vector(32, 8),
54057 => conv_std_logic_vector(33, 8),
54058 => conv_std_logic_vector(34, 8),
54059 => conv_std_logic_vector(35, 8),
54060 => conv_std_logic_vector(36, 8),
54061 => conv_std_logic_vector(37, 8),
54062 => conv_std_logic_vector(37, 8),
54063 => conv_std_logic_vector(38, 8),
54064 => conv_std_logic_vector(39, 8),
54065 => conv_std_logic_vector(40, 8),
54066 => conv_std_logic_vector(41, 8),
54067 => conv_std_logic_vector(42, 8),
54068 => conv_std_logic_vector(42, 8),
54069 => conv_std_logic_vector(43, 8),
54070 => conv_std_logic_vector(44, 8),
54071 => conv_std_logic_vector(45, 8),
54072 => conv_std_logic_vector(46, 8),
54073 => conv_std_logic_vector(46, 8),
54074 => conv_std_logic_vector(47, 8),
54075 => conv_std_logic_vector(48, 8),
54076 => conv_std_logic_vector(49, 8),
54077 => conv_std_logic_vector(50, 8),
54078 => conv_std_logic_vector(51, 8),
54079 => conv_std_logic_vector(51, 8),
54080 => conv_std_logic_vector(52, 8),
54081 => conv_std_logic_vector(53, 8),
54082 => conv_std_logic_vector(54, 8),
54083 => conv_std_logic_vector(55, 8),
54084 => conv_std_logic_vector(56, 8),
54085 => conv_std_logic_vector(56, 8),
54086 => conv_std_logic_vector(57, 8),
54087 => conv_std_logic_vector(58, 8),
54088 => conv_std_logic_vector(59, 8),
54089 => conv_std_logic_vector(60, 8),
54090 => conv_std_logic_vector(60, 8),
54091 => conv_std_logic_vector(61, 8),
54092 => conv_std_logic_vector(62, 8),
54093 => conv_std_logic_vector(63, 8),
54094 => conv_std_logic_vector(64, 8),
54095 => conv_std_logic_vector(65, 8),
54096 => conv_std_logic_vector(65, 8),
54097 => conv_std_logic_vector(66, 8),
54098 => conv_std_logic_vector(67, 8),
54099 => conv_std_logic_vector(68, 8),
54100 => conv_std_logic_vector(69, 8),
54101 => conv_std_logic_vector(70, 8),
54102 => conv_std_logic_vector(70, 8),
54103 => conv_std_logic_vector(71, 8),
54104 => conv_std_logic_vector(72, 8),
54105 => conv_std_logic_vector(73, 8),
54106 => conv_std_logic_vector(74, 8),
54107 => conv_std_logic_vector(75, 8),
54108 => conv_std_logic_vector(75, 8),
54109 => conv_std_logic_vector(76, 8),
54110 => conv_std_logic_vector(77, 8),
54111 => conv_std_logic_vector(78, 8),
54112 => conv_std_logic_vector(79, 8),
54113 => conv_std_logic_vector(79, 8),
54114 => conv_std_logic_vector(80, 8),
54115 => conv_std_logic_vector(81, 8),
54116 => conv_std_logic_vector(82, 8),
54117 => conv_std_logic_vector(83, 8),
54118 => conv_std_logic_vector(84, 8),
54119 => conv_std_logic_vector(84, 8),
54120 => conv_std_logic_vector(85, 8),
54121 => conv_std_logic_vector(86, 8),
54122 => conv_std_logic_vector(87, 8),
54123 => conv_std_logic_vector(88, 8),
54124 => conv_std_logic_vector(89, 8),
54125 => conv_std_logic_vector(89, 8),
54126 => conv_std_logic_vector(90, 8),
54127 => conv_std_logic_vector(91, 8),
54128 => conv_std_logic_vector(92, 8),
54129 => conv_std_logic_vector(93, 8),
54130 => conv_std_logic_vector(93, 8),
54131 => conv_std_logic_vector(94, 8),
54132 => conv_std_logic_vector(95, 8),
54133 => conv_std_logic_vector(96, 8),
54134 => conv_std_logic_vector(97, 8),
54135 => conv_std_logic_vector(98, 8),
54136 => conv_std_logic_vector(98, 8),
54137 => conv_std_logic_vector(99, 8),
54138 => conv_std_logic_vector(100, 8),
54139 => conv_std_logic_vector(101, 8),
54140 => conv_std_logic_vector(102, 8),
54141 => conv_std_logic_vector(103, 8),
54142 => conv_std_logic_vector(103, 8),
54143 => conv_std_logic_vector(104, 8),
54144 => conv_std_logic_vector(105, 8),
54145 => conv_std_logic_vector(106, 8),
54146 => conv_std_logic_vector(107, 8),
54147 => conv_std_logic_vector(107, 8),
54148 => conv_std_logic_vector(108, 8),
54149 => conv_std_logic_vector(109, 8),
54150 => conv_std_logic_vector(110, 8),
54151 => conv_std_logic_vector(111, 8),
54152 => conv_std_logic_vector(112, 8),
54153 => conv_std_logic_vector(112, 8),
54154 => conv_std_logic_vector(113, 8),
54155 => conv_std_logic_vector(114, 8),
54156 => conv_std_logic_vector(115, 8),
54157 => conv_std_logic_vector(116, 8),
54158 => conv_std_logic_vector(117, 8),
54159 => conv_std_logic_vector(117, 8),
54160 => conv_std_logic_vector(118, 8),
54161 => conv_std_logic_vector(119, 8),
54162 => conv_std_logic_vector(120, 8),
54163 => conv_std_logic_vector(121, 8),
54164 => conv_std_logic_vector(121, 8),
54165 => conv_std_logic_vector(122, 8),
54166 => conv_std_logic_vector(123, 8),
54167 => conv_std_logic_vector(124, 8),
54168 => conv_std_logic_vector(125, 8),
54169 => conv_std_logic_vector(126, 8),
54170 => conv_std_logic_vector(126, 8),
54171 => conv_std_logic_vector(127, 8),
54172 => conv_std_logic_vector(128, 8),
54173 => conv_std_logic_vector(129, 8),
54174 => conv_std_logic_vector(130, 8),
54175 => conv_std_logic_vector(131, 8),
54176 => conv_std_logic_vector(131, 8),
54177 => conv_std_logic_vector(132, 8),
54178 => conv_std_logic_vector(133, 8),
54179 => conv_std_logic_vector(134, 8),
54180 => conv_std_logic_vector(135, 8),
54181 => conv_std_logic_vector(135, 8),
54182 => conv_std_logic_vector(136, 8),
54183 => conv_std_logic_vector(137, 8),
54184 => conv_std_logic_vector(138, 8),
54185 => conv_std_logic_vector(139, 8),
54186 => conv_std_logic_vector(140, 8),
54187 => conv_std_logic_vector(140, 8),
54188 => conv_std_logic_vector(141, 8),
54189 => conv_std_logic_vector(142, 8),
54190 => conv_std_logic_vector(143, 8),
54191 => conv_std_logic_vector(144, 8),
54192 => conv_std_logic_vector(145, 8),
54193 => conv_std_logic_vector(145, 8),
54194 => conv_std_logic_vector(146, 8),
54195 => conv_std_logic_vector(147, 8),
54196 => conv_std_logic_vector(148, 8),
54197 => conv_std_logic_vector(149, 8),
54198 => conv_std_logic_vector(150, 8),
54199 => conv_std_logic_vector(150, 8),
54200 => conv_std_logic_vector(151, 8),
54201 => conv_std_logic_vector(152, 8),
54202 => conv_std_logic_vector(153, 8),
54203 => conv_std_logic_vector(154, 8),
54204 => conv_std_logic_vector(154, 8),
54205 => conv_std_logic_vector(155, 8),
54206 => conv_std_logic_vector(156, 8),
54207 => conv_std_logic_vector(157, 8),
54208 => conv_std_logic_vector(158, 8),
54209 => conv_std_logic_vector(159, 8),
54210 => conv_std_logic_vector(159, 8),
54211 => conv_std_logic_vector(160, 8),
54212 => conv_std_logic_vector(161, 8),
54213 => conv_std_logic_vector(162, 8),
54214 => conv_std_logic_vector(163, 8),
54215 => conv_std_logic_vector(164, 8),
54216 => conv_std_logic_vector(164, 8),
54217 => conv_std_logic_vector(165, 8),
54218 => conv_std_logic_vector(166, 8),
54219 => conv_std_logic_vector(167, 8),
54220 => conv_std_logic_vector(168, 8),
54221 => conv_std_logic_vector(168, 8),
54222 => conv_std_logic_vector(169, 8),
54223 => conv_std_logic_vector(170, 8),
54224 => conv_std_logic_vector(171, 8),
54225 => conv_std_logic_vector(172, 8),
54226 => conv_std_logic_vector(173, 8),
54227 => conv_std_logic_vector(173, 8),
54228 => conv_std_logic_vector(174, 8),
54229 => conv_std_logic_vector(175, 8),
54230 => conv_std_logic_vector(176, 8),
54231 => conv_std_logic_vector(177, 8),
54232 => conv_std_logic_vector(178, 8),
54233 => conv_std_logic_vector(178, 8),
54234 => conv_std_logic_vector(179, 8),
54235 => conv_std_logic_vector(180, 8),
54236 => conv_std_logic_vector(181, 8),
54237 => conv_std_logic_vector(182, 8),
54238 => conv_std_logic_vector(182, 8),
54239 => conv_std_logic_vector(183, 8),
54240 => conv_std_logic_vector(184, 8),
54241 => conv_std_logic_vector(185, 8),
54242 => conv_std_logic_vector(186, 8),
54243 => conv_std_logic_vector(187, 8),
54244 => conv_std_logic_vector(187, 8),
54245 => conv_std_logic_vector(188, 8),
54246 => conv_std_logic_vector(189, 8),
54247 => conv_std_logic_vector(190, 8),
54248 => conv_std_logic_vector(191, 8),
54249 => conv_std_logic_vector(192, 8),
54250 => conv_std_logic_vector(192, 8),
54251 => conv_std_logic_vector(193, 8),
54252 => conv_std_logic_vector(194, 8),
54253 => conv_std_logic_vector(195, 8),
54254 => conv_std_logic_vector(196, 8),
54255 => conv_std_logic_vector(196, 8),
54256 => conv_std_logic_vector(197, 8),
54257 => conv_std_logic_vector(198, 8),
54258 => conv_std_logic_vector(199, 8),
54259 => conv_std_logic_vector(200, 8),
54260 => conv_std_logic_vector(201, 8),
54261 => conv_std_logic_vector(201, 8),
54262 => conv_std_logic_vector(202, 8),
54263 => conv_std_logic_vector(203, 8),
54264 => conv_std_logic_vector(204, 8),
54265 => conv_std_logic_vector(205, 8),
54266 => conv_std_logic_vector(206, 8),
54267 => conv_std_logic_vector(206, 8),
54268 => conv_std_logic_vector(207, 8),
54269 => conv_std_logic_vector(208, 8),
54270 => conv_std_logic_vector(209, 8),
54271 => conv_std_logic_vector(210, 8),
54272 => conv_std_logic_vector(0, 8),
54273 => conv_std_logic_vector(0, 8),
54274 => conv_std_logic_vector(1, 8),
54275 => conv_std_logic_vector(2, 8),
54276 => conv_std_logic_vector(3, 8),
54277 => conv_std_logic_vector(4, 8),
54278 => conv_std_logic_vector(4, 8),
54279 => conv_std_logic_vector(5, 8),
54280 => conv_std_logic_vector(6, 8),
54281 => conv_std_logic_vector(7, 8),
54282 => conv_std_logic_vector(8, 8),
54283 => conv_std_logic_vector(9, 8),
54284 => conv_std_logic_vector(9, 8),
54285 => conv_std_logic_vector(10, 8),
54286 => conv_std_logic_vector(11, 8),
54287 => conv_std_logic_vector(12, 8),
54288 => conv_std_logic_vector(13, 8),
54289 => conv_std_logic_vector(14, 8),
54290 => conv_std_logic_vector(14, 8),
54291 => conv_std_logic_vector(15, 8),
54292 => conv_std_logic_vector(16, 8),
54293 => conv_std_logic_vector(17, 8),
54294 => conv_std_logic_vector(18, 8),
54295 => conv_std_logic_vector(19, 8),
54296 => conv_std_logic_vector(19, 8),
54297 => conv_std_logic_vector(20, 8),
54298 => conv_std_logic_vector(21, 8),
54299 => conv_std_logic_vector(22, 8),
54300 => conv_std_logic_vector(23, 8),
54301 => conv_std_logic_vector(24, 8),
54302 => conv_std_logic_vector(24, 8),
54303 => conv_std_logic_vector(25, 8),
54304 => conv_std_logic_vector(26, 8),
54305 => conv_std_logic_vector(27, 8),
54306 => conv_std_logic_vector(28, 8),
54307 => conv_std_logic_vector(28, 8),
54308 => conv_std_logic_vector(29, 8),
54309 => conv_std_logic_vector(30, 8),
54310 => conv_std_logic_vector(31, 8),
54311 => conv_std_logic_vector(32, 8),
54312 => conv_std_logic_vector(33, 8),
54313 => conv_std_logic_vector(33, 8),
54314 => conv_std_logic_vector(34, 8),
54315 => conv_std_logic_vector(35, 8),
54316 => conv_std_logic_vector(36, 8),
54317 => conv_std_logic_vector(37, 8),
54318 => conv_std_logic_vector(38, 8),
54319 => conv_std_logic_vector(38, 8),
54320 => conv_std_logic_vector(39, 8),
54321 => conv_std_logic_vector(40, 8),
54322 => conv_std_logic_vector(41, 8),
54323 => conv_std_logic_vector(42, 8),
54324 => conv_std_logic_vector(43, 8),
54325 => conv_std_logic_vector(43, 8),
54326 => conv_std_logic_vector(44, 8),
54327 => conv_std_logic_vector(45, 8),
54328 => conv_std_logic_vector(46, 8),
54329 => conv_std_logic_vector(47, 8),
54330 => conv_std_logic_vector(48, 8),
54331 => conv_std_logic_vector(48, 8),
54332 => conv_std_logic_vector(49, 8),
54333 => conv_std_logic_vector(50, 8),
54334 => conv_std_logic_vector(51, 8),
54335 => conv_std_logic_vector(52, 8),
54336 => conv_std_logic_vector(53, 8),
54337 => conv_std_logic_vector(53, 8),
54338 => conv_std_logic_vector(54, 8),
54339 => conv_std_logic_vector(55, 8),
54340 => conv_std_logic_vector(56, 8),
54341 => conv_std_logic_vector(57, 8),
54342 => conv_std_logic_vector(57, 8),
54343 => conv_std_logic_vector(58, 8),
54344 => conv_std_logic_vector(59, 8),
54345 => conv_std_logic_vector(60, 8),
54346 => conv_std_logic_vector(61, 8),
54347 => conv_std_logic_vector(62, 8),
54348 => conv_std_logic_vector(62, 8),
54349 => conv_std_logic_vector(63, 8),
54350 => conv_std_logic_vector(64, 8),
54351 => conv_std_logic_vector(65, 8),
54352 => conv_std_logic_vector(66, 8),
54353 => conv_std_logic_vector(67, 8),
54354 => conv_std_logic_vector(67, 8),
54355 => conv_std_logic_vector(68, 8),
54356 => conv_std_logic_vector(69, 8),
54357 => conv_std_logic_vector(70, 8),
54358 => conv_std_logic_vector(71, 8),
54359 => conv_std_logic_vector(72, 8),
54360 => conv_std_logic_vector(72, 8),
54361 => conv_std_logic_vector(73, 8),
54362 => conv_std_logic_vector(74, 8),
54363 => conv_std_logic_vector(75, 8),
54364 => conv_std_logic_vector(76, 8),
54365 => conv_std_logic_vector(77, 8),
54366 => conv_std_logic_vector(77, 8),
54367 => conv_std_logic_vector(78, 8),
54368 => conv_std_logic_vector(79, 8),
54369 => conv_std_logic_vector(80, 8),
54370 => conv_std_logic_vector(81, 8),
54371 => conv_std_logic_vector(81, 8),
54372 => conv_std_logic_vector(82, 8),
54373 => conv_std_logic_vector(83, 8),
54374 => conv_std_logic_vector(84, 8),
54375 => conv_std_logic_vector(85, 8),
54376 => conv_std_logic_vector(86, 8),
54377 => conv_std_logic_vector(86, 8),
54378 => conv_std_logic_vector(87, 8),
54379 => conv_std_logic_vector(88, 8),
54380 => conv_std_logic_vector(89, 8),
54381 => conv_std_logic_vector(90, 8),
54382 => conv_std_logic_vector(91, 8),
54383 => conv_std_logic_vector(91, 8),
54384 => conv_std_logic_vector(92, 8),
54385 => conv_std_logic_vector(93, 8),
54386 => conv_std_logic_vector(94, 8),
54387 => conv_std_logic_vector(95, 8),
54388 => conv_std_logic_vector(96, 8),
54389 => conv_std_logic_vector(96, 8),
54390 => conv_std_logic_vector(97, 8),
54391 => conv_std_logic_vector(98, 8),
54392 => conv_std_logic_vector(99, 8),
54393 => conv_std_logic_vector(100, 8),
54394 => conv_std_logic_vector(101, 8),
54395 => conv_std_logic_vector(101, 8),
54396 => conv_std_logic_vector(102, 8),
54397 => conv_std_logic_vector(103, 8),
54398 => conv_std_logic_vector(104, 8),
54399 => conv_std_logic_vector(105, 8),
54400 => conv_std_logic_vector(106, 8),
54401 => conv_std_logic_vector(106, 8),
54402 => conv_std_logic_vector(107, 8),
54403 => conv_std_logic_vector(108, 8),
54404 => conv_std_logic_vector(109, 8),
54405 => conv_std_logic_vector(110, 8),
54406 => conv_std_logic_vector(110, 8),
54407 => conv_std_logic_vector(111, 8),
54408 => conv_std_logic_vector(112, 8),
54409 => conv_std_logic_vector(113, 8),
54410 => conv_std_logic_vector(114, 8),
54411 => conv_std_logic_vector(115, 8),
54412 => conv_std_logic_vector(115, 8),
54413 => conv_std_logic_vector(116, 8),
54414 => conv_std_logic_vector(117, 8),
54415 => conv_std_logic_vector(118, 8),
54416 => conv_std_logic_vector(119, 8),
54417 => conv_std_logic_vector(120, 8),
54418 => conv_std_logic_vector(120, 8),
54419 => conv_std_logic_vector(121, 8),
54420 => conv_std_logic_vector(122, 8),
54421 => conv_std_logic_vector(123, 8),
54422 => conv_std_logic_vector(124, 8),
54423 => conv_std_logic_vector(125, 8),
54424 => conv_std_logic_vector(125, 8),
54425 => conv_std_logic_vector(126, 8),
54426 => conv_std_logic_vector(127, 8),
54427 => conv_std_logic_vector(128, 8),
54428 => conv_std_logic_vector(129, 8),
54429 => conv_std_logic_vector(130, 8),
54430 => conv_std_logic_vector(130, 8),
54431 => conv_std_logic_vector(131, 8),
54432 => conv_std_logic_vector(132, 8),
54433 => conv_std_logic_vector(133, 8),
54434 => conv_std_logic_vector(134, 8),
54435 => conv_std_logic_vector(134, 8),
54436 => conv_std_logic_vector(135, 8),
54437 => conv_std_logic_vector(136, 8),
54438 => conv_std_logic_vector(137, 8),
54439 => conv_std_logic_vector(138, 8),
54440 => conv_std_logic_vector(139, 8),
54441 => conv_std_logic_vector(139, 8),
54442 => conv_std_logic_vector(140, 8),
54443 => conv_std_logic_vector(141, 8),
54444 => conv_std_logic_vector(142, 8),
54445 => conv_std_logic_vector(143, 8),
54446 => conv_std_logic_vector(144, 8),
54447 => conv_std_logic_vector(144, 8),
54448 => conv_std_logic_vector(145, 8),
54449 => conv_std_logic_vector(146, 8),
54450 => conv_std_logic_vector(147, 8),
54451 => conv_std_logic_vector(148, 8),
54452 => conv_std_logic_vector(149, 8),
54453 => conv_std_logic_vector(149, 8),
54454 => conv_std_logic_vector(150, 8),
54455 => conv_std_logic_vector(151, 8),
54456 => conv_std_logic_vector(152, 8),
54457 => conv_std_logic_vector(153, 8),
54458 => conv_std_logic_vector(154, 8),
54459 => conv_std_logic_vector(154, 8),
54460 => conv_std_logic_vector(155, 8),
54461 => conv_std_logic_vector(156, 8),
54462 => conv_std_logic_vector(157, 8),
54463 => conv_std_logic_vector(158, 8),
54464 => conv_std_logic_vector(159, 8),
54465 => conv_std_logic_vector(159, 8),
54466 => conv_std_logic_vector(160, 8),
54467 => conv_std_logic_vector(161, 8),
54468 => conv_std_logic_vector(162, 8),
54469 => conv_std_logic_vector(163, 8),
54470 => conv_std_logic_vector(163, 8),
54471 => conv_std_logic_vector(164, 8),
54472 => conv_std_logic_vector(165, 8),
54473 => conv_std_logic_vector(166, 8),
54474 => conv_std_logic_vector(167, 8),
54475 => conv_std_logic_vector(168, 8),
54476 => conv_std_logic_vector(168, 8),
54477 => conv_std_logic_vector(169, 8),
54478 => conv_std_logic_vector(170, 8),
54479 => conv_std_logic_vector(171, 8),
54480 => conv_std_logic_vector(172, 8),
54481 => conv_std_logic_vector(173, 8),
54482 => conv_std_logic_vector(173, 8),
54483 => conv_std_logic_vector(174, 8),
54484 => conv_std_logic_vector(175, 8),
54485 => conv_std_logic_vector(176, 8),
54486 => conv_std_logic_vector(177, 8),
54487 => conv_std_logic_vector(178, 8),
54488 => conv_std_logic_vector(178, 8),
54489 => conv_std_logic_vector(179, 8),
54490 => conv_std_logic_vector(180, 8),
54491 => conv_std_logic_vector(181, 8),
54492 => conv_std_logic_vector(182, 8),
54493 => conv_std_logic_vector(183, 8),
54494 => conv_std_logic_vector(183, 8),
54495 => conv_std_logic_vector(184, 8),
54496 => conv_std_logic_vector(185, 8),
54497 => conv_std_logic_vector(186, 8),
54498 => conv_std_logic_vector(187, 8),
54499 => conv_std_logic_vector(187, 8),
54500 => conv_std_logic_vector(188, 8),
54501 => conv_std_logic_vector(189, 8),
54502 => conv_std_logic_vector(190, 8),
54503 => conv_std_logic_vector(191, 8),
54504 => conv_std_logic_vector(192, 8),
54505 => conv_std_logic_vector(192, 8),
54506 => conv_std_logic_vector(193, 8),
54507 => conv_std_logic_vector(194, 8),
54508 => conv_std_logic_vector(195, 8),
54509 => conv_std_logic_vector(196, 8),
54510 => conv_std_logic_vector(197, 8),
54511 => conv_std_logic_vector(197, 8),
54512 => conv_std_logic_vector(198, 8),
54513 => conv_std_logic_vector(199, 8),
54514 => conv_std_logic_vector(200, 8),
54515 => conv_std_logic_vector(201, 8),
54516 => conv_std_logic_vector(202, 8),
54517 => conv_std_logic_vector(202, 8),
54518 => conv_std_logic_vector(203, 8),
54519 => conv_std_logic_vector(204, 8),
54520 => conv_std_logic_vector(205, 8),
54521 => conv_std_logic_vector(206, 8),
54522 => conv_std_logic_vector(207, 8),
54523 => conv_std_logic_vector(207, 8),
54524 => conv_std_logic_vector(208, 8),
54525 => conv_std_logic_vector(209, 8),
54526 => conv_std_logic_vector(210, 8),
54527 => conv_std_logic_vector(211, 8),
54528 => conv_std_logic_vector(0, 8),
54529 => conv_std_logic_vector(0, 8),
54530 => conv_std_logic_vector(1, 8),
54531 => conv_std_logic_vector(2, 8),
54532 => conv_std_logic_vector(3, 8),
54533 => conv_std_logic_vector(4, 8),
54534 => conv_std_logic_vector(4, 8),
54535 => conv_std_logic_vector(5, 8),
54536 => conv_std_logic_vector(6, 8),
54537 => conv_std_logic_vector(7, 8),
54538 => conv_std_logic_vector(8, 8),
54539 => conv_std_logic_vector(9, 8),
54540 => conv_std_logic_vector(9, 8),
54541 => conv_std_logic_vector(10, 8),
54542 => conv_std_logic_vector(11, 8),
54543 => conv_std_logic_vector(12, 8),
54544 => conv_std_logic_vector(13, 8),
54545 => conv_std_logic_vector(14, 8),
54546 => conv_std_logic_vector(14, 8),
54547 => conv_std_logic_vector(15, 8),
54548 => conv_std_logic_vector(16, 8),
54549 => conv_std_logic_vector(17, 8),
54550 => conv_std_logic_vector(18, 8),
54551 => conv_std_logic_vector(19, 8),
54552 => conv_std_logic_vector(19, 8),
54553 => conv_std_logic_vector(20, 8),
54554 => conv_std_logic_vector(21, 8),
54555 => conv_std_logic_vector(22, 8),
54556 => conv_std_logic_vector(23, 8),
54557 => conv_std_logic_vector(24, 8),
54558 => conv_std_logic_vector(24, 8),
54559 => conv_std_logic_vector(25, 8),
54560 => conv_std_logic_vector(26, 8),
54561 => conv_std_logic_vector(27, 8),
54562 => conv_std_logic_vector(28, 8),
54563 => conv_std_logic_vector(29, 8),
54564 => conv_std_logic_vector(29, 8),
54565 => conv_std_logic_vector(30, 8),
54566 => conv_std_logic_vector(31, 8),
54567 => conv_std_logic_vector(32, 8),
54568 => conv_std_logic_vector(33, 8),
54569 => conv_std_logic_vector(34, 8),
54570 => conv_std_logic_vector(34, 8),
54571 => conv_std_logic_vector(35, 8),
54572 => conv_std_logic_vector(36, 8),
54573 => conv_std_logic_vector(37, 8),
54574 => conv_std_logic_vector(38, 8),
54575 => conv_std_logic_vector(39, 8),
54576 => conv_std_logic_vector(39, 8),
54577 => conv_std_logic_vector(40, 8),
54578 => conv_std_logic_vector(41, 8),
54579 => conv_std_logic_vector(42, 8),
54580 => conv_std_logic_vector(43, 8),
54581 => conv_std_logic_vector(44, 8),
54582 => conv_std_logic_vector(44, 8),
54583 => conv_std_logic_vector(45, 8),
54584 => conv_std_logic_vector(46, 8),
54585 => conv_std_logic_vector(47, 8),
54586 => conv_std_logic_vector(48, 8),
54587 => conv_std_logic_vector(49, 8),
54588 => conv_std_logic_vector(49, 8),
54589 => conv_std_logic_vector(50, 8),
54590 => conv_std_logic_vector(51, 8),
54591 => conv_std_logic_vector(52, 8),
54592 => conv_std_logic_vector(53, 8),
54593 => conv_std_logic_vector(54, 8),
54594 => conv_std_logic_vector(54, 8),
54595 => conv_std_logic_vector(55, 8),
54596 => conv_std_logic_vector(56, 8),
54597 => conv_std_logic_vector(57, 8),
54598 => conv_std_logic_vector(58, 8),
54599 => conv_std_logic_vector(59, 8),
54600 => conv_std_logic_vector(59, 8),
54601 => conv_std_logic_vector(60, 8),
54602 => conv_std_logic_vector(61, 8),
54603 => conv_std_logic_vector(62, 8),
54604 => conv_std_logic_vector(63, 8),
54605 => conv_std_logic_vector(64, 8),
54606 => conv_std_logic_vector(64, 8),
54607 => conv_std_logic_vector(65, 8),
54608 => conv_std_logic_vector(66, 8),
54609 => conv_std_logic_vector(67, 8),
54610 => conv_std_logic_vector(68, 8),
54611 => conv_std_logic_vector(69, 8),
54612 => conv_std_logic_vector(69, 8),
54613 => conv_std_logic_vector(70, 8),
54614 => conv_std_logic_vector(71, 8),
54615 => conv_std_logic_vector(72, 8),
54616 => conv_std_logic_vector(73, 8),
54617 => conv_std_logic_vector(74, 8),
54618 => conv_std_logic_vector(74, 8),
54619 => conv_std_logic_vector(75, 8),
54620 => conv_std_logic_vector(76, 8),
54621 => conv_std_logic_vector(77, 8),
54622 => conv_std_logic_vector(78, 8),
54623 => conv_std_logic_vector(79, 8),
54624 => conv_std_logic_vector(79, 8),
54625 => conv_std_logic_vector(80, 8),
54626 => conv_std_logic_vector(81, 8),
54627 => conv_std_logic_vector(82, 8),
54628 => conv_std_logic_vector(83, 8),
54629 => conv_std_logic_vector(84, 8),
54630 => conv_std_logic_vector(84, 8),
54631 => conv_std_logic_vector(85, 8),
54632 => conv_std_logic_vector(86, 8),
54633 => conv_std_logic_vector(87, 8),
54634 => conv_std_logic_vector(88, 8),
54635 => conv_std_logic_vector(89, 8),
54636 => conv_std_logic_vector(89, 8),
54637 => conv_std_logic_vector(90, 8),
54638 => conv_std_logic_vector(91, 8),
54639 => conv_std_logic_vector(92, 8),
54640 => conv_std_logic_vector(93, 8),
54641 => conv_std_logic_vector(94, 8),
54642 => conv_std_logic_vector(94, 8),
54643 => conv_std_logic_vector(95, 8),
54644 => conv_std_logic_vector(96, 8),
54645 => conv_std_logic_vector(97, 8),
54646 => conv_std_logic_vector(98, 8),
54647 => conv_std_logic_vector(99, 8),
54648 => conv_std_logic_vector(99, 8),
54649 => conv_std_logic_vector(100, 8),
54650 => conv_std_logic_vector(101, 8),
54651 => conv_std_logic_vector(102, 8),
54652 => conv_std_logic_vector(103, 8),
54653 => conv_std_logic_vector(104, 8),
54654 => conv_std_logic_vector(104, 8),
54655 => conv_std_logic_vector(105, 8),
54656 => conv_std_logic_vector(106, 8),
54657 => conv_std_logic_vector(107, 8),
54658 => conv_std_logic_vector(108, 8),
54659 => conv_std_logic_vector(108, 8),
54660 => conv_std_logic_vector(109, 8),
54661 => conv_std_logic_vector(110, 8),
54662 => conv_std_logic_vector(111, 8),
54663 => conv_std_logic_vector(112, 8),
54664 => conv_std_logic_vector(113, 8),
54665 => conv_std_logic_vector(113, 8),
54666 => conv_std_logic_vector(114, 8),
54667 => conv_std_logic_vector(115, 8),
54668 => conv_std_logic_vector(116, 8),
54669 => conv_std_logic_vector(117, 8),
54670 => conv_std_logic_vector(118, 8),
54671 => conv_std_logic_vector(118, 8),
54672 => conv_std_logic_vector(119, 8),
54673 => conv_std_logic_vector(120, 8),
54674 => conv_std_logic_vector(121, 8),
54675 => conv_std_logic_vector(122, 8),
54676 => conv_std_logic_vector(123, 8),
54677 => conv_std_logic_vector(123, 8),
54678 => conv_std_logic_vector(124, 8),
54679 => conv_std_logic_vector(125, 8),
54680 => conv_std_logic_vector(126, 8),
54681 => conv_std_logic_vector(127, 8),
54682 => conv_std_logic_vector(128, 8),
54683 => conv_std_logic_vector(128, 8),
54684 => conv_std_logic_vector(129, 8),
54685 => conv_std_logic_vector(130, 8),
54686 => conv_std_logic_vector(131, 8),
54687 => conv_std_logic_vector(132, 8),
54688 => conv_std_logic_vector(133, 8),
54689 => conv_std_logic_vector(133, 8),
54690 => conv_std_logic_vector(134, 8),
54691 => conv_std_logic_vector(135, 8),
54692 => conv_std_logic_vector(136, 8),
54693 => conv_std_logic_vector(137, 8),
54694 => conv_std_logic_vector(138, 8),
54695 => conv_std_logic_vector(138, 8),
54696 => conv_std_logic_vector(139, 8),
54697 => conv_std_logic_vector(140, 8),
54698 => conv_std_logic_vector(141, 8),
54699 => conv_std_logic_vector(142, 8),
54700 => conv_std_logic_vector(143, 8),
54701 => conv_std_logic_vector(143, 8),
54702 => conv_std_logic_vector(144, 8),
54703 => conv_std_logic_vector(145, 8),
54704 => conv_std_logic_vector(146, 8),
54705 => conv_std_logic_vector(147, 8),
54706 => conv_std_logic_vector(148, 8),
54707 => conv_std_logic_vector(148, 8),
54708 => conv_std_logic_vector(149, 8),
54709 => conv_std_logic_vector(150, 8),
54710 => conv_std_logic_vector(151, 8),
54711 => conv_std_logic_vector(152, 8),
54712 => conv_std_logic_vector(153, 8),
54713 => conv_std_logic_vector(153, 8),
54714 => conv_std_logic_vector(154, 8),
54715 => conv_std_logic_vector(155, 8),
54716 => conv_std_logic_vector(156, 8),
54717 => conv_std_logic_vector(157, 8),
54718 => conv_std_logic_vector(158, 8),
54719 => conv_std_logic_vector(158, 8),
54720 => conv_std_logic_vector(159, 8),
54721 => conv_std_logic_vector(160, 8),
54722 => conv_std_logic_vector(161, 8),
54723 => conv_std_logic_vector(162, 8),
54724 => conv_std_logic_vector(163, 8),
54725 => conv_std_logic_vector(163, 8),
54726 => conv_std_logic_vector(164, 8),
54727 => conv_std_logic_vector(165, 8),
54728 => conv_std_logic_vector(166, 8),
54729 => conv_std_logic_vector(167, 8),
54730 => conv_std_logic_vector(168, 8),
54731 => conv_std_logic_vector(168, 8),
54732 => conv_std_logic_vector(169, 8),
54733 => conv_std_logic_vector(170, 8),
54734 => conv_std_logic_vector(171, 8),
54735 => conv_std_logic_vector(172, 8),
54736 => conv_std_logic_vector(173, 8),
54737 => conv_std_logic_vector(173, 8),
54738 => conv_std_logic_vector(174, 8),
54739 => conv_std_logic_vector(175, 8),
54740 => conv_std_logic_vector(176, 8),
54741 => conv_std_logic_vector(177, 8),
54742 => conv_std_logic_vector(178, 8),
54743 => conv_std_logic_vector(178, 8),
54744 => conv_std_logic_vector(179, 8),
54745 => conv_std_logic_vector(180, 8),
54746 => conv_std_logic_vector(181, 8),
54747 => conv_std_logic_vector(182, 8),
54748 => conv_std_logic_vector(183, 8),
54749 => conv_std_logic_vector(183, 8),
54750 => conv_std_logic_vector(184, 8),
54751 => conv_std_logic_vector(185, 8),
54752 => conv_std_logic_vector(186, 8),
54753 => conv_std_logic_vector(187, 8),
54754 => conv_std_logic_vector(188, 8),
54755 => conv_std_logic_vector(188, 8),
54756 => conv_std_logic_vector(189, 8),
54757 => conv_std_logic_vector(190, 8),
54758 => conv_std_logic_vector(191, 8),
54759 => conv_std_logic_vector(192, 8),
54760 => conv_std_logic_vector(193, 8),
54761 => conv_std_logic_vector(193, 8),
54762 => conv_std_logic_vector(194, 8),
54763 => conv_std_logic_vector(195, 8),
54764 => conv_std_logic_vector(196, 8),
54765 => conv_std_logic_vector(197, 8),
54766 => conv_std_logic_vector(198, 8),
54767 => conv_std_logic_vector(198, 8),
54768 => conv_std_logic_vector(199, 8),
54769 => conv_std_logic_vector(200, 8),
54770 => conv_std_logic_vector(201, 8),
54771 => conv_std_logic_vector(202, 8),
54772 => conv_std_logic_vector(203, 8),
54773 => conv_std_logic_vector(203, 8),
54774 => conv_std_logic_vector(204, 8),
54775 => conv_std_logic_vector(205, 8),
54776 => conv_std_logic_vector(206, 8),
54777 => conv_std_logic_vector(207, 8),
54778 => conv_std_logic_vector(208, 8),
54779 => conv_std_logic_vector(208, 8),
54780 => conv_std_logic_vector(209, 8),
54781 => conv_std_logic_vector(210, 8),
54782 => conv_std_logic_vector(211, 8),
54783 => conv_std_logic_vector(212, 8),
54784 => conv_std_logic_vector(0, 8),
54785 => conv_std_logic_vector(0, 8),
54786 => conv_std_logic_vector(1, 8),
54787 => conv_std_logic_vector(2, 8),
54788 => conv_std_logic_vector(3, 8),
54789 => conv_std_logic_vector(4, 8),
54790 => conv_std_logic_vector(5, 8),
54791 => conv_std_logic_vector(5, 8),
54792 => conv_std_logic_vector(6, 8),
54793 => conv_std_logic_vector(7, 8),
54794 => conv_std_logic_vector(8, 8),
54795 => conv_std_logic_vector(9, 8),
54796 => conv_std_logic_vector(10, 8),
54797 => conv_std_logic_vector(10, 8),
54798 => conv_std_logic_vector(11, 8),
54799 => conv_std_logic_vector(12, 8),
54800 => conv_std_logic_vector(13, 8),
54801 => conv_std_logic_vector(14, 8),
54802 => conv_std_logic_vector(15, 8),
54803 => conv_std_logic_vector(15, 8),
54804 => conv_std_logic_vector(16, 8),
54805 => conv_std_logic_vector(17, 8),
54806 => conv_std_logic_vector(18, 8),
54807 => conv_std_logic_vector(19, 8),
54808 => conv_std_logic_vector(20, 8),
54809 => conv_std_logic_vector(20, 8),
54810 => conv_std_logic_vector(21, 8),
54811 => conv_std_logic_vector(22, 8),
54812 => conv_std_logic_vector(23, 8),
54813 => conv_std_logic_vector(24, 8),
54814 => conv_std_logic_vector(25, 8),
54815 => conv_std_logic_vector(25, 8),
54816 => conv_std_logic_vector(26, 8),
54817 => conv_std_logic_vector(27, 8),
54818 => conv_std_logic_vector(28, 8),
54819 => conv_std_logic_vector(29, 8),
54820 => conv_std_logic_vector(30, 8),
54821 => conv_std_logic_vector(30, 8),
54822 => conv_std_logic_vector(31, 8),
54823 => conv_std_logic_vector(32, 8),
54824 => conv_std_logic_vector(33, 8),
54825 => conv_std_logic_vector(34, 8),
54826 => conv_std_logic_vector(35, 8),
54827 => conv_std_logic_vector(35, 8),
54828 => conv_std_logic_vector(36, 8),
54829 => conv_std_logic_vector(37, 8),
54830 => conv_std_logic_vector(38, 8),
54831 => conv_std_logic_vector(39, 8),
54832 => conv_std_logic_vector(40, 8),
54833 => conv_std_logic_vector(40, 8),
54834 => conv_std_logic_vector(41, 8),
54835 => conv_std_logic_vector(42, 8),
54836 => conv_std_logic_vector(43, 8),
54837 => conv_std_logic_vector(44, 8),
54838 => conv_std_logic_vector(45, 8),
54839 => conv_std_logic_vector(45, 8),
54840 => conv_std_logic_vector(46, 8),
54841 => conv_std_logic_vector(47, 8),
54842 => conv_std_logic_vector(48, 8),
54843 => conv_std_logic_vector(49, 8),
54844 => conv_std_logic_vector(50, 8),
54845 => conv_std_logic_vector(50, 8),
54846 => conv_std_logic_vector(51, 8),
54847 => conv_std_logic_vector(52, 8),
54848 => conv_std_logic_vector(53, 8),
54849 => conv_std_logic_vector(54, 8),
54850 => conv_std_logic_vector(55, 8),
54851 => conv_std_logic_vector(56, 8),
54852 => conv_std_logic_vector(56, 8),
54853 => conv_std_logic_vector(57, 8),
54854 => conv_std_logic_vector(58, 8),
54855 => conv_std_logic_vector(59, 8),
54856 => conv_std_logic_vector(60, 8),
54857 => conv_std_logic_vector(61, 8),
54858 => conv_std_logic_vector(61, 8),
54859 => conv_std_logic_vector(62, 8),
54860 => conv_std_logic_vector(63, 8),
54861 => conv_std_logic_vector(64, 8),
54862 => conv_std_logic_vector(65, 8),
54863 => conv_std_logic_vector(66, 8),
54864 => conv_std_logic_vector(66, 8),
54865 => conv_std_logic_vector(67, 8),
54866 => conv_std_logic_vector(68, 8),
54867 => conv_std_logic_vector(69, 8),
54868 => conv_std_logic_vector(70, 8),
54869 => conv_std_logic_vector(71, 8),
54870 => conv_std_logic_vector(71, 8),
54871 => conv_std_logic_vector(72, 8),
54872 => conv_std_logic_vector(73, 8),
54873 => conv_std_logic_vector(74, 8),
54874 => conv_std_logic_vector(75, 8),
54875 => conv_std_logic_vector(76, 8),
54876 => conv_std_logic_vector(76, 8),
54877 => conv_std_logic_vector(77, 8),
54878 => conv_std_logic_vector(78, 8),
54879 => conv_std_logic_vector(79, 8),
54880 => conv_std_logic_vector(80, 8),
54881 => conv_std_logic_vector(81, 8),
54882 => conv_std_logic_vector(81, 8),
54883 => conv_std_logic_vector(82, 8),
54884 => conv_std_logic_vector(83, 8),
54885 => conv_std_logic_vector(84, 8),
54886 => conv_std_logic_vector(85, 8),
54887 => conv_std_logic_vector(86, 8),
54888 => conv_std_logic_vector(86, 8),
54889 => conv_std_logic_vector(87, 8),
54890 => conv_std_logic_vector(88, 8),
54891 => conv_std_logic_vector(89, 8),
54892 => conv_std_logic_vector(90, 8),
54893 => conv_std_logic_vector(91, 8),
54894 => conv_std_logic_vector(91, 8),
54895 => conv_std_logic_vector(92, 8),
54896 => conv_std_logic_vector(93, 8),
54897 => conv_std_logic_vector(94, 8),
54898 => conv_std_logic_vector(95, 8),
54899 => conv_std_logic_vector(96, 8),
54900 => conv_std_logic_vector(96, 8),
54901 => conv_std_logic_vector(97, 8),
54902 => conv_std_logic_vector(98, 8),
54903 => conv_std_logic_vector(99, 8),
54904 => conv_std_logic_vector(100, 8),
54905 => conv_std_logic_vector(101, 8),
54906 => conv_std_logic_vector(101, 8),
54907 => conv_std_logic_vector(102, 8),
54908 => conv_std_logic_vector(103, 8),
54909 => conv_std_logic_vector(104, 8),
54910 => conv_std_logic_vector(105, 8),
54911 => conv_std_logic_vector(106, 8),
54912 => conv_std_logic_vector(107, 8),
54913 => conv_std_logic_vector(107, 8),
54914 => conv_std_logic_vector(108, 8),
54915 => conv_std_logic_vector(109, 8),
54916 => conv_std_logic_vector(110, 8),
54917 => conv_std_logic_vector(111, 8),
54918 => conv_std_logic_vector(112, 8),
54919 => conv_std_logic_vector(112, 8),
54920 => conv_std_logic_vector(113, 8),
54921 => conv_std_logic_vector(114, 8),
54922 => conv_std_logic_vector(115, 8),
54923 => conv_std_logic_vector(116, 8),
54924 => conv_std_logic_vector(117, 8),
54925 => conv_std_logic_vector(117, 8),
54926 => conv_std_logic_vector(118, 8),
54927 => conv_std_logic_vector(119, 8),
54928 => conv_std_logic_vector(120, 8),
54929 => conv_std_logic_vector(121, 8),
54930 => conv_std_logic_vector(122, 8),
54931 => conv_std_logic_vector(122, 8),
54932 => conv_std_logic_vector(123, 8),
54933 => conv_std_logic_vector(124, 8),
54934 => conv_std_logic_vector(125, 8),
54935 => conv_std_logic_vector(126, 8),
54936 => conv_std_logic_vector(127, 8),
54937 => conv_std_logic_vector(127, 8),
54938 => conv_std_logic_vector(128, 8),
54939 => conv_std_logic_vector(129, 8),
54940 => conv_std_logic_vector(130, 8),
54941 => conv_std_logic_vector(131, 8),
54942 => conv_std_logic_vector(132, 8),
54943 => conv_std_logic_vector(132, 8),
54944 => conv_std_logic_vector(133, 8),
54945 => conv_std_logic_vector(134, 8),
54946 => conv_std_logic_vector(135, 8),
54947 => conv_std_logic_vector(136, 8),
54948 => conv_std_logic_vector(137, 8),
54949 => conv_std_logic_vector(137, 8),
54950 => conv_std_logic_vector(138, 8),
54951 => conv_std_logic_vector(139, 8),
54952 => conv_std_logic_vector(140, 8),
54953 => conv_std_logic_vector(141, 8),
54954 => conv_std_logic_vector(142, 8),
54955 => conv_std_logic_vector(142, 8),
54956 => conv_std_logic_vector(143, 8),
54957 => conv_std_logic_vector(144, 8),
54958 => conv_std_logic_vector(145, 8),
54959 => conv_std_logic_vector(146, 8),
54960 => conv_std_logic_vector(147, 8),
54961 => conv_std_logic_vector(147, 8),
54962 => conv_std_logic_vector(148, 8),
54963 => conv_std_logic_vector(149, 8),
54964 => conv_std_logic_vector(150, 8),
54965 => conv_std_logic_vector(151, 8),
54966 => conv_std_logic_vector(152, 8),
54967 => conv_std_logic_vector(152, 8),
54968 => conv_std_logic_vector(153, 8),
54969 => conv_std_logic_vector(154, 8),
54970 => conv_std_logic_vector(155, 8),
54971 => conv_std_logic_vector(156, 8),
54972 => conv_std_logic_vector(157, 8),
54973 => conv_std_logic_vector(157, 8),
54974 => conv_std_logic_vector(158, 8),
54975 => conv_std_logic_vector(159, 8),
54976 => conv_std_logic_vector(160, 8),
54977 => conv_std_logic_vector(161, 8),
54978 => conv_std_logic_vector(162, 8),
54979 => conv_std_logic_vector(163, 8),
54980 => conv_std_logic_vector(163, 8),
54981 => conv_std_logic_vector(164, 8),
54982 => conv_std_logic_vector(165, 8),
54983 => conv_std_logic_vector(166, 8),
54984 => conv_std_logic_vector(167, 8),
54985 => conv_std_logic_vector(168, 8),
54986 => conv_std_logic_vector(168, 8),
54987 => conv_std_logic_vector(169, 8),
54988 => conv_std_logic_vector(170, 8),
54989 => conv_std_logic_vector(171, 8),
54990 => conv_std_logic_vector(172, 8),
54991 => conv_std_logic_vector(173, 8),
54992 => conv_std_logic_vector(173, 8),
54993 => conv_std_logic_vector(174, 8),
54994 => conv_std_logic_vector(175, 8),
54995 => conv_std_logic_vector(176, 8),
54996 => conv_std_logic_vector(177, 8),
54997 => conv_std_logic_vector(178, 8),
54998 => conv_std_logic_vector(178, 8),
54999 => conv_std_logic_vector(179, 8),
55000 => conv_std_logic_vector(180, 8),
55001 => conv_std_logic_vector(181, 8),
55002 => conv_std_logic_vector(182, 8),
55003 => conv_std_logic_vector(183, 8),
55004 => conv_std_logic_vector(183, 8),
55005 => conv_std_logic_vector(184, 8),
55006 => conv_std_logic_vector(185, 8),
55007 => conv_std_logic_vector(186, 8),
55008 => conv_std_logic_vector(187, 8),
55009 => conv_std_logic_vector(188, 8),
55010 => conv_std_logic_vector(188, 8),
55011 => conv_std_logic_vector(189, 8),
55012 => conv_std_logic_vector(190, 8),
55013 => conv_std_logic_vector(191, 8),
55014 => conv_std_logic_vector(192, 8),
55015 => conv_std_logic_vector(193, 8),
55016 => conv_std_logic_vector(193, 8),
55017 => conv_std_logic_vector(194, 8),
55018 => conv_std_logic_vector(195, 8),
55019 => conv_std_logic_vector(196, 8),
55020 => conv_std_logic_vector(197, 8),
55021 => conv_std_logic_vector(198, 8),
55022 => conv_std_logic_vector(198, 8),
55023 => conv_std_logic_vector(199, 8),
55024 => conv_std_logic_vector(200, 8),
55025 => conv_std_logic_vector(201, 8),
55026 => conv_std_logic_vector(202, 8),
55027 => conv_std_logic_vector(203, 8),
55028 => conv_std_logic_vector(203, 8),
55029 => conv_std_logic_vector(204, 8),
55030 => conv_std_logic_vector(205, 8),
55031 => conv_std_logic_vector(206, 8),
55032 => conv_std_logic_vector(207, 8),
55033 => conv_std_logic_vector(208, 8),
55034 => conv_std_logic_vector(208, 8),
55035 => conv_std_logic_vector(209, 8),
55036 => conv_std_logic_vector(210, 8),
55037 => conv_std_logic_vector(211, 8),
55038 => conv_std_logic_vector(212, 8),
55039 => conv_std_logic_vector(213, 8),
55040 => conv_std_logic_vector(0, 8),
55041 => conv_std_logic_vector(0, 8),
55042 => conv_std_logic_vector(1, 8),
55043 => conv_std_logic_vector(2, 8),
55044 => conv_std_logic_vector(3, 8),
55045 => conv_std_logic_vector(4, 8),
55046 => conv_std_logic_vector(5, 8),
55047 => conv_std_logic_vector(5, 8),
55048 => conv_std_logic_vector(6, 8),
55049 => conv_std_logic_vector(7, 8),
55050 => conv_std_logic_vector(8, 8),
55051 => conv_std_logic_vector(9, 8),
55052 => conv_std_logic_vector(10, 8),
55053 => conv_std_logic_vector(10, 8),
55054 => conv_std_logic_vector(11, 8),
55055 => conv_std_logic_vector(12, 8),
55056 => conv_std_logic_vector(13, 8),
55057 => conv_std_logic_vector(14, 8),
55058 => conv_std_logic_vector(15, 8),
55059 => conv_std_logic_vector(15, 8),
55060 => conv_std_logic_vector(16, 8),
55061 => conv_std_logic_vector(17, 8),
55062 => conv_std_logic_vector(18, 8),
55063 => conv_std_logic_vector(19, 8),
55064 => conv_std_logic_vector(20, 8),
55065 => conv_std_logic_vector(20, 8),
55066 => conv_std_logic_vector(21, 8),
55067 => conv_std_logic_vector(22, 8),
55068 => conv_std_logic_vector(23, 8),
55069 => conv_std_logic_vector(24, 8),
55070 => conv_std_logic_vector(25, 8),
55071 => conv_std_logic_vector(26, 8),
55072 => conv_std_logic_vector(26, 8),
55073 => conv_std_logic_vector(27, 8),
55074 => conv_std_logic_vector(28, 8),
55075 => conv_std_logic_vector(29, 8),
55076 => conv_std_logic_vector(30, 8),
55077 => conv_std_logic_vector(31, 8),
55078 => conv_std_logic_vector(31, 8),
55079 => conv_std_logic_vector(32, 8),
55080 => conv_std_logic_vector(33, 8),
55081 => conv_std_logic_vector(34, 8),
55082 => conv_std_logic_vector(35, 8),
55083 => conv_std_logic_vector(36, 8),
55084 => conv_std_logic_vector(36, 8),
55085 => conv_std_logic_vector(37, 8),
55086 => conv_std_logic_vector(38, 8),
55087 => conv_std_logic_vector(39, 8),
55088 => conv_std_logic_vector(40, 8),
55089 => conv_std_logic_vector(41, 8),
55090 => conv_std_logic_vector(41, 8),
55091 => conv_std_logic_vector(42, 8),
55092 => conv_std_logic_vector(43, 8),
55093 => conv_std_logic_vector(44, 8),
55094 => conv_std_logic_vector(45, 8),
55095 => conv_std_logic_vector(46, 8),
55096 => conv_std_logic_vector(47, 8),
55097 => conv_std_logic_vector(47, 8),
55098 => conv_std_logic_vector(48, 8),
55099 => conv_std_logic_vector(49, 8),
55100 => conv_std_logic_vector(50, 8),
55101 => conv_std_logic_vector(51, 8),
55102 => conv_std_logic_vector(52, 8),
55103 => conv_std_logic_vector(52, 8),
55104 => conv_std_logic_vector(53, 8),
55105 => conv_std_logic_vector(54, 8),
55106 => conv_std_logic_vector(55, 8),
55107 => conv_std_logic_vector(56, 8),
55108 => conv_std_logic_vector(57, 8),
55109 => conv_std_logic_vector(57, 8),
55110 => conv_std_logic_vector(58, 8),
55111 => conv_std_logic_vector(59, 8),
55112 => conv_std_logic_vector(60, 8),
55113 => conv_std_logic_vector(61, 8),
55114 => conv_std_logic_vector(62, 8),
55115 => conv_std_logic_vector(62, 8),
55116 => conv_std_logic_vector(63, 8),
55117 => conv_std_logic_vector(64, 8),
55118 => conv_std_logic_vector(65, 8),
55119 => conv_std_logic_vector(66, 8),
55120 => conv_std_logic_vector(67, 8),
55121 => conv_std_logic_vector(68, 8),
55122 => conv_std_logic_vector(68, 8),
55123 => conv_std_logic_vector(69, 8),
55124 => conv_std_logic_vector(70, 8),
55125 => conv_std_logic_vector(71, 8),
55126 => conv_std_logic_vector(72, 8),
55127 => conv_std_logic_vector(73, 8),
55128 => conv_std_logic_vector(73, 8),
55129 => conv_std_logic_vector(74, 8),
55130 => conv_std_logic_vector(75, 8),
55131 => conv_std_logic_vector(76, 8),
55132 => conv_std_logic_vector(77, 8),
55133 => conv_std_logic_vector(78, 8),
55134 => conv_std_logic_vector(78, 8),
55135 => conv_std_logic_vector(79, 8),
55136 => conv_std_logic_vector(80, 8),
55137 => conv_std_logic_vector(81, 8),
55138 => conv_std_logic_vector(82, 8),
55139 => conv_std_logic_vector(83, 8),
55140 => conv_std_logic_vector(83, 8),
55141 => conv_std_logic_vector(84, 8),
55142 => conv_std_logic_vector(85, 8),
55143 => conv_std_logic_vector(86, 8),
55144 => conv_std_logic_vector(87, 8),
55145 => conv_std_logic_vector(88, 8),
55146 => conv_std_logic_vector(89, 8),
55147 => conv_std_logic_vector(89, 8),
55148 => conv_std_logic_vector(90, 8),
55149 => conv_std_logic_vector(91, 8),
55150 => conv_std_logic_vector(92, 8),
55151 => conv_std_logic_vector(93, 8),
55152 => conv_std_logic_vector(94, 8),
55153 => conv_std_logic_vector(94, 8),
55154 => conv_std_logic_vector(95, 8),
55155 => conv_std_logic_vector(96, 8),
55156 => conv_std_logic_vector(97, 8),
55157 => conv_std_logic_vector(98, 8),
55158 => conv_std_logic_vector(99, 8),
55159 => conv_std_logic_vector(99, 8),
55160 => conv_std_logic_vector(100, 8),
55161 => conv_std_logic_vector(101, 8),
55162 => conv_std_logic_vector(102, 8),
55163 => conv_std_logic_vector(103, 8),
55164 => conv_std_logic_vector(104, 8),
55165 => conv_std_logic_vector(104, 8),
55166 => conv_std_logic_vector(105, 8),
55167 => conv_std_logic_vector(106, 8),
55168 => conv_std_logic_vector(107, 8),
55169 => conv_std_logic_vector(108, 8),
55170 => conv_std_logic_vector(109, 8),
55171 => conv_std_logic_vector(110, 8),
55172 => conv_std_logic_vector(110, 8),
55173 => conv_std_logic_vector(111, 8),
55174 => conv_std_logic_vector(112, 8),
55175 => conv_std_logic_vector(113, 8),
55176 => conv_std_logic_vector(114, 8),
55177 => conv_std_logic_vector(115, 8),
55178 => conv_std_logic_vector(115, 8),
55179 => conv_std_logic_vector(116, 8),
55180 => conv_std_logic_vector(117, 8),
55181 => conv_std_logic_vector(118, 8),
55182 => conv_std_logic_vector(119, 8),
55183 => conv_std_logic_vector(120, 8),
55184 => conv_std_logic_vector(120, 8),
55185 => conv_std_logic_vector(121, 8),
55186 => conv_std_logic_vector(122, 8),
55187 => conv_std_logic_vector(123, 8),
55188 => conv_std_logic_vector(124, 8),
55189 => conv_std_logic_vector(125, 8),
55190 => conv_std_logic_vector(125, 8),
55191 => conv_std_logic_vector(126, 8),
55192 => conv_std_logic_vector(127, 8),
55193 => conv_std_logic_vector(128, 8),
55194 => conv_std_logic_vector(129, 8),
55195 => conv_std_logic_vector(130, 8),
55196 => conv_std_logic_vector(131, 8),
55197 => conv_std_logic_vector(131, 8),
55198 => conv_std_logic_vector(132, 8),
55199 => conv_std_logic_vector(133, 8),
55200 => conv_std_logic_vector(134, 8),
55201 => conv_std_logic_vector(135, 8),
55202 => conv_std_logic_vector(136, 8),
55203 => conv_std_logic_vector(136, 8),
55204 => conv_std_logic_vector(137, 8),
55205 => conv_std_logic_vector(138, 8),
55206 => conv_std_logic_vector(139, 8),
55207 => conv_std_logic_vector(140, 8),
55208 => conv_std_logic_vector(141, 8),
55209 => conv_std_logic_vector(141, 8),
55210 => conv_std_logic_vector(142, 8),
55211 => conv_std_logic_vector(143, 8),
55212 => conv_std_logic_vector(144, 8),
55213 => conv_std_logic_vector(145, 8),
55214 => conv_std_logic_vector(146, 8),
55215 => conv_std_logic_vector(146, 8),
55216 => conv_std_logic_vector(147, 8),
55217 => conv_std_logic_vector(148, 8),
55218 => conv_std_logic_vector(149, 8),
55219 => conv_std_logic_vector(150, 8),
55220 => conv_std_logic_vector(151, 8),
55221 => conv_std_logic_vector(152, 8),
55222 => conv_std_logic_vector(152, 8),
55223 => conv_std_logic_vector(153, 8),
55224 => conv_std_logic_vector(154, 8),
55225 => conv_std_logic_vector(155, 8),
55226 => conv_std_logic_vector(156, 8),
55227 => conv_std_logic_vector(157, 8),
55228 => conv_std_logic_vector(157, 8),
55229 => conv_std_logic_vector(158, 8),
55230 => conv_std_logic_vector(159, 8),
55231 => conv_std_logic_vector(160, 8),
55232 => conv_std_logic_vector(161, 8),
55233 => conv_std_logic_vector(162, 8),
55234 => conv_std_logic_vector(162, 8),
55235 => conv_std_logic_vector(163, 8),
55236 => conv_std_logic_vector(164, 8),
55237 => conv_std_logic_vector(165, 8),
55238 => conv_std_logic_vector(166, 8),
55239 => conv_std_logic_vector(167, 8),
55240 => conv_std_logic_vector(167, 8),
55241 => conv_std_logic_vector(168, 8),
55242 => conv_std_logic_vector(169, 8),
55243 => conv_std_logic_vector(170, 8),
55244 => conv_std_logic_vector(171, 8),
55245 => conv_std_logic_vector(172, 8),
55246 => conv_std_logic_vector(173, 8),
55247 => conv_std_logic_vector(173, 8),
55248 => conv_std_logic_vector(174, 8),
55249 => conv_std_logic_vector(175, 8),
55250 => conv_std_logic_vector(176, 8),
55251 => conv_std_logic_vector(177, 8),
55252 => conv_std_logic_vector(178, 8),
55253 => conv_std_logic_vector(178, 8),
55254 => conv_std_logic_vector(179, 8),
55255 => conv_std_logic_vector(180, 8),
55256 => conv_std_logic_vector(181, 8),
55257 => conv_std_logic_vector(182, 8),
55258 => conv_std_logic_vector(183, 8),
55259 => conv_std_logic_vector(183, 8),
55260 => conv_std_logic_vector(184, 8),
55261 => conv_std_logic_vector(185, 8),
55262 => conv_std_logic_vector(186, 8),
55263 => conv_std_logic_vector(187, 8),
55264 => conv_std_logic_vector(188, 8),
55265 => conv_std_logic_vector(188, 8),
55266 => conv_std_logic_vector(189, 8),
55267 => conv_std_logic_vector(190, 8),
55268 => conv_std_logic_vector(191, 8),
55269 => conv_std_logic_vector(192, 8),
55270 => conv_std_logic_vector(193, 8),
55271 => conv_std_logic_vector(194, 8),
55272 => conv_std_logic_vector(194, 8),
55273 => conv_std_logic_vector(195, 8),
55274 => conv_std_logic_vector(196, 8),
55275 => conv_std_logic_vector(197, 8),
55276 => conv_std_logic_vector(198, 8),
55277 => conv_std_logic_vector(199, 8),
55278 => conv_std_logic_vector(199, 8),
55279 => conv_std_logic_vector(200, 8),
55280 => conv_std_logic_vector(201, 8),
55281 => conv_std_logic_vector(202, 8),
55282 => conv_std_logic_vector(203, 8),
55283 => conv_std_logic_vector(204, 8),
55284 => conv_std_logic_vector(204, 8),
55285 => conv_std_logic_vector(205, 8),
55286 => conv_std_logic_vector(206, 8),
55287 => conv_std_logic_vector(207, 8),
55288 => conv_std_logic_vector(208, 8),
55289 => conv_std_logic_vector(209, 8),
55290 => conv_std_logic_vector(209, 8),
55291 => conv_std_logic_vector(210, 8),
55292 => conv_std_logic_vector(211, 8),
55293 => conv_std_logic_vector(212, 8),
55294 => conv_std_logic_vector(213, 8),
55295 => conv_std_logic_vector(214, 8),
55296 => conv_std_logic_vector(0, 8),
55297 => conv_std_logic_vector(0, 8),
55298 => conv_std_logic_vector(1, 8),
55299 => conv_std_logic_vector(2, 8),
55300 => conv_std_logic_vector(3, 8),
55301 => conv_std_logic_vector(4, 8),
55302 => conv_std_logic_vector(5, 8),
55303 => conv_std_logic_vector(5, 8),
55304 => conv_std_logic_vector(6, 8),
55305 => conv_std_logic_vector(7, 8),
55306 => conv_std_logic_vector(8, 8),
55307 => conv_std_logic_vector(9, 8),
55308 => conv_std_logic_vector(10, 8),
55309 => conv_std_logic_vector(10, 8),
55310 => conv_std_logic_vector(11, 8),
55311 => conv_std_logic_vector(12, 8),
55312 => conv_std_logic_vector(13, 8),
55313 => conv_std_logic_vector(14, 8),
55314 => conv_std_logic_vector(15, 8),
55315 => conv_std_logic_vector(16, 8),
55316 => conv_std_logic_vector(16, 8),
55317 => conv_std_logic_vector(17, 8),
55318 => conv_std_logic_vector(18, 8),
55319 => conv_std_logic_vector(19, 8),
55320 => conv_std_logic_vector(20, 8),
55321 => conv_std_logic_vector(21, 8),
55322 => conv_std_logic_vector(21, 8),
55323 => conv_std_logic_vector(22, 8),
55324 => conv_std_logic_vector(23, 8),
55325 => conv_std_logic_vector(24, 8),
55326 => conv_std_logic_vector(25, 8),
55327 => conv_std_logic_vector(26, 8),
55328 => conv_std_logic_vector(27, 8),
55329 => conv_std_logic_vector(27, 8),
55330 => conv_std_logic_vector(28, 8),
55331 => conv_std_logic_vector(29, 8),
55332 => conv_std_logic_vector(30, 8),
55333 => conv_std_logic_vector(31, 8),
55334 => conv_std_logic_vector(32, 8),
55335 => conv_std_logic_vector(32, 8),
55336 => conv_std_logic_vector(33, 8),
55337 => conv_std_logic_vector(34, 8),
55338 => conv_std_logic_vector(35, 8),
55339 => conv_std_logic_vector(36, 8),
55340 => conv_std_logic_vector(37, 8),
55341 => conv_std_logic_vector(37, 8),
55342 => conv_std_logic_vector(38, 8),
55343 => conv_std_logic_vector(39, 8),
55344 => conv_std_logic_vector(40, 8),
55345 => conv_std_logic_vector(41, 8),
55346 => conv_std_logic_vector(42, 8),
55347 => conv_std_logic_vector(43, 8),
55348 => conv_std_logic_vector(43, 8),
55349 => conv_std_logic_vector(44, 8),
55350 => conv_std_logic_vector(45, 8),
55351 => conv_std_logic_vector(46, 8),
55352 => conv_std_logic_vector(47, 8),
55353 => conv_std_logic_vector(48, 8),
55354 => conv_std_logic_vector(48, 8),
55355 => conv_std_logic_vector(49, 8),
55356 => conv_std_logic_vector(50, 8),
55357 => conv_std_logic_vector(51, 8),
55358 => conv_std_logic_vector(52, 8),
55359 => conv_std_logic_vector(53, 8),
55360 => conv_std_logic_vector(54, 8),
55361 => conv_std_logic_vector(54, 8),
55362 => conv_std_logic_vector(55, 8),
55363 => conv_std_logic_vector(56, 8),
55364 => conv_std_logic_vector(57, 8),
55365 => conv_std_logic_vector(58, 8),
55366 => conv_std_logic_vector(59, 8),
55367 => conv_std_logic_vector(59, 8),
55368 => conv_std_logic_vector(60, 8),
55369 => conv_std_logic_vector(61, 8),
55370 => conv_std_logic_vector(62, 8),
55371 => conv_std_logic_vector(63, 8),
55372 => conv_std_logic_vector(64, 8),
55373 => conv_std_logic_vector(64, 8),
55374 => conv_std_logic_vector(65, 8),
55375 => conv_std_logic_vector(66, 8),
55376 => conv_std_logic_vector(67, 8),
55377 => conv_std_logic_vector(68, 8),
55378 => conv_std_logic_vector(69, 8),
55379 => conv_std_logic_vector(70, 8),
55380 => conv_std_logic_vector(70, 8),
55381 => conv_std_logic_vector(71, 8),
55382 => conv_std_logic_vector(72, 8),
55383 => conv_std_logic_vector(73, 8),
55384 => conv_std_logic_vector(74, 8),
55385 => conv_std_logic_vector(75, 8),
55386 => conv_std_logic_vector(75, 8),
55387 => conv_std_logic_vector(76, 8),
55388 => conv_std_logic_vector(77, 8),
55389 => conv_std_logic_vector(78, 8),
55390 => conv_std_logic_vector(79, 8),
55391 => conv_std_logic_vector(80, 8),
55392 => conv_std_logic_vector(81, 8),
55393 => conv_std_logic_vector(81, 8),
55394 => conv_std_logic_vector(82, 8),
55395 => conv_std_logic_vector(83, 8),
55396 => conv_std_logic_vector(84, 8),
55397 => conv_std_logic_vector(85, 8),
55398 => conv_std_logic_vector(86, 8),
55399 => conv_std_logic_vector(86, 8),
55400 => conv_std_logic_vector(87, 8),
55401 => conv_std_logic_vector(88, 8),
55402 => conv_std_logic_vector(89, 8),
55403 => conv_std_logic_vector(90, 8),
55404 => conv_std_logic_vector(91, 8),
55405 => conv_std_logic_vector(91, 8),
55406 => conv_std_logic_vector(92, 8),
55407 => conv_std_logic_vector(93, 8),
55408 => conv_std_logic_vector(94, 8),
55409 => conv_std_logic_vector(95, 8),
55410 => conv_std_logic_vector(96, 8),
55411 => conv_std_logic_vector(97, 8),
55412 => conv_std_logic_vector(97, 8),
55413 => conv_std_logic_vector(98, 8),
55414 => conv_std_logic_vector(99, 8),
55415 => conv_std_logic_vector(100, 8),
55416 => conv_std_logic_vector(101, 8),
55417 => conv_std_logic_vector(102, 8),
55418 => conv_std_logic_vector(102, 8),
55419 => conv_std_logic_vector(103, 8),
55420 => conv_std_logic_vector(104, 8),
55421 => conv_std_logic_vector(105, 8),
55422 => conv_std_logic_vector(106, 8),
55423 => conv_std_logic_vector(107, 8),
55424 => conv_std_logic_vector(108, 8),
55425 => conv_std_logic_vector(108, 8),
55426 => conv_std_logic_vector(109, 8),
55427 => conv_std_logic_vector(110, 8),
55428 => conv_std_logic_vector(111, 8),
55429 => conv_std_logic_vector(112, 8),
55430 => conv_std_logic_vector(113, 8),
55431 => conv_std_logic_vector(113, 8),
55432 => conv_std_logic_vector(114, 8),
55433 => conv_std_logic_vector(115, 8),
55434 => conv_std_logic_vector(116, 8),
55435 => conv_std_logic_vector(117, 8),
55436 => conv_std_logic_vector(118, 8),
55437 => conv_std_logic_vector(118, 8),
55438 => conv_std_logic_vector(119, 8),
55439 => conv_std_logic_vector(120, 8),
55440 => conv_std_logic_vector(121, 8),
55441 => conv_std_logic_vector(122, 8),
55442 => conv_std_logic_vector(123, 8),
55443 => conv_std_logic_vector(124, 8),
55444 => conv_std_logic_vector(124, 8),
55445 => conv_std_logic_vector(125, 8),
55446 => conv_std_logic_vector(126, 8),
55447 => conv_std_logic_vector(127, 8),
55448 => conv_std_logic_vector(128, 8),
55449 => conv_std_logic_vector(129, 8),
55450 => conv_std_logic_vector(129, 8),
55451 => conv_std_logic_vector(130, 8),
55452 => conv_std_logic_vector(131, 8),
55453 => conv_std_logic_vector(132, 8),
55454 => conv_std_logic_vector(133, 8),
55455 => conv_std_logic_vector(134, 8),
55456 => conv_std_logic_vector(135, 8),
55457 => conv_std_logic_vector(135, 8),
55458 => conv_std_logic_vector(136, 8),
55459 => conv_std_logic_vector(137, 8),
55460 => conv_std_logic_vector(138, 8),
55461 => conv_std_logic_vector(139, 8),
55462 => conv_std_logic_vector(140, 8),
55463 => conv_std_logic_vector(140, 8),
55464 => conv_std_logic_vector(141, 8),
55465 => conv_std_logic_vector(142, 8),
55466 => conv_std_logic_vector(143, 8),
55467 => conv_std_logic_vector(144, 8),
55468 => conv_std_logic_vector(145, 8),
55469 => conv_std_logic_vector(145, 8),
55470 => conv_std_logic_vector(146, 8),
55471 => conv_std_logic_vector(147, 8),
55472 => conv_std_logic_vector(148, 8),
55473 => conv_std_logic_vector(149, 8),
55474 => conv_std_logic_vector(150, 8),
55475 => conv_std_logic_vector(151, 8),
55476 => conv_std_logic_vector(151, 8),
55477 => conv_std_logic_vector(152, 8),
55478 => conv_std_logic_vector(153, 8),
55479 => conv_std_logic_vector(154, 8),
55480 => conv_std_logic_vector(155, 8),
55481 => conv_std_logic_vector(156, 8),
55482 => conv_std_logic_vector(156, 8),
55483 => conv_std_logic_vector(157, 8),
55484 => conv_std_logic_vector(158, 8),
55485 => conv_std_logic_vector(159, 8),
55486 => conv_std_logic_vector(160, 8),
55487 => conv_std_logic_vector(161, 8),
55488 => conv_std_logic_vector(162, 8),
55489 => conv_std_logic_vector(162, 8),
55490 => conv_std_logic_vector(163, 8),
55491 => conv_std_logic_vector(164, 8),
55492 => conv_std_logic_vector(165, 8),
55493 => conv_std_logic_vector(166, 8),
55494 => conv_std_logic_vector(167, 8),
55495 => conv_std_logic_vector(167, 8),
55496 => conv_std_logic_vector(168, 8),
55497 => conv_std_logic_vector(169, 8),
55498 => conv_std_logic_vector(170, 8),
55499 => conv_std_logic_vector(171, 8),
55500 => conv_std_logic_vector(172, 8),
55501 => conv_std_logic_vector(172, 8),
55502 => conv_std_logic_vector(173, 8),
55503 => conv_std_logic_vector(174, 8),
55504 => conv_std_logic_vector(175, 8),
55505 => conv_std_logic_vector(176, 8),
55506 => conv_std_logic_vector(177, 8),
55507 => conv_std_logic_vector(178, 8),
55508 => conv_std_logic_vector(178, 8),
55509 => conv_std_logic_vector(179, 8),
55510 => conv_std_logic_vector(180, 8),
55511 => conv_std_logic_vector(181, 8),
55512 => conv_std_logic_vector(182, 8),
55513 => conv_std_logic_vector(183, 8),
55514 => conv_std_logic_vector(183, 8),
55515 => conv_std_logic_vector(184, 8),
55516 => conv_std_logic_vector(185, 8),
55517 => conv_std_logic_vector(186, 8),
55518 => conv_std_logic_vector(187, 8),
55519 => conv_std_logic_vector(188, 8),
55520 => conv_std_logic_vector(189, 8),
55521 => conv_std_logic_vector(189, 8),
55522 => conv_std_logic_vector(190, 8),
55523 => conv_std_logic_vector(191, 8),
55524 => conv_std_logic_vector(192, 8),
55525 => conv_std_logic_vector(193, 8),
55526 => conv_std_logic_vector(194, 8),
55527 => conv_std_logic_vector(194, 8),
55528 => conv_std_logic_vector(195, 8),
55529 => conv_std_logic_vector(196, 8),
55530 => conv_std_logic_vector(197, 8),
55531 => conv_std_logic_vector(198, 8),
55532 => conv_std_logic_vector(199, 8),
55533 => conv_std_logic_vector(199, 8),
55534 => conv_std_logic_vector(200, 8),
55535 => conv_std_logic_vector(201, 8),
55536 => conv_std_logic_vector(202, 8),
55537 => conv_std_logic_vector(203, 8),
55538 => conv_std_logic_vector(204, 8),
55539 => conv_std_logic_vector(205, 8),
55540 => conv_std_logic_vector(205, 8),
55541 => conv_std_logic_vector(206, 8),
55542 => conv_std_logic_vector(207, 8),
55543 => conv_std_logic_vector(208, 8),
55544 => conv_std_logic_vector(209, 8),
55545 => conv_std_logic_vector(210, 8),
55546 => conv_std_logic_vector(210, 8),
55547 => conv_std_logic_vector(211, 8),
55548 => conv_std_logic_vector(212, 8),
55549 => conv_std_logic_vector(213, 8),
55550 => conv_std_logic_vector(214, 8),
55551 => conv_std_logic_vector(215, 8),
55552 => conv_std_logic_vector(0, 8),
55553 => conv_std_logic_vector(0, 8),
55554 => conv_std_logic_vector(1, 8),
55555 => conv_std_logic_vector(2, 8),
55556 => conv_std_logic_vector(3, 8),
55557 => conv_std_logic_vector(4, 8),
55558 => conv_std_logic_vector(5, 8),
55559 => conv_std_logic_vector(5, 8),
55560 => conv_std_logic_vector(6, 8),
55561 => conv_std_logic_vector(7, 8),
55562 => conv_std_logic_vector(8, 8),
55563 => conv_std_logic_vector(9, 8),
55564 => conv_std_logic_vector(10, 8),
55565 => conv_std_logic_vector(11, 8),
55566 => conv_std_logic_vector(11, 8),
55567 => conv_std_logic_vector(12, 8),
55568 => conv_std_logic_vector(13, 8),
55569 => conv_std_logic_vector(14, 8),
55570 => conv_std_logic_vector(15, 8),
55571 => conv_std_logic_vector(16, 8),
55572 => conv_std_logic_vector(16, 8),
55573 => conv_std_logic_vector(17, 8),
55574 => conv_std_logic_vector(18, 8),
55575 => conv_std_logic_vector(19, 8),
55576 => conv_std_logic_vector(20, 8),
55577 => conv_std_logic_vector(21, 8),
55578 => conv_std_logic_vector(22, 8),
55579 => conv_std_logic_vector(22, 8),
55580 => conv_std_logic_vector(23, 8),
55581 => conv_std_logic_vector(24, 8),
55582 => conv_std_logic_vector(25, 8),
55583 => conv_std_logic_vector(26, 8),
55584 => conv_std_logic_vector(27, 8),
55585 => conv_std_logic_vector(27, 8),
55586 => conv_std_logic_vector(28, 8),
55587 => conv_std_logic_vector(29, 8),
55588 => conv_std_logic_vector(30, 8),
55589 => conv_std_logic_vector(31, 8),
55590 => conv_std_logic_vector(32, 8),
55591 => conv_std_logic_vector(33, 8),
55592 => conv_std_logic_vector(33, 8),
55593 => conv_std_logic_vector(34, 8),
55594 => conv_std_logic_vector(35, 8),
55595 => conv_std_logic_vector(36, 8),
55596 => conv_std_logic_vector(37, 8),
55597 => conv_std_logic_vector(38, 8),
55598 => conv_std_logic_vector(38, 8),
55599 => conv_std_logic_vector(39, 8),
55600 => conv_std_logic_vector(40, 8),
55601 => conv_std_logic_vector(41, 8),
55602 => conv_std_logic_vector(42, 8),
55603 => conv_std_logic_vector(43, 8),
55604 => conv_std_logic_vector(44, 8),
55605 => conv_std_logic_vector(44, 8),
55606 => conv_std_logic_vector(45, 8),
55607 => conv_std_logic_vector(46, 8),
55608 => conv_std_logic_vector(47, 8),
55609 => conv_std_logic_vector(48, 8),
55610 => conv_std_logic_vector(49, 8),
55611 => conv_std_logic_vector(50, 8),
55612 => conv_std_logic_vector(50, 8),
55613 => conv_std_logic_vector(51, 8),
55614 => conv_std_logic_vector(52, 8),
55615 => conv_std_logic_vector(53, 8),
55616 => conv_std_logic_vector(54, 8),
55617 => conv_std_logic_vector(55, 8),
55618 => conv_std_logic_vector(55, 8),
55619 => conv_std_logic_vector(56, 8),
55620 => conv_std_logic_vector(57, 8),
55621 => conv_std_logic_vector(58, 8),
55622 => conv_std_logic_vector(59, 8),
55623 => conv_std_logic_vector(60, 8),
55624 => conv_std_logic_vector(61, 8),
55625 => conv_std_logic_vector(61, 8),
55626 => conv_std_logic_vector(62, 8),
55627 => conv_std_logic_vector(63, 8),
55628 => conv_std_logic_vector(64, 8),
55629 => conv_std_logic_vector(65, 8),
55630 => conv_std_logic_vector(66, 8),
55631 => conv_std_logic_vector(66, 8),
55632 => conv_std_logic_vector(67, 8),
55633 => conv_std_logic_vector(68, 8),
55634 => conv_std_logic_vector(69, 8),
55635 => conv_std_logic_vector(70, 8),
55636 => conv_std_logic_vector(71, 8),
55637 => conv_std_logic_vector(72, 8),
55638 => conv_std_logic_vector(72, 8),
55639 => conv_std_logic_vector(73, 8),
55640 => conv_std_logic_vector(74, 8),
55641 => conv_std_logic_vector(75, 8),
55642 => conv_std_logic_vector(76, 8),
55643 => conv_std_logic_vector(77, 8),
55644 => conv_std_logic_vector(77, 8),
55645 => conv_std_logic_vector(78, 8),
55646 => conv_std_logic_vector(79, 8),
55647 => conv_std_logic_vector(80, 8),
55648 => conv_std_logic_vector(81, 8),
55649 => conv_std_logic_vector(82, 8),
55650 => conv_std_logic_vector(83, 8),
55651 => conv_std_logic_vector(83, 8),
55652 => conv_std_logic_vector(84, 8),
55653 => conv_std_logic_vector(85, 8),
55654 => conv_std_logic_vector(86, 8),
55655 => conv_std_logic_vector(87, 8),
55656 => conv_std_logic_vector(88, 8),
55657 => conv_std_logic_vector(89, 8),
55658 => conv_std_logic_vector(89, 8),
55659 => conv_std_logic_vector(90, 8),
55660 => conv_std_logic_vector(91, 8),
55661 => conv_std_logic_vector(92, 8),
55662 => conv_std_logic_vector(93, 8),
55663 => conv_std_logic_vector(94, 8),
55664 => conv_std_logic_vector(94, 8),
55665 => conv_std_logic_vector(95, 8),
55666 => conv_std_logic_vector(96, 8),
55667 => conv_std_logic_vector(97, 8),
55668 => conv_std_logic_vector(98, 8),
55669 => conv_std_logic_vector(99, 8),
55670 => conv_std_logic_vector(100, 8),
55671 => conv_std_logic_vector(100, 8),
55672 => conv_std_logic_vector(101, 8),
55673 => conv_std_logic_vector(102, 8),
55674 => conv_std_logic_vector(103, 8),
55675 => conv_std_logic_vector(104, 8),
55676 => conv_std_logic_vector(105, 8),
55677 => conv_std_logic_vector(105, 8),
55678 => conv_std_logic_vector(106, 8),
55679 => conv_std_logic_vector(107, 8),
55680 => conv_std_logic_vector(108, 8),
55681 => conv_std_logic_vector(109, 8),
55682 => conv_std_logic_vector(110, 8),
55683 => conv_std_logic_vector(111, 8),
55684 => conv_std_logic_vector(111, 8),
55685 => conv_std_logic_vector(112, 8),
55686 => conv_std_logic_vector(113, 8),
55687 => conv_std_logic_vector(114, 8),
55688 => conv_std_logic_vector(115, 8),
55689 => conv_std_logic_vector(116, 8),
55690 => conv_std_logic_vector(116, 8),
55691 => conv_std_logic_vector(117, 8),
55692 => conv_std_logic_vector(118, 8),
55693 => conv_std_logic_vector(119, 8),
55694 => conv_std_logic_vector(120, 8),
55695 => conv_std_logic_vector(121, 8),
55696 => conv_std_logic_vector(122, 8),
55697 => conv_std_logic_vector(122, 8),
55698 => conv_std_logic_vector(123, 8),
55699 => conv_std_logic_vector(124, 8),
55700 => conv_std_logic_vector(125, 8),
55701 => conv_std_logic_vector(126, 8),
55702 => conv_std_logic_vector(127, 8),
55703 => conv_std_logic_vector(127, 8),
55704 => conv_std_logic_vector(128, 8),
55705 => conv_std_logic_vector(129, 8),
55706 => conv_std_logic_vector(130, 8),
55707 => conv_std_logic_vector(131, 8),
55708 => conv_std_logic_vector(132, 8),
55709 => conv_std_logic_vector(133, 8),
55710 => conv_std_logic_vector(133, 8),
55711 => conv_std_logic_vector(134, 8),
55712 => conv_std_logic_vector(135, 8),
55713 => conv_std_logic_vector(136, 8),
55714 => conv_std_logic_vector(137, 8),
55715 => conv_std_logic_vector(138, 8),
55716 => conv_std_logic_vector(139, 8),
55717 => conv_std_logic_vector(139, 8),
55718 => conv_std_logic_vector(140, 8),
55719 => conv_std_logic_vector(141, 8),
55720 => conv_std_logic_vector(142, 8),
55721 => conv_std_logic_vector(143, 8),
55722 => conv_std_logic_vector(144, 8),
55723 => conv_std_logic_vector(144, 8),
55724 => conv_std_logic_vector(145, 8),
55725 => conv_std_logic_vector(146, 8),
55726 => conv_std_logic_vector(147, 8),
55727 => conv_std_logic_vector(148, 8),
55728 => conv_std_logic_vector(149, 8),
55729 => conv_std_logic_vector(150, 8),
55730 => conv_std_logic_vector(150, 8),
55731 => conv_std_logic_vector(151, 8),
55732 => conv_std_logic_vector(152, 8),
55733 => conv_std_logic_vector(153, 8),
55734 => conv_std_logic_vector(154, 8),
55735 => conv_std_logic_vector(155, 8),
55736 => conv_std_logic_vector(155, 8),
55737 => conv_std_logic_vector(156, 8),
55738 => conv_std_logic_vector(157, 8),
55739 => conv_std_logic_vector(158, 8),
55740 => conv_std_logic_vector(159, 8),
55741 => conv_std_logic_vector(160, 8),
55742 => conv_std_logic_vector(161, 8),
55743 => conv_std_logic_vector(161, 8),
55744 => conv_std_logic_vector(162, 8),
55745 => conv_std_logic_vector(163, 8),
55746 => conv_std_logic_vector(164, 8),
55747 => conv_std_logic_vector(165, 8),
55748 => conv_std_logic_vector(166, 8),
55749 => conv_std_logic_vector(166, 8),
55750 => conv_std_logic_vector(167, 8),
55751 => conv_std_logic_vector(168, 8),
55752 => conv_std_logic_vector(169, 8),
55753 => conv_std_logic_vector(170, 8),
55754 => conv_std_logic_vector(171, 8),
55755 => conv_std_logic_vector(172, 8),
55756 => conv_std_logic_vector(172, 8),
55757 => conv_std_logic_vector(173, 8),
55758 => conv_std_logic_vector(174, 8),
55759 => conv_std_logic_vector(175, 8),
55760 => conv_std_logic_vector(176, 8),
55761 => conv_std_logic_vector(177, 8),
55762 => conv_std_logic_vector(178, 8),
55763 => conv_std_logic_vector(178, 8),
55764 => conv_std_logic_vector(179, 8),
55765 => conv_std_logic_vector(180, 8),
55766 => conv_std_logic_vector(181, 8),
55767 => conv_std_logic_vector(182, 8),
55768 => conv_std_logic_vector(183, 8),
55769 => conv_std_logic_vector(183, 8),
55770 => conv_std_logic_vector(184, 8),
55771 => conv_std_logic_vector(185, 8),
55772 => conv_std_logic_vector(186, 8),
55773 => conv_std_logic_vector(187, 8),
55774 => conv_std_logic_vector(188, 8),
55775 => conv_std_logic_vector(189, 8),
55776 => conv_std_logic_vector(189, 8),
55777 => conv_std_logic_vector(190, 8),
55778 => conv_std_logic_vector(191, 8),
55779 => conv_std_logic_vector(192, 8),
55780 => conv_std_logic_vector(193, 8),
55781 => conv_std_logic_vector(194, 8),
55782 => conv_std_logic_vector(194, 8),
55783 => conv_std_logic_vector(195, 8),
55784 => conv_std_logic_vector(196, 8),
55785 => conv_std_logic_vector(197, 8),
55786 => conv_std_logic_vector(198, 8),
55787 => conv_std_logic_vector(199, 8),
55788 => conv_std_logic_vector(200, 8),
55789 => conv_std_logic_vector(200, 8),
55790 => conv_std_logic_vector(201, 8),
55791 => conv_std_logic_vector(202, 8),
55792 => conv_std_logic_vector(203, 8),
55793 => conv_std_logic_vector(204, 8),
55794 => conv_std_logic_vector(205, 8),
55795 => conv_std_logic_vector(205, 8),
55796 => conv_std_logic_vector(206, 8),
55797 => conv_std_logic_vector(207, 8),
55798 => conv_std_logic_vector(208, 8),
55799 => conv_std_logic_vector(209, 8),
55800 => conv_std_logic_vector(210, 8),
55801 => conv_std_logic_vector(211, 8),
55802 => conv_std_logic_vector(211, 8),
55803 => conv_std_logic_vector(212, 8),
55804 => conv_std_logic_vector(213, 8),
55805 => conv_std_logic_vector(214, 8),
55806 => conv_std_logic_vector(215, 8),
55807 => conv_std_logic_vector(216, 8),
55808 => conv_std_logic_vector(0, 8),
55809 => conv_std_logic_vector(0, 8),
55810 => conv_std_logic_vector(1, 8),
55811 => conv_std_logic_vector(2, 8),
55812 => conv_std_logic_vector(3, 8),
55813 => conv_std_logic_vector(4, 8),
55814 => conv_std_logic_vector(5, 8),
55815 => conv_std_logic_vector(5, 8),
55816 => conv_std_logic_vector(6, 8),
55817 => conv_std_logic_vector(7, 8),
55818 => conv_std_logic_vector(8, 8),
55819 => conv_std_logic_vector(9, 8),
55820 => conv_std_logic_vector(10, 8),
55821 => conv_std_logic_vector(11, 8),
55822 => conv_std_logic_vector(11, 8),
55823 => conv_std_logic_vector(12, 8),
55824 => conv_std_logic_vector(13, 8),
55825 => conv_std_logic_vector(14, 8),
55826 => conv_std_logic_vector(15, 8),
55827 => conv_std_logic_vector(16, 8),
55828 => conv_std_logic_vector(17, 8),
55829 => conv_std_logic_vector(17, 8),
55830 => conv_std_logic_vector(18, 8),
55831 => conv_std_logic_vector(19, 8),
55832 => conv_std_logic_vector(20, 8),
55833 => conv_std_logic_vector(21, 8),
55834 => conv_std_logic_vector(22, 8),
55835 => conv_std_logic_vector(22, 8),
55836 => conv_std_logic_vector(23, 8),
55837 => conv_std_logic_vector(24, 8),
55838 => conv_std_logic_vector(25, 8),
55839 => conv_std_logic_vector(26, 8),
55840 => conv_std_logic_vector(27, 8),
55841 => conv_std_logic_vector(28, 8),
55842 => conv_std_logic_vector(28, 8),
55843 => conv_std_logic_vector(29, 8),
55844 => conv_std_logic_vector(30, 8),
55845 => conv_std_logic_vector(31, 8),
55846 => conv_std_logic_vector(32, 8),
55847 => conv_std_logic_vector(33, 8),
55848 => conv_std_logic_vector(34, 8),
55849 => conv_std_logic_vector(34, 8),
55850 => conv_std_logic_vector(35, 8),
55851 => conv_std_logic_vector(36, 8),
55852 => conv_std_logic_vector(37, 8),
55853 => conv_std_logic_vector(38, 8),
55854 => conv_std_logic_vector(39, 8),
55855 => conv_std_logic_vector(40, 8),
55856 => conv_std_logic_vector(40, 8),
55857 => conv_std_logic_vector(41, 8),
55858 => conv_std_logic_vector(42, 8),
55859 => conv_std_logic_vector(43, 8),
55860 => conv_std_logic_vector(44, 8),
55861 => conv_std_logic_vector(45, 8),
55862 => conv_std_logic_vector(45, 8),
55863 => conv_std_logic_vector(46, 8),
55864 => conv_std_logic_vector(47, 8),
55865 => conv_std_logic_vector(48, 8),
55866 => conv_std_logic_vector(49, 8),
55867 => conv_std_logic_vector(50, 8),
55868 => conv_std_logic_vector(51, 8),
55869 => conv_std_logic_vector(51, 8),
55870 => conv_std_logic_vector(52, 8),
55871 => conv_std_logic_vector(53, 8),
55872 => conv_std_logic_vector(54, 8),
55873 => conv_std_logic_vector(55, 8),
55874 => conv_std_logic_vector(56, 8),
55875 => conv_std_logic_vector(57, 8),
55876 => conv_std_logic_vector(57, 8),
55877 => conv_std_logic_vector(58, 8),
55878 => conv_std_logic_vector(59, 8),
55879 => conv_std_logic_vector(60, 8),
55880 => conv_std_logic_vector(61, 8),
55881 => conv_std_logic_vector(62, 8),
55882 => conv_std_logic_vector(63, 8),
55883 => conv_std_logic_vector(63, 8),
55884 => conv_std_logic_vector(64, 8),
55885 => conv_std_logic_vector(65, 8),
55886 => conv_std_logic_vector(66, 8),
55887 => conv_std_logic_vector(67, 8),
55888 => conv_std_logic_vector(68, 8),
55889 => conv_std_logic_vector(68, 8),
55890 => conv_std_logic_vector(69, 8),
55891 => conv_std_logic_vector(70, 8),
55892 => conv_std_logic_vector(71, 8),
55893 => conv_std_logic_vector(72, 8),
55894 => conv_std_logic_vector(73, 8),
55895 => conv_std_logic_vector(74, 8),
55896 => conv_std_logic_vector(74, 8),
55897 => conv_std_logic_vector(75, 8),
55898 => conv_std_logic_vector(76, 8),
55899 => conv_std_logic_vector(77, 8),
55900 => conv_std_logic_vector(78, 8),
55901 => conv_std_logic_vector(79, 8),
55902 => conv_std_logic_vector(80, 8),
55903 => conv_std_logic_vector(80, 8),
55904 => conv_std_logic_vector(81, 8),
55905 => conv_std_logic_vector(82, 8),
55906 => conv_std_logic_vector(83, 8),
55907 => conv_std_logic_vector(84, 8),
55908 => conv_std_logic_vector(85, 8),
55909 => conv_std_logic_vector(86, 8),
55910 => conv_std_logic_vector(86, 8),
55911 => conv_std_logic_vector(87, 8),
55912 => conv_std_logic_vector(88, 8),
55913 => conv_std_logic_vector(89, 8),
55914 => conv_std_logic_vector(90, 8),
55915 => conv_std_logic_vector(91, 8),
55916 => conv_std_logic_vector(91, 8),
55917 => conv_std_logic_vector(92, 8),
55918 => conv_std_logic_vector(93, 8),
55919 => conv_std_logic_vector(94, 8),
55920 => conv_std_logic_vector(95, 8),
55921 => conv_std_logic_vector(96, 8),
55922 => conv_std_logic_vector(97, 8),
55923 => conv_std_logic_vector(97, 8),
55924 => conv_std_logic_vector(98, 8),
55925 => conv_std_logic_vector(99, 8),
55926 => conv_std_logic_vector(100, 8),
55927 => conv_std_logic_vector(101, 8),
55928 => conv_std_logic_vector(102, 8),
55929 => conv_std_logic_vector(103, 8),
55930 => conv_std_logic_vector(103, 8),
55931 => conv_std_logic_vector(104, 8),
55932 => conv_std_logic_vector(105, 8),
55933 => conv_std_logic_vector(106, 8),
55934 => conv_std_logic_vector(107, 8),
55935 => conv_std_logic_vector(108, 8),
55936 => conv_std_logic_vector(109, 8),
55937 => conv_std_logic_vector(109, 8),
55938 => conv_std_logic_vector(110, 8),
55939 => conv_std_logic_vector(111, 8),
55940 => conv_std_logic_vector(112, 8),
55941 => conv_std_logic_vector(113, 8),
55942 => conv_std_logic_vector(114, 8),
55943 => conv_std_logic_vector(114, 8),
55944 => conv_std_logic_vector(115, 8),
55945 => conv_std_logic_vector(116, 8),
55946 => conv_std_logic_vector(117, 8),
55947 => conv_std_logic_vector(118, 8),
55948 => conv_std_logic_vector(119, 8),
55949 => conv_std_logic_vector(120, 8),
55950 => conv_std_logic_vector(120, 8),
55951 => conv_std_logic_vector(121, 8),
55952 => conv_std_logic_vector(122, 8),
55953 => conv_std_logic_vector(123, 8),
55954 => conv_std_logic_vector(124, 8),
55955 => conv_std_logic_vector(125, 8),
55956 => conv_std_logic_vector(126, 8),
55957 => conv_std_logic_vector(126, 8),
55958 => conv_std_logic_vector(127, 8),
55959 => conv_std_logic_vector(128, 8),
55960 => conv_std_logic_vector(129, 8),
55961 => conv_std_logic_vector(130, 8),
55962 => conv_std_logic_vector(131, 8),
55963 => conv_std_logic_vector(131, 8),
55964 => conv_std_logic_vector(132, 8),
55965 => conv_std_logic_vector(133, 8),
55966 => conv_std_logic_vector(134, 8),
55967 => conv_std_logic_vector(135, 8),
55968 => conv_std_logic_vector(136, 8),
55969 => conv_std_logic_vector(137, 8),
55970 => conv_std_logic_vector(137, 8),
55971 => conv_std_logic_vector(138, 8),
55972 => conv_std_logic_vector(139, 8),
55973 => conv_std_logic_vector(140, 8),
55974 => conv_std_logic_vector(141, 8),
55975 => conv_std_logic_vector(142, 8),
55976 => conv_std_logic_vector(143, 8),
55977 => conv_std_logic_vector(143, 8),
55978 => conv_std_logic_vector(144, 8),
55979 => conv_std_logic_vector(145, 8),
55980 => conv_std_logic_vector(146, 8),
55981 => conv_std_logic_vector(147, 8),
55982 => conv_std_logic_vector(148, 8),
55983 => conv_std_logic_vector(149, 8),
55984 => conv_std_logic_vector(149, 8),
55985 => conv_std_logic_vector(150, 8),
55986 => conv_std_logic_vector(151, 8),
55987 => conv_std_logic_vector(152, 8),
55988 => conv_std_logic_vector(153, 8),
55989 => conv_std_logic_vector(154, 8),
55990 => conv_std_logic_vector(154, 8),
55991 => conv_std_logic_vector(155, 8),
55992 => conv_std_logic_vector(156, 8),
55993 => conv_std_logic_vector(157, 8),
55994 => conv_std_logic_vector(158, 8),
55995 => conv_std_logic_vector(159, 8),
55996 => conv_std_logic_vector(160, 8),
55997 => conv_std_logic_vector(160, 8),
55998 => conv_std_logic_vector(161, 8),
55999 => conv_std_logic_vector(162, 8),
56000 => conv_std_logic_vector(163, 8),
56001 => conv_std_logic_vector(164, 8),
56002 => conv_std_logic_vector(165, 8),
56003 => conv_std_logic_vector(166, 8),
56004 => conv_std_logic_vector(166, 8),
56005 => conv_std_logic_vector(167, 8),
56006 => conv_std_logic_vector(168, 8),
56007 => conv_std_logic_vector(169, 8),
56008 => conv_std_logic_vector(170, 8),
56009 => conv_std_logic_vector(171, 8),
56010 => conv_std_logic_vector(172, 8),
56011 => conv_std_logic_vector(172, 8),
56012 => conv_std_logic_vector(173, 8),
56013 => conv_std_logic_vector(174, 8),
56014 => conv_std_logic_vector(175, 8),
56015 => conv_std_logic_vector(176, 8),
56016 => conv_std_logic_vector(177, 8),
56017 => conv_std_logic_vector(177, 8),
56018 => conv_std_logic_vector(178, 8),
56019 => conv_std_logic_vector(179, 8),
56020 => conv_std_logic_vector(180, 8),
56021 => conv_std_logic_vector(181, 8),
56022 => conv_std_logic_vector(182, 8),
56023 => conv_std_logic_vector(183, 8),
56024 => conv_std_logic_vector(183, 8),
56025 => conv_std_logic_vector(184, 8),
56026 => conv_std_logic_vector(185, 8),
56027 => conv_std_logic_vector(186, 8),
56028 => conv_std_logic_vector(187, 8),
56029 => conv_std_logic_vector(188, 8),
56030 => conv_std_logic_vector(189, 8),
56031 => conv_std_logic_vector(189, 8),
56032 => conv_std_logic_vector(190, 8),
56033 => conv_std_logic_vector(191, 8),
56034 => conv_std_logic_vector(192, 8),
56035 => conv_std_logic_vector(193, 8),
56036 => conv_std_logic_vector(194, 8),
56037 => conv_std_logic_vector(195, 8),
56038 => conv_std_logic_vector(195, 8),
56039 => conv_std_logic_vector(196, 8),
56040 => conv_std_logic_vector(197, 8),
56041 => conv_std_logic_vector(198, 8),
56042 => conv_std_logic_vector(199, 8),
56043 => conv_std_logic_vector(200, 8),
56044 => conv_std_logic_vector(200, 8),
56045 => conv_std_logic_vector(201, 8),
56046 => conv_std_logic_vector(202, 8),
56047 => conv_std_logic_vector(203, 8),
56048 => conv_std_logic_vector(204, 8),
56049 => conv_std_logic_vector(205, 8),
56050 => conv_std_logic_vector(206, 8),
56051 => conv_std_logic_vector(206, 8),
56052 => conv_std_logic_vector(207, 8),
56053 => conv_std_logic_vector(208, 8),
56054 => conv_std_logic_vector(209, 8),
56055 => conv_std_logic_vector(210, 8),
56056 => conv_std_logic_vector(211, 8),
56057 => conv_std_logic_vector(212, 8),
56058 => conv_std_logic_vector(212, 8),
56059 => conv_std_logic_vector(213, 8),
56060 => conv_std_logic_vector(214, 8),
56061 => conv_std_logic_vector(215, 8),
56062 => conv_std_logic_vector(216, 8),
56063 => conv_std_logic_vector(217, 8),
56064 => conv_std_logic_vector(0, 8),
56065 => conv_std_logic_vector(0, 8),
56066 => conv_std_logic_vector(1, 8),
56067 => conv_std_logic_vector(2, 8),
56068 => conv_std_logic_vector(3, 8),
56069 => conv_std_logic_vector(4, 8),
56070 => conv_std_logic_vector(5, 8),
56071 => conv_std_logic_vector(5, 8),
56072 => conv_std_logic_vector(6, 8),
56073 => conv_std_logic_vector(7, 8),
56074 => conv_std_logic_vector(8, 8),
56075 => conv_std_logic_vector(9, 8),
56076 => conv_std_logic_vector(10, 8),
56077 => conv_std_logic_vector(11, 8),
56078 => conv_std_logic_vector(11, 8),
56079 => conv_std_logic_vector(12, 8),
56080 => conv_std_logic_vector(13, 8),
56081 => conv_std_logic_vector(14, 8),
56082 => conv_std_logic_vector(15, 8),
56083 => conv_std_logic_vector(16, 8),
56084 => conv_std_logic_vector(17, 8),
56085 => conv_std_logic_vector(17, 8),
56086 => conv_std_logic_vector(18, 8),
56087 => conv_std_logic_vector(19, 8),
56088 => conv_std_logic_vector(20, 8),
56089 => conv_std_logic_vector(21, 8),
56090 => conv_std_logic_vector(22, 8),
56091 => conv_std_logic_vector(23, 8),
56092 => conv_std_logic_vector(23, 8),
56093 => conv_std_logic_vector(24, 8),
56094 => conv_std_logic_vector(25, 8),
56095 => conv_std_logic_vector(26, 8),
56096 => conv_std_logic_vector(27, 8),
56097 => conv_std_logic_vector(28, 8),
56098 => conv_std_logic_vector(29, 8),
56099 => conv_std_logic_vector(29, 8),
56100 => conv_std_logic_vector(30, 8),
56101 => conv_std_logic_vector(31, 8),
56102 => conv_std_logic_vector(32, 8),
56103 => conv_std_logic_vector(33, 8),
56104 => conv_std_logic_vector(34, 8),
56105 => conv_std_logic_vector(35, 8),
56106 => conv_std_logic_vector(35, 8),
56107 => conv_std_logic_vector(36, 8),
56108 => conv_std_logic_vector(37, 8),
56109 => conv_std_logic_vector(38, 8),
56110 => conv_std_logic_vector(39, 8),
56111 => conv_std_logic_vector(40, 8),
56112 => conv_std_logic_vector(41, 8),
56113 => conv_std_logic_vector(41, 8),
56114 => conv_std_logic_vector(42, 8),
56115 => conv_std_logic_vector(43, 8),
56116 => conv_std_logic_vector(44, 8),
56117 => conv_std_logic_vector(45, 8),
56118 => conv_std_logic_vector(46, 8),
56119 => conv_std_logic_vector(47, 8),
56120 => conv_std_logic_vector(47, 8),
56121 => conv_std_logic_vector(48, 8),
56122 => conv_std_logic_vector(49, 8),
56123 => conv_std_logic_vector(50, 8),
56124 => conv_std_logic_vector(51, 8),
56125 => conv_std_logic_vector(52, 8),
56126 => conv_std_logic_vector(53, 8),
56127 => conv_std_logic_vector(53, 8),
56128 => conv_std_logic_vector(54, 8),
56129 => conv_std_logic_vector(55, 8),
56130 => conv_std_logic_vector(56, 8),
56131 => conv_std_logic_vector(57, 8),
56132 => conv_std_logic_vector(58, 8),
56133 => conv_std_logic_vector(59, 8),
56134 => conv_std_logic_vector(59, 8),
56135 => conv_std_logic_vector(60, 8),
56136 => conv_std_logic_vector(61, 8),
56137 => conv_std_logic_vector(62, 8),
56138 => conv_std_logic_vector(63, 8),
56139 => conv_std_logic_vector(64, 8),
56140 => conv_std_logic_vector(65, 8),
56141 => conv_std_logic_vector(65, 8),
56142 => conv_std_logic_vector(66, 8),
56143 => conv_std_logic_vector(67, 8),
56144 => conv_std_logic_vector(68, 8),
56145 => conv_std_logic_vector(69, 8),
56146 => conv_std_logic_vector(70, 8),
56147 => conv_std_logic_vector(71, 8),
56148 => conv_std_logic_vector(71, 8),
56149 => conv_std_logic_vector(72, 8),
56150 => conv_std_logic_vector(73, 8),
56151 => conv_std_logic_vector(74, 8),
56152 => conv_std_logic_vector(75, 8),
56153 => conv_std_logic_vector(76, 8),
56154 => conv_std_logic_vector(76, 8),
56155 => conv_std_logic_vector(77, 8),
56156 => conv_std_logic_vector(78, 8),
56157 => conv_std_logic_vector(79, 8),
56158 => conv_std_logic_vector(80, 8),
56159 => conv_std_logic_vector(81, 8),
56160 => conv_std_logic_vector(82, 8),
56161 => conv_std_logic_vector(82, 8),
56162 => conv_std_logic_vector(83, 8),
56163 => conv_std_logic_vector(84, 8),
56164 => conv_std_logic_vector(85, 8),
56165 => conv_std_logic_vector(86, 8),
56166 => conv_std_logic_vector(87, 8),
56167 => conv_std_logic_vector(88, 8),
56168 => conv_std_logic_vector(88, 8),
56169 => conv_std_logic_vector(89, 8),
56170 => conv_std_logic_vector(90, 8),
56171 => conv_std_logic_vector(91, 8),
56172 => conv_std_logic_vector(92, 8),
56173 => conv_std_logic_vector(93, 8),
56174 => conv_std_logic_vector(94, 8),
56175 => conv_std_logic_vector(94, 8),
56176 => conv_std_logic_vector(95, 8),
56177 => conv_std_logic_vector(96, 8),
56178 => conv_std_logic_vector(97, 8),
56179 => conv_std_logic_vector(98, 8),
56180 => conv_std_logic_vector(99, 8),
56181 => conv_std_logic_vector(100, 8),
56182 => conv_std_logic_vector(100, 8),
56183 => conv_std_logic_vector(101, 8),
56184 => conv_std_logic_vector(102, 8),
56185 => conv_std_logic_vector(103, 8),
56186 => conv_std_logic_vector(104, 8),
56187 => conv_std_logic_vector(105, 8),
56188 => conv_std_logic_vector(106, 8),
56189 => conv_std_logic_vector(106, 8),
56190 => conv_std_logic_vector(107, 8),
56191 => conv_std_logic_vector(108, 8),
56192 => conv_std_logic_vector(109, 8),
56193 => conv_std_logic_vector(110, 8),
56194 => conv_std_logic_vector(111, 8),
56195 => conv_std_logic_vector(112, 8),
56196 => conv_std_logic_vector(112, 8),
56197 => conv_std_logic_vector(113, 8),
56198 => conv_std_logic_vector(114, 8),
56199 => conv_std_logic_vector(115, 8),
56200 => conv_std_logic_vector(116, 8),
56201 => conv_std_logic_vector(117, 8),
56202 => conv_std_logic_vector(118, 8),
56203 => conv_std_logic_vector(118, 8),
56204 => conv_std_logic_vector(119, 8),
56205 => conv_std_logic_vector(120, 8),
56206 => conv_std_logic_vector(121, 8),
56207 => conv_std_logic_vector(122, 8),
56208 => conv_std_logic_vector(123, 8),
56209 => conv_std_logic_vector(124, 8),
56210 => conv_std_logic_vector(124, 8),
56211 => conv_std_logic_vector(125, 8),
56212 => conv_std_logic_vector(126, 8),
56213 => conv_std_logic_vector(127, 8),
56214 => conv_std_logic_vector(128, 8),
56215 => conv_std_logic_vector(129, 8),
56216 => conv_std_logic_vector(130, 8),
56217 => conv_std_logic_vector(130, 8),
56218 => conv_std_logic_vector(131, 8),
56219 => conv_std_logic_vector(132, 8),
56220 => conv_std_logic_vector(133, 8),
56221 => conv_std_logic_vector(134, 8),
56222 => conv_std_logic_vector(135, 8),
56223 => conv_std_logic_vector(136, 8),
56224 => conv_std_logic_vector(136, 8),
56225 => conv_std_logic_vector(137, 8),
56226 => conv_std_logic_vector(138, 8),
56227 => conv_std_logic_vector(139, 8),
56228 => conv_std_logic_vector(140, 8),
56229 => conv_std_logic_vector(141, 8),
56230 => conv_std_logic_vector(142, 8),
56231 => conv_std_logic_vector(142, 8),
56232 => conv_std_logic_vector(143, 8),
56233 => conv_std_logic_vector(144, 8),
56234 => conv_std_logic_vector(145, 8),
56235 => conv_std_logic_vector(146, 8),
56236 => conv_std_logic_vector(147, 8),
56237 => conv_std_logic_vector(147, 8),
56238 => conv_std_logic_vector(148, 8),
56239 => conv_std_logic_vector(149, 8),
56240 => conv_std_logic_vector(150, 8),
56241 => conv_std_logic_vector(151, 8),
56242 => conv_std_logic_vector(152, 8),
56243 => conv_std_logic_vector(153, 8),
56244 => conv_std_logic_vector(153, 8),
56245 => conv_std_logic_vector(154, 8),
56246 => conv_std_logic_vector(155, 8),
56247 => conv_std_logic_vector(156, 8),
56248 => conv_std_logic_vector(157, 8),
56249 => conv_std_logic_vector(158, 8),
56250 => conv_std_logic_vector(159, 8),
56251 => conv_std_logic_vector(159, 8),
56252 => conv_std_logic_vector(160, 8),
56253 => conv_std_logic_vector(161, 8),
56254 => conv_std_logic_vector(162, 8),
56255 => conv_std_logic_vector(163, 8),
56256 => conv_std_logic_vector(164, 8),
56257 => conv_std_logic_vector(165, 8),
56258 => conv_std_logic_vector(165, 8),
56259 => conv_std_logic_vector(166, 8),
56260 => conv_std_logic_vector(167, 8),
56261 => conv_std_logic_vector(168, 8),
56262 => conv_std_logic_vector(169, 8),
56263 => conv_std_logic_vector(170, 8),
56264 => conv_std_logic_vector(171, 8),
56265 => conv_std_logic_vector(171, 8),
56266 => conv_std_logic_vector(172, 8),
56267 => conv_std_logic_vector(173, 8),
56268 => conv_std_logic_vector(174, 8),
56269 => conv_std_logic_vector(175, 8),
56270 => conv_std_logic_vector(176, 8),
56271 => conv_std_logic_vector(177, 8),
56272 => conv_std_logic_vector(177, 8),
56273 => conv_std_logic_vector(178, 8),
56274 => conv_std_logic_vector(179, 8),
56275 => conv_std_logic_vector(180, 8),
56276 => conv_std_logic_vector(181, 8),
56277 => conv_std_logic_vector(182, 8),
56278 => conv_std_logic_vector(183, 8),
56279 => conv_std_logic_vector(183, 8),
56280 => conv_std_logic_vector(184, 8),
56281 => conv_std_logic_vector(185, 8),
56282 => conv_std_logic_vector(186, 8),
56283 => conv_std_logic_vector(187, 8),
56284 => conv_std_logic_vector(188, 8),
56285 => conv_std_logic_vector(189, 8),
56286 => conv_std_logic_vector(189, 8),
56287 => conv_std_logic_vector(190, 8),
56288 => conv_std_logic_vector(191, 8),
56289 => conv_std_logic_vector(192, 8),
56290 => conv_std_logic_vector(193, 8),
56291 => conv_std_logic_vector(194, 8),
56292 => conv_std_logic_vector(195, 8),
56293 => conv_std_logic_vector(195, 8),
56294 => conv_std_logic_vector(196, 8),
56295 => conv_std_logic_vector(197, 8),
56296 => conv_std_logic_vector(198, 8),
56297 => conv_std_logic_vector(199, 8),
56298 => conv_std_logic_vector(200, 8),
56299 => conv_std_logic_vector(201, 8),
56300 => conv_std_logic_vector(201, 8),
56301 => conv_std_logic_vector(202, 8),
56302 => conv_std_logic_vector(203, 8),
56303 => conv_std_logic_vector(204, 8),
56304 => conv_std_logic_vector(205, 8),
56305 => conv_std_logic_vector(206, 8),
56306 => conv_std_logic_vector(207, 8),
56307 => conv_std_logic_vector(207, 8),
56308 => conv_std_logic_vector(208, 8),
56309 => conv_std_logic_vector(209, 8),
56310 => conv_std_logic_vector(210, 8),
56311 => conv_std_logic_vector(211, 8),
56312 => conv_std_logic_vector(212, 8),
56313 => conv_std_logic_vector(213, 8),
56314 => conv_std_logic_vector(213, 8),
56315 => conv_std_logic_vector(214, 8),
56316 => conv_std_logic_vector(215, 8),
56317 => conv_std_logic_vector(216, 8),
56318 => conv_std_logic_vector(217, 8),
56319 => conv_std_logic_vector(218, 8),
56320 => conv_std_logic_vector(0, 8),
56321 => conv_std_logic_vector(0, 8),
56322 => conv_std_logic_vector(1, 8),
56323 => conv_std_logic_vector(2, 8),
56324 => conv_std_logic_vector(3, 8),
56325 => conv_std_logic_vector(4, 8),
56326 => conv_std_logic_vector(5, 8),
56327 => conv_std_logic_vector(6, 8),
56328 => conv_std_logic_vector(6, 8),
56329 => conv_std_logic_vector(7, 8),
56330 => conv_std_logic_vector(8, 8),
56331 => conv_std_logic_vector(9, 8),
56332 => conv_std_logic_vector(10, 8),
56333 => conv_std_logic_vector(11, 8),
56334 => conv_std_logic_vector(12, 8),
56335 => conv_std_logic_vector(12, 8),
56336 => conv_std_logic_vector(13, 8),
56337 => conv_std_logic_vector(14, 8),
56338 => conv_std_logic_vector(15, 8),
56339 => conv_std_logic_vector(16, 8),
56340 => conv_std_logic_vector(17, 8),
56341 => conv_std_logic_vector(18, 8),
56342 => conv_std_logic_vector(18, 8),
56343 => conv_std_logic_vector(19, 8),
56344 => conv_std_logic_vector(20, 8),
56345 => conv_std_logic_vector(21, 8),
56346 => conv_std_logic_vector(22, 8),
56347 => conv_std_logic_vector(23, 8),
56348 => conv_std_logic_vector(24, 8),
56349 => conv_std_logic_vector(24, 8),
56350 => conv_std_logic_vector(25, 8),
56351 => conv_std_logic_vector(26, 8),
56352 => conv_std_logic_vector(27, 8),
56353 => conv_std_logic_vector(28, 8),
56354 => conv_std_logic_vector(29, 8),
56355 => conv_std_logic_vector(30, 8),
56356 => conv_std_logic_vector(30, 8),
56357 => conv_std_logic_vector(31, 8),
56358 => conv_std_logic_vector(32, 8),
56359 => conv_std_logic_vector(33, 8),
56360 => conv_std_logic_vector(34, 8),
56361 => conv_std_logic_vector(35, 8),
56362 => conv_std_logic_vector(36, 8),
56363 => conv_std_logic_vector(36, 8),
56364 => conv_std_logic_vector(37, 8),
56365 => conv_std_logic_vector(38, 8),
56366 => conv_std_logic_vector(39, 8),
56367 => conv_std_logic_vector(40, 8),
56368 => conv_std_logic_vector(41, 8),
56369 => conv_std_logic_vector(42, 8),
56370 => conv_std_logic_vector(42, 8),
56371 => conv_std_logic_vector(43, 8),
56372 => conv_std_logic_vector(44, 8),
56373 => conv_std_logic_vector(45, 8),
56374 => conv_std_logic_vector(46, 8),
56375 => conv_std_logic_vector(47, 8),
56376 => conv_std_logic_vector(48, 8),
56377 => conv_std_logic_vector(48, 8),
56378 => conv_std_logic_vector(49, 8),
56379 => conv_std_logic_vector(50, 8),
56380 => conv_std_logic_vector(51, 8),
56381 => conv_std_logic_vector(52, 8),
56382 => conv_std_logic_vector(53, 8),
56383 => conv_std_logic_vector(54, 8),
56384 => conv_std_logic_vector(55, 8),
56385 => conv_std_logic_vector(55, 8),
56386 => conv_std_logic_vector(56, 8),
56387 => conv_std_logic_vector(57, 8),
56388 => conv_std_logic_vector(58, 8),
56389 => conv_std_logic_vector(59, 8),
56390 => conv_std_logic_vector(60, 8),
56391 => conv_std_logic_vector(61, 8),
56392 => conv_std_logic_vector(61, 8),
56393 => conv_std_logic_vector(62, 8),
56394 => conv_std_logic_vector(63, 8),
56395 => conv_std_logic_vector(64, 8),
56396 => conv_std_logic_vector(65, 8),
56397 => conv_std_logic_vector(66, 8),
56398 => conv_std_logic_vector(67, 8),
56399 => conv_std_logic_vector(67, 8),
56400 => conv_std_logic_vector(68, 8),
56401 => conv_std_logic_vector(69, 8),
56402 => conv_std_logic_vector(70, 8),
56403 => conv_std_logic_vector(71, 8),
56404 => conv_std_logic_vector(72, 8),
56405 => conv_std_logic_vector(73, 8),
56406 => conv_std_logic_vector(73, 8),
56407 => conv_std_logic_vector(74, 8),
56408 => conv_std_logic_vector(75, 8),
56409 => conv_std_logic_vector(76, 8),
56410 => conv_std_logic_vector(77, 8),
56411 => conv_std_logic_vector(78, 8),
56412 => conv_std_logic_vector(79, 8),
56413 => conv_std_logic_vector(79, 8),
56414 => conv_std_logic_vector(80, 8),
56415 => conv_std_logic_vector(81, 8),
56416 => conv_std_logic_vector(82, 8),
56417 => conv_std_logic_vector(83, 8),
56418 => conv_std_logic_vector(84, 8),
56419 => conv_std_logic_vector(85, 8),
56420 => conv_std_logic_vector(85, 8),
56421 => conv_std_logic_vector(86, 8),
56422 => conv_std_logic_vector(87, 8),
56423 => conv_std_logic_vector(88, 8),
56424 => conv_std_logic_vector(89, 8),
56425 => conv_std_logic_vector(90, 8),
56426 => conv_std_logic_vector(91, 8),
56427 => conv_std_logic_vector(91, 8),
56428 => conv_std_logic_vector(92, 8),
56429 => conv_std_logic_vector(93, 8),
56430 => conv_std_logic_vector(94, 8),
56431 => conv_std_logic_vector(95, 8),
56432 => conv_std_logic_vector(96, 8),
56433 => conv_std_logic_vector(97, 8),
56434 => conv_std_logic_vector(97, 8),
56435 => conv_std_logic_vector(98, 8),
56436 => conv_std_logic_vector(99, 8),
56437 => conv_std_logic_vector(100, 8),
56438 => conv_std_logic_vector(101, 8),
56439 => conv_std_logic_vector(102, 8),
56440 => conv_std_logic_vector(103, 8),
56441 => conv_std_logic_vector(103, 8),
56442 => conv_std_logic_vector(104, 8),
56443 => conv_std_logic_vector(105, 8),
56444 => conv_std_logic_vector(106, 8),
56445 => conv_std_logic_vector(107, 8),
56446 => conv_std_logic_vector(108, 8),
56447 => conv_std_logic_vector(109, 8),
56448 => conv_std_logic_vector(110, 8),
56449 => conv_std_logic_vector(110, 8),
56450 => conv_std_logic_vector(111, 8),
56451 => conv_std_logic_vector(112, 8),
56452 => conv_std_logic_vector(113, 8),
56453 => conv_std_logic_vector(114, 8),
56454 => conv_std_logic_vector(115, 8),
56455 => conv_std_logic_vector(116, 8),
56456 => conv_std_logic_vector(116, 8),
56457 => conv_std_logic_vector(117, 8),
56458 => conv_std_logic_vector(118, 8),
56459 => conv_std_logic_vector(119, 8),
56460 => conv_std_logic_vector(120, 8),
56461 => conv_std_logic_vector(121, 8),
56462 => conv_std_logic_vector(122, 8),
56463 => conv_std_logic_vector(122, 8),
56464 => conv_std_logic_vector(123, 8),
56465 => conv_std_logic_vector(124, 8),
56466 => conv_std_logic_vector(125, 8),
56467 => conv_std_logic_vector(126, 8),
56468 => conv_std_logic_vector(127, 8),
56469 => conv_std_logic_vector(128, 8),
56470 => conv_std_logic_vector(128, 8),
56471 => conv_std_logic_vector(129, 8),
56472 => conv_std_logic_vector(130, 8),
56473 => conv_std_logic_vector(131, 8),
56474 => conv_std_logic_vector(132, 8),
56475 => conv_std_logic_vector(133, 8),
56476 => conv_std_logic_vector(134, 8),
56477 => conv_std_logic_vector(134, 8),
56478 => conv_std_logic_vector(135, 8),
56479 => conv_std_logic_vector(136, 8),
56480 => conv_std_logic_vector(137, 8),
56481 => conv_std_logic_vector(138, 8),
56482 => conv_std_logic_vector(139, 8),
56483 => conv_std_logic_vector(140, 8),
56484 => conv_std_logic_vector(140, 8),
56485 => conv_std_logic_vector(141, 8),
56486 => conv_std_logic_vector(142, 8),
56487 => conv_std_logic_vector(143, 8),
56488 => conv_std_logic_vector(144, 8),
56489 => conv_std_logic_vector(145, 8),
56490 => conv_std_logic_vector(146, 8),
56491 => conv_std_logic_vector(146, 8),
56492 => conv_std_logic_vector(147, 8),
56493 => conv_std_logic_vector(148, 8),
56494 => conv_std_logic_vector(149, 8),
56495 => conv_std_logic_vector(150, 8),
56496 => conv_std_logic_vector(151, 8),
56497 => conv_std_logic_vector(152, 8),
56498 => conv_std_logic_vector(152, 8),
56499 => conv_std_logic_vector(153, 8),
56500 => conv_std_logic_vector(154, 8),
56501 => conv_std_logic_vector(155, 8),
56502 => conv_std_logic_vector(156, 8),
56503 => conv_std_logic_vector(157, 8),
56504 => conv_std_logic_vector(158, 8),
56505 => conv_std_logic_vector(158, 8),
56506 => conv_std_logic_vector(159, 8),
56507 => conv_std_logic_vector(160, 8),
56508 => conv_std_logic_vector(161, 8),
56509 => conv_std_logic_vector(162, 8),
56510 => conv_std_logic_vector(163, 8),
56511 => conv_std_logic_vector(164, 8),
56512 => conv_std_logic_vector(165, 8),
56513 => conv_std_logic_vector(165, 8),
56514 => conv_std_logic_vector(166, 8),
56515 => conv_std_logic_vector(167, 8),
56516 => conv_std_logic_vector(168, 8),
56517 => conv_std_logic_vector(169, 8),
56518 => conv_std_logic_vector(170, 8),
56519 => conv_std_logic_vector(171, 8),
56520 => conv_std_logic_vector(171, 8),
56521 => conv_std_logic_vector(172, 8),
56522 => conv_std_logic_vector(173, 8),
56523 => conv_std_logic_vector(174, 8),
56524 => conv_std_logic_vector(175, 8),
56525 => conv_std_logic_vector(176, 8),
56526 => conv_std_logic_vector(177, 8),
56527 => conv_std_logic_vector(177, 8),
56528 => conv_std_logic_vector(178, 8),
56529 => conv_std_logic_vector(179, 8),
56530 => conv_std_logic_vector(180, 8),
56531 => conv_std_logic_vector(181, 8),
56532 => conv_std_logic_vector(182, 8),
56533 => conv_std_logic_vector(183, 8),
56534 => conv_std_logic_vector(183, 8),
56535 => conv_std_logic_vector(184, 8),
56536 => conv_std_logic_vector(185, 8),
56537 => conv_std_logic_vector(186, 8),
56538 => conv_std_logic_vector(187, 8),
56539 => conv_std_logic_vector(188, 8),
56540 => conv_std_logic_vector(189, 8),
56541 => conv_std_logic_vector(189, 8),
56542 => conv_std_logic_vector(190, 8),
56543 => conv_std_logic_vector(191, 8),
56544 => conv_std_logic_vector(192, 8),
56545 => conv_std_logic_vector(193, 8),
56546 => conv_std_logic_vector(194, 8),
56547 => conv_std_logic_vector(195, 8),
56548 => conv_std_logic_vector(195, 8),
56549 => conv_std_logic_vector(196, 8),
56550 => conv_std_logic_vector(197, 8),
56551 => conv_std_logic_vector(198, 8),
56552 => conv_std_logic_vector(199, 8),
56553 => conv_std_logic_vector(200, 8),
56554 => conv_std_logic_vector(201, 8),
56555 => conv_std_logic_vector(201, 8),
56556 => conv_std_logic_vector(202, 8),
56557 => conv_std_logic_vector(203, 8),
56558 => conv_std_logic_vector(204, 8),
56559 => conv_std_logic_vector(205, 8),
56560 => conv_std_logic_vector(206, 8),
56561 => conv_std_logic_vector(207, 8),
56562 => conv_std_logic_vector(207, 8),
56563 => conv_std_logic_vector(208, 8),
56564 => conv_std_logic_vector(209, 8),
56565 => conv_std_logic_vector(210, 8),
56566 => conv_std_logic_vector(211, 8),
56567 => conv_std_logic_vector(212, 8),
56568 => conv_std_logic_vector(213, 8),
56569 => conv_std_logic_vector(213, 8),
56570 => conv_std_logic_vector(214, 8),
56571 => conv_std_logic_vector(215, 8),
56572 => conv_std_logic_vector(216, 8),
56573 => conv_std_logic_vector(217, 8),
56574 => conv_std_logic_vector(218, 8),
56575 => conv_std_logic_vector(219, 8),
56576 => conv_std_logic_vector(0, 8),
56577 => conv_std_logic_vector(0, 8),
56578 => conv_std_logic_vector(1, 8),
56579 => conv_std_logic_vector(2, 8),
56580 => conv_std_logic_vector(3, 8),
56581 => conv_std_logic_vector(4, 8),
56582 => conv_std_logic_vector(5, 8),
56583 => conv_std_logic_vector(6, 8),
56584 => conv_std_logic_vector(6, 8),
56585 => conv_std_logic_vector(7, 8),
56586 => conv_std_logic_vector(8, 8),
56587 => conv_std_logic_vector(9, 8),
56588 => conv_std_logic_vector(10, 8),
56589 => conv_std_logic_vector(11, 8),
56590 => conv_std_logic_vector(12, 8),
56591 => conv_std_logic_vector(12, 8),
56592 => conv_std_logic_vector(13, 8),
56593 => conv_std_logic_vector(14, 8),
56594 => conv_std_logic_vector(15, 8),
56595 => conv_std_logic_vector(16, 8),
56596 => conv_std_logic_vector(17, 8),
56597 => conv_std_logic_vector(18, 8),
56598 => conv_std_logic_vector(18, 8),
56599 => conv_std_logic_vector(19, 8),
56600 => conv_std_logic_vector(20, 8),
56601 => conv_std_logic_vector(21, 8),
56602 => conv_std_logic_vector(22, 8),
56603 => conv_std_logic_vector(23, 8),
56604 => conv_std_logic_vector(24, 8),
56605 => conv_std_logic_vector(25, 8),
56606 => conv_std_logic_vector(25, 8),
56607 => conv_std_logic_vector(26, 8),
56608 => conv_std_logic_vector(27, 8),
56609 => conv_std_logic_vector(28, 8),
56610 => conv_std_logic_vector(29, 8),
56611 => conv_std_logic_vector(30, 8),
56612 => conv_std_logic_vector(31, 8),
56613 => conv_std_logic_vector(31, 8),
56614 => conv_std_logic_vector(32, 8),
56615 => conv_std_logic_vector(33, 8),
56616 => conv_std_logic_vector(34, 8),
56617 => conv_std_logic_vector(35, 8),
56618 => conv_std_logic_vector(36, 8),
56619 => conv_std_logic_vector(37, 8),
56620 => conv_std_logic_vector(37, 8),
56621 => conv_std_logic_vector(38, 8),
56622 => conv_std_logic_vector(39, 8),
56623 => conv_std_logic_vector(40, 8),
56624 => conv_std_logic_vector(41, 8),
56625 => conv_std_logic_vector(42, 8),
56626 => conv_std_logic_vector(43, 8),
56627 => conv_std_logic_vector(44, 8),
56628 => conv_std_logic_vector(44, 8),
56629 => conv_std_logic_vector(45, 8),
56630 => conv_std_logic_vector(46, 8),
56631 => conv_std_logic_vector(47, 8),
56632 => conv_std_logic_vector(48, 8),
56633 => conv_std_logic_vector(49, 8),
56634 => conv_std_logic_vector(50, 8),
56635 => conv_std_logic_vector(50, 8),
56636 => conv_std_logic_vector(51, 8),
56637 => conv_std_logic_vector(52, 8),
56638 => conv_std_logic_vector(53, 8),
56639 => conv_std_logic_vector(54, 8),
56640 => conv_std_logic_vector(55, 8),
56641 => conv_std_logic_vector(56, 8),
56642 => conv_std_logic_vector(56, 8),
56643 => conv_std_logic_vector(57, 8),
56644 => conv_std_logic_vector(58, 8),
56645 => conv_std_logic_vector(59, 8),
56646 => conv_std_logic_vector(60, 8),
56647 => conv_std_logic_vector(61, 8),
56648 => conv_std_logic_vector(62, 8),
56649 => conv_std_logic_vector(63, 8),
56650 => conv_std_logic_vector(63, 8),
56651 => conv_std_logic_vector(64, 8),
56652 => conv_std_logic_vector(65, 8),
56653 => conv_std_logic_vector(66, 8),
56654 => conv_std_logic_vector(67, 8),
56655 => conv_std_logic_vector(68, 8),
56656 => conv_std_logic_vector(69, 8),
56657 => conv_std_logic_vector(69, 8),
56658 => conv_std_logic_vector(70, 8),
56659 => conv_std_logic_vector(71, 8),
56660 => conv_std_logic_vector(72, 8),
56661 => conv_std_logic_vector(73, 8),
56662 => conv_std_logic_vector(74, 8),
56663 => conv_std_logic_vector(75, 8),
56664 => conv_std_logic_vector(75, 8),
56665 => conv_std_logic_vector(76, 8),
56666 => conv_std_logic_vector(77, 8),
56667 => conv_std_logic_vector(78, 8),
56668 => conv_std_logic_vector(79, 8),
56669 => conv_std_logic_vector(80, 8),
56670 => conv_std_logic_vector(81, 8),
56671 => conv_std_logic_vector(82, 8),
56672 => conv_std_logic_vector(82, 8),
56673 => conv_std_logic_vector(83, 8),
56674 => conv_std_logic_vector(84, 8),
56675 => conv_std_logic_vector(85, 8),
56676 => conv_std_logic_vector(86, 8),
56677 => conv_std_logic_vector(87, 8),
56678 => conv_std_logic_vector(88, 8),
56679 => conv_std_logic_vector(88, 8),
56680 => conv_std_logic_vector(89, 8),
56681 => conv_std_logic_vector(90, 8),
56682 => conv_std_logic_vector(91, 8),
56683 => conv_std_logic_vector(92, 8),
56684 => conv_std_logic_vector(93, 8),
56685 => conv_std_logic_vector(94, 8),
56686 => conv_std_logic_vector(94, 8),
56687 => conv_std_logic_vector(95, 8),
56688 => conv_std_logic_vector(96, 8),
56689 => conv_std_logic_vector(97, 8),
56690 => conv_std_logic_vector(98, 8),
56691 => conv_std_logic_vector(99, 8),
56692 => conv_std_logic_vector(100, 8),
56693 => conv_std_logic_vector(101, 8),
56694 => conv_std_logic_vector(101, 8),
56695 => conv_std_logic_vector(102, 8),
56696 => conv_std_logic_vector(103, 8),
56697 => conv_std_logic_vector(104, 8),
56698 => conv_std_logic_vector(105, 8),
56699 => conv_std_logic_vector(106, 8),
56700 => conv_std_logic_vector(107, 8),
56701 => conv_std_logic_vector(107, 8),
56702 => conv_std_logic_vector(108, 8),
56703 => conv_std_logic_vector(109, 8),
56704 => conv_std_logic_vector(110, 8),
56705 => conv_std_logic_vector(111, 8),
56706 => conv_std_logic_vector(112, 8),
56707 => conv_std_logic_vector(113, 8),
56708 => conv_std_logic_vector(113, 8),
56709 => conv_std_logic_vector(114, 8),
56710 => conv_std_logic_vector(115, 8),
56711 => conv_std_logic_vector(116, 8),
56712 => conv_std_logic_vector(117, 8),
56713 => conv_std_logic_vector(118, 8),
56714 => conv_std_logic_vector(119, 8),
56715 => conv_std_logic_vector(119, 8),
56716 => conv_std_logic_vector(120, 8),
56717 => conv_std_logic_vector(121, 8),
56718 => conv_std_logic_vector(122, 8),
56719 => conv_std_logic_vector(123, 8),
56720 => conv_std_logic_vector(124, 8),
56721 => conv_std_logic_vector(125, 8),
56722 => conv_std_logic_vector(126, 8),
56723 => conv_std_logic_vector(126, 8),
56724 => conv_std_logic_vector(127, 8),
56725 => conv_std_logic_vector(128, 8),
56726 => conv_std_logic_vector(129, 8),
56727 => conv_std_logic_vector(130, 8),
56728 => conv_std_logic_vector(131, 8),
56729 => conv_std_logic_vector(132, 8),
56730 => conv_std_logic_vector(132, 8),
56731 => conv_std_logic_vector(133, 8),
56732 => conv_std_logic_vector(134, 8),
56733 => conv_std_logic_vector(135, 8),
56734 => conv_std_logic_vector(136, 8),
56735 => conv_std_logic_vector(137, 8),
56736 => conv_std_logic_vector(138, 8),
56737 => conv_std_logic_vector(138, 8),
56738 => conv_std_logic_vector(139, 8),
56739 => conv_std_logic_vector(140, 8),
56740 => conv_std_logic_vector(141, 8),
56741 => conv_std_logic_vector(142, 8),
56742 => conv_std_logic_vector(143, 8),
56743 => conv_std_logic_vector(144, 8),
56744 => conv_std_logic_vector(145, 8),
56745 => conv_std_logic_vector(145, 8),
56746 => conv_std_logic_vector(146, 8),
56747 => conv_std_logic_vector(147, 8),
56748 => conv_std_logic_vector(148, 8),
56749 => conv_std_logic_vector(149, 8),
56750 => conv_std_logic_vector(150, 8),
56751 => conv_std_logic_vector(151, 8),
56752 => conv_std_logic_vector(151, 8),
56753 => conv_std_logic_vector(152, 8),
56754 => conv_std_logic_vector(153, 8),
56755 => conv_std_logic_vector(154, 8),
56756 => conv_std_logic_vector(155, 8),
56757 => conv_std_logic_vector(156, 8),
56758 => conv_std_logic_vector(157, 8),
56759 => conv_std_logic_vector(157, 8),
56760 => conv_std_logic_vector(158, 8),
56761 => conv_std_logic_vector(159, 8),
56762 => conv_std_logic_vector(160, 8),
56763 => conv_std_logic_vector(161, 8),
56764 => conv_std_logic_vector(162, 8),
56765 => conv_std_logic_vector(163, 8),
56766 => conv_std_logic_vector(164, 8),
56767 => conv_std_logic_vector(164, 8),
56768 => conv_std_logic_vector(165, 8),
56769 => conv_std_logic_vector(166, 8),
56770 => conv_std_logic_vector(167, 8),
56771 => conv_std_logic_vector(168, 8),
56772 => conv_std_logic_vector(169, 8),
56773 => conv_std_logic_vector(170, 8),
56774 => conv_std_logic_vector(170, 8),
56775 => conv_std_logic_vector(171, 8),
56776 => conv_std_logic_vector(172, 8),
56777 => conv_std_logic_vector(173, 8),
56778 => conv_std_logic_vector(174, 8),
56779 => conv_std_logic_vector(175, 8),
56780 => conv_std_logic_vector(176, 8),
56781 => conv_std_logic_vector(176, 8),
56782 => conv_std_logic_vector(177, 8),
56783 => conv_std_logic_vector(178, 8),
56784 => conv_std_logic_vector(179, 8),
56785 => conv_std_logic_vector(180, 8),
56786 => conv_std_logic_vector(181, 8),
56787 => conv_std_logic_vector(182, 8),
56788 => conv_std_logic_vector(183, 8),
56789 => conv_std_logic_vector(183, 8),
56790 => conv_std_logic_vector(184, 8),
56791 => conv_std_logic_vector(185, 8),
56792 => conv_std_logic_vector(186, 8),
56793 => conv_std_logic_vector(187, 8),
56794 => conv_std_logic_vector(188, 8),
56795 => conv_std_logic_vector(189, 8),
56796 => conv_std_logic_vector(189, 8),
56797 => conv_std_logic_vector(190, 8),
56798 => conv_std_logic_vector(191, 8),
56799 => conv_std_logic_vector(192, 8),
56800 => conv_std_logic_vector(193, 8),
56801 => conv_std_logic_vector(194, 8),
56802 => conv_std_logic_vector(195, 8),
56803 => conv_std_logic_vector(195, 8),
56804 => conv_std_logic_vector(196, 8),
56805 => conv_std_logic_vector(197, 8),
56806 => conv_std_logic_vector(198, 8),
56807 => conv_std_logic_vector(199, 8),
56808 => conv_std_logic_vector(200, 8),
56809 => conv_std_logic_vector(201, 8),
56810 => conv_std_logic_vector(202, 8),
56811 => conv_std_logic_vector(202, 8),
56812 => conv_std_logic_vector(203, 8),
56813 => conv_std_logic_vector(204, 8),
56814 => conv_std_logic_vector(205, 8),
56815 => conv_std_logic_vector(206, 8),
56816 => conv_std_logic_vector(207, 8),
56817 => conv_std_logic_vector(208, 8),
56818 => conv_std_logic_vector(208, 8),
56819 => conv_std_logic_vector(209, 8),
56820 => conv_std_logic_vector(210, 8),
56821 => conv_std_logic_vector(211, 8),
56822 => conv_std_logic_vector(212, 8),
56823 => conv_std_logic_vector(213, 8),
56824 => conv_std_logic_vector(214, 8),
56825 => conv_std_logic_vector(214, 8),
56826 => conv_std_logic_vector(215, 8),
56827 => conv_std_logic_vector(216, 8),
56828 => conv_std_logic_vector(217, 8),
56829 => conv_std_logic_vector(218, 8),
56830 => conv_std_logic_vector(219, 8),
56831 => conv_std_logic_vector(220, 8),
56832 => conv_std_logic_vector(0, 8),
56833 => conv_std_logic_vector(0, 8),
56834 => conv_std_logic_vector(1, 8),
56835 => conv_std_logic_vector(2, 8),
56836 => conv_std_logic_vector(3, 8),
56837 => conv_std_logic_vector(4, 8),
56838 => conv_std_logic_vector(5, 8),
56839 => conv_std_logic_vector(6, 8),
56840 => conv_std_logic_vector(6, 8),
56841 => conv_std_logic_vector(7, 8),
56842 => conv_std_logic_vector(8, 8),
56843 => conv_std_logic_vector(9, 8),
56844 => conv_std_logic_vector(10, 8),
56845 => conv_std_logic_vector(11, 8),
56846 => conv_std_logic_vector(12, 8),
56847 => conv_std_logic_vector(13, 8),
56848 => conv_std_logic_vector(13, 8),
56849 => conv_std_logic_vector(14, 8),
56850 => conv_std_logic_vector(15, 8),
56851 => conv_std_logic_vector(16, 8),
56852 => conv_std_logic_vector(17, 8),
56853 => conv_std_logic_vector(18, 8),
56854 => conv_std_logic_vector(19, 8),
56855 => conv_std_logic_vector(19, 8),
56856 => conv_std_logic_vector(20, 8),
56857 => conv_std_logic_vector(21, 8),
56858 => conv_std_logic_vector(22, 8),
56859 => conv_std_logic_vector(23, 8),
56860 => conv_std_logic_vector(24, 8),
56861 => conv_std_logic_vector(25, 8),
56862 => conv_std_logic_vector(26, 8),
56863 => conv_std_logic_vector(26, 8),
56864 => conv_std_logic_vector(27, 8),
56865 => conv_std_logic_vector(28, 8),
56866 => conv_std_logic_vector(29, 8),
56867 => conv_std_logic_vector(30, 8),
56868 => conv_std_logic_vector(31, 8),
56869 => conv_std_logic_vector(32, 8),
56870 => conv_std_logic_vector(32, 8),
56871 => conv_std_logic_vector(33, 8),
56872 => conv_std_logic_vector(34, 8),
56873 => conv_std_logic_vector(35, 8),
56874 => conv_std_logic_vector(36, 8),
56875 => conv_std_logic_vector(37, 8),
56876 => conv_std_logic_vector(38, 8),
56877 => conv_std_logic_vector(39, 8),
56878 => conv_std_logic_vector(39, 8),
56879 => conv_std_logic_vector(40, 8),
56880 => conv_std_logic_vector(41, 8),
56881 => conv_std_logic_vector(42, 8),
56882 => conv_std_logic_vector(43, 8),
56883 => conv_std_logic_vector(44, 8),
56884 => conv_std_logic_vector(45, 8),
56885 => conv_std_logic_vector(45, 8),
56886 => conv_std_logic_vector(46, 8),
56887 => conv_std_logic_vector(47, 8),
56888 => conv_std_logic_vector(48, 8),
56889 => conv_std_logic_vector(49, 8),
56890 => conv_std_logic_vector(50, 8),
56891 => conv_std_logic_vector(51, 8),
56892 => conv_std_logic_vector(52, 8),
56893 => conv_std_logic_vector(52, 8),
56894 => conv_std_logic_vector(53, 8),
56895 => conv_std_logic_vector(54, 8),
56896 => conv_std_logic_vector(55, 8),
56897 => conv_std_logic_vector(56, 8),
56898 => conv_std_logic_vector(57, 8),
56899 => conv_std_logic_vector(58, 8),
56900 => conv_std_logic_vector(58, 8),
56901 => conv_std_logic_vector(59, 8),
56902 => conv_std_logic_vector(60, 8),
56903 => conv_std_logic_vector(61, 8),
56904 => conv_std_logic_vector(62, 8),
56905 => conv_std_logic_vector(63, 8),
56906 => conv_std_logic_vector(64, 8),
56907 => conv_std_logic_vector(65, 8),
56908 => conv_std_logic_vector(65, 8),
56909 => conv_std_logic_vector(66, 8),
56910 => conv_std_logic_vector(67, 8),
56911 => conv_std_logic_vector(68, 8),
56912 => conv_std_logic_vector(69, 8),
56913 => conv_std_logic_vector(70, 8),
56914 => conv_std_logic_vector(71, 8),
56915 => conv_std_logic_vector(71, 8),
56916 => conv_std_logic_vector(72, 8),
56917 => conv_std_logic_vector(73, 8),
56918 => conv_std_logic_vector(74, 8),
56919 => conv_std_logic_vector(75, 8),
56920 => conv_std_logic_vector(76, 8),
56921 => conv_std_logic_vector(77, 8),
56922 => conv_std_logic_vector(78, 8),
56923 => conv_std_logic_vector(78, 8),
56924 => conv_std_logic_vector(79, 8),
56925 => conv_std_logic_vector(80, 8),
56926 => conv_std_logic_vector(81, 8),
56927 => conv_std_logic_vector(82, 8),
56928 => conv_std_logic_vector(83, 8),
56929 => conv_std_logic_vector(84, 8),
56930 => conv_std_logic_vector(84, 8),
56931 => conv_std_logic_vector(85, 8),
56932 => conv_std_logic_vector(86, 8),
56933 => conv_std_logic_vector(87, 8),
56934 => conv_std_logic_vector(88, 8),
56935 => conv_std_logic_vector(89, 8),
56936 => conv_std_logic_vector(90, 8),
56937 => conv_std_logic_vector(91, 8),
56938 => conv_std_logic_vector(91, 8),
56939 => conv_std_logic_vector(92, 8),
56940 => conv_std_logic_vector(93, 8),
56941 => conv_std_logic_vector(94, 8),
56942 => conv_std_logic_vector(95, 8),
56943 => conv_std_logic_vector(96, 8),
56944 => conv_std_logic_vector(97, 8),
56945 => conv_std_logic_vector(97, 8),
56946 => conv_std_logic_vector(98, 8),
56947 => conv_std_logic_vector(99, 8),
56948 => conv_std_logic_vector(100, 8),
56949 => conv_std_logic_vector(101, 8),
56950 => conv_std_logic_vector(102, 8),
56951 => conv_std_logic_vector(103, 8),
56952 => conv_std_logic_vector(104, 8),
56953 => conv_std_logic_vector(104, 8),
56954 => conv_std_logic_vector(105, 8),
56955 => conv_std_logic_vector(106, 8),
56956 => conv_std_logic_vector(107, 8),
56957 => conv_std_logic_vector(108, 8),
56958 => conv_std_logic_vector(109, 8),
56959 => conv_std_logic_vector(110, 8),
56960 => conv_std_logic_vector(111, 8),
56961 => conv_std_logic_vector(111, 8),
56962 => conv_std_logic_vector(112, 8),
56963 => conv_std_logic_vector(113, 8),
56964 => conv_std_logic_vector(114, 8),
56965 => conv_std_logic_vector(115, 8),
56966 => conv_std_logic_vector(116, 8),
56967 => conv_std_logic_vector(117, 8),
56968 => conv_std_logic_vector(117, 8),
56969 => conv_std_logic_vector(118, 8),
56970 => conv_std_logic_vector(119, 8),
56971 => conv_std_logic_vector(120, 8),
56972 => conv_std_logic_vector(121, 8),
56973 => conv_std_logic_vector(122, 8),
56974 => conv_std_logic_vector(123, 8),
56975 => conv_std_logic_vector(124, 8),
56976 => conv_std_logic_vector(124, 8),
56977 => conv_std_logic_vector(125, 8),
56978 => conv_std_logic_vector(126, 8),
56979 => conv_std_logic_vector(127, 8),
56980 => conv_std_logic_vector(128, 8),
56981 => conv_std_logic_vector(129, 8),
56982 => conv_std_logic_vector(130, 8),
56983 => conv_std_logic_vector(130, 8),
56984 => conv_std_logic_vector(131, 8),
56985 => conv_std_logic_vector(132, 8),
56986 => conv_std_logic_vector(133, 8),
56987 => conv_std_logic_vector(134, 8),
56988 => conv_std_logic_vector(135, 8),
56989 => conv_std_logic_vector(136, 8),
56990 => conv_std_logic_vector(137, 8),
56991 => conv_std_logic_vector(137, 8),
56992 => conv_std_logic_vector(138, 8),
56993 => conv_std_logic_vector(139, 8),
56994 => conv_std_logic_vector(140, 8),
56995 => conv_std_logic_vector(141, 8),
56996 => conv_std_logic_vector(142, 8),
56997 => conv_std_logic_vector(143, 8),
56998 => conv_std_logic_vector(143, 8),
56999 => conv_std_logic_vector(144, 8),
57000 => conv_std_logic_vector(145, 8),
57001 => conv_std_logic_vector(146, 8),
57002 => conv_std_logic_vector(147, 8),
57003 => conv_std_logic_vector(148, 8),
57004 => conv_std_logic_vector(149, 8),
57005 => conv_std_logic_vector(150, 8),
57006 => conv_std_logic_vector(150, 8),
57007 => conv_std_logic_vector(151, 8),
57008 => conv_std_logic_vector(152, 8),
57009 => conv_std_logic_vector(153, 8),
57010 => conv_std_logic_vector(154, 8),
57011 => conv_std_logic_vector(155, 8),
57012 => conv_std_logic_vector(156, 8),
57013 => conv_std_logic_vector(156, 8),
57014 => conv_std_logic_vector(157, 8),
57015 => conv_std_logic_vector(158, 8),
57016 => conv_std_logic_vector(159, 8),
57017 => conv_std_logic_vector(160, 8),
57018 => conv_std_logic_vector(161, 8),
57019 => conv_std_logic_vector(162, 8),
57020 => conv_std_logic_vector(163, 8),
57021 => conv_std_logic_vector(163, 8),
57022 => conv_std_logic_vector(164, 8),
57023 => conv_std_logic_vector(165, 8),
57024 => conv_std_logic_vector(166, 8),
57025 => conv_std_logic_vector(167, 8),
57026 => conv_std_logic_vector(168, 8),
57027 => conv_std_logic_vector(169, 8),
57028 => conv_std_logic_vector(169, 8),
57029 => conv_std_logic_vector(170, 8),
57030 => conv_std_logic_vector(171, 8),
57031 => conv_std_logic_vector(172, 8),
57032 => conv_std_logic_vector(173, 8),
57033 => conv_std_logic_vector(174, 8),
57034 => conv_std_logic_vector(175, 8),
57035 => conv_std_logic_vector(176, 8),
57036 => conv_std_logic_vector(176, 8),
57037 => conv_std_logic_vector(177, 8),
57038 => conv_std_logic_vector(178, 8),
57039 => conv_std_logic_vector(179, 8),
57040 => conv_std_logic_vector(180, 8),
57041 => conv_std_logic_vector(181, 8),
57042 => conv_std_logic_vector(182, 8),
57043 => conv_std_logic_vector(182, 8),
57044 => conv_std_logic_vector(183, 8),
57045 => conv_std_logic_vector(184, 8),
57046 => conv_std_logic_vector(185, 8),
57047 => conv_std_logic_vector(186, 8),
57048 => conv_std_logic_vector(187, 8),
57049 => conv_std_logic_vector(188, 8),
57050 => conv_std_logic_vector(189, 8),
57051 => conv_std_logic_vector(189, 8),
57052 => conv_std_logic_vector(190, 8),
57053 => conv_std_logic_vector(191, 8),
57054 => conv_std_logic_vector(192, 8),
57055 => conv_std_logic_vector(193, 8),
57056 => conv_std_logic_vector(194, 8),
57057 => conv_std_logic_vector(195, 8),
57058 => conv_std_logic_vector(195, 8),
57059 => conv_std_logic_vector(196, 8),
57060 => conv_std_logic_vector(197, 8),
57061 => conv_std_logic_vector(198, 8),
57062 => conv_std_logic_vector(199, 8),
57063 => conv_std_logic_vector(200, 8),
57064 => conv_std_logic_vector(201, 8),
57065 => conv_std_logic_vector(202, 8),
57066 => conv_std_logic_vector(202, 8),
57067 => conv_std_logic_vector(203, 8),
57068 => conv_std_logic_vector(204, 8),
57069 => conv_std_logic_vector(205, 8),
57070 => conv_std_logic_vector(206, 8),
57071 => conv_std_logic_vector(207, 8),
57072 => conv_std_logic_vector(208, 8),
57073 => conv_std_logic_vector(208, 8),
57074 => conv_std_logic_vector(209, 8),
57075 => conv_std_logic_vector(210, 8),
57076 => conv_std_logic_vector(211, 8),
57077 => conv_std_logic_vector(212, 8),
57078 => conv_std_logic_vector(213, 8),
57079 => conv_std_logic_vector(214, 8),
57080 => conv_std_logic_vector(215, 8),
57081 => conv_std_logic_vector(215, 8),
57082 => conv_std_logic_vector(216, 8),
57083 => conv_std_logic_vector(217, 8),
57084 => conv_std_logic_vector(218, 8),
57085 => conv_std_logic_vector(219, 8),
57086 => conv_std_logic_vector(220, 8),
57087 => conv_std_logic_vector(221, 8),
57088 => conv_std_logic_vector(0, 8),
57089 => conv_std_logic_vector(0, 8),
57090 => conv_std_logic_vector(1, 8),
57091 => conv_std_logic_vector(2, 8),
57092 => conv_std_logic_vector(3, 8),
57093 => conv_std_logic_vector(4, 8),
57094 => conv_std_logic_vector(5, 8),
57095 => conv_std_logic_vector(6, 8),
57096 => conv_std_logic_vector(6, 8),
57097 => conv_std_logic_vector(7, 8),
57098 => conv_std_logic_vector(8, 8),
57099 => conv_std_logic_vector(9, 8),
57100 => conv_std_logic_vector(10, 8),
57101 => conv_std_logic_vector(11, 8),
57102 => conv_std_logic_vector(12, 8),
57103 => conv_std_logic_vector(13, 8),
57104 => conv_std_logic_vector(13, 8),
57105 => conv_std_logic_vector(14, 8),
57106 => conv_std_logic_vector(15, 8),
57107 => conv_std_logic_vector(16, 8),
57108 => conv_std_logic_vector(17, 8),
57109 => conv_std_logic_vector(18, 8),
57110 => conv_std_logic_vector(19, 8),
57111 => conv_std_logic_vector(20, 8),
57112 => conv_std_logic_vector(20, 8),
57113 => conv_std_logic_vector(21, 8),
57114 => conv_std_logic_vector(22, 8),
57115 => conv_std_logic_vector(23, 8),
57116 => conv_std_logic_vector(24, 8),
57117 => conv_std_logic_vector(25, 8),
57118 => conv_std_logic_vector(26, 8),
57119 => conv_std_logic_vector(27, 8),
57120 => conv_std_logic_vector(27, 8),
57121 => conv_std_logic_vector(28, 8),
57122 => conv_std_logic_vector(29, 8),
57123 => conv_std_logic_vector(30, 8),
57124 => conv_std_logic_vector(31, 8),
57125 => conv_std_logic_vector(32, 8),
57126 => conv_std_logic_vector(33, 8),
57127 => conv_std_logic_vector(33, 8),
57128 => conv_std_logic_vector(34, 8),
57129 => conv_std_logic_vector(35, 8),
57130 => conv_std_logic_vector(36, 8),
57131 => conv_std_logic_vector(37, 8),
57132 => conv_std_logic_vector(38, 8),
57133 => conv_std_logic_vector(39, 8),
57134 => conv_std_logic_vector(40, 8),
57135 => conv_std_logic_vector(40, 8),
57136 => conv_std_logic_vector(41, 8),
57137 => conv_std_logic_vector(42, 8),
57138 => conv_std_logic_vector(43, 8),
57139 => conv_std_logic_vector(44, 8),
57140 => conv_std_logic_vector(45, 8),
57141 => conv_std_logic_vector(46, 8),
57142 => conv_std_logic_vector(47, 8),
57143 => conv_std_logic_vector(47, 8),
57144 => conv_std_logic_vector(48, 8),
57145 => conv_std_logic_vector(49, 8),
57146 => conv_std_logic_vector(50, 8),
57147 => conv_std_logic_vector(51, 8),
57148 => conv_std_logic_vector(52, 8),
57149 => conv_std_logic_vector(53, 8),
57150 => conv_std_logic_vector(54, 8),
57151 => conv_std_logic_vector(54, 8),
57152 => conv_std_logic_vector(55, 8),
57153 => conv_std_logic_vector(56, 8),
57154 => conv_std_logic_vector(57, 8),
57155 => conv_std_logic_vector(58, 8),
57156 => conv_std_logic_vector(59, 8),
57157 => conv_std_logic_vector(60, 8),
57158 => conv_std_logic_vector(60, 8),
57159 => conv_std_logic_vector(61, 8),
57160 => conv_std_logic_vector(62, 8),
57161 => conv_std_logic_vector(63, 8),
57162 => conv_std_logic_vector(64, 8),
57163 => conv_std_logic_vector(65, 8),
57164 => conv_std_logic_vector(66, 8),
57165 => conv_std_logic_vector(67, 8),
57166 => conv_std_logic_vector(67, 8),
57167 => conv_std_logic_vector(68, 8),
57168 => conv_std_logic_vector(69, 8),
57169 => conv_std_logic_vector(70, 8),
57170 => conv_std_logic_vector(71, 8),
57171 => conv_std_logic_vector(72, 8),
57172 => conv_std_logic_vector(73, 8),
57173 => conv_std_logic_vector(74, 8),
57174 => conv_std_logic_vector(74, 8),
57175 => conv_std_logic_vector(75, 8),
57176 => conv_std_logic_vector(76, 8),
57177 => conv_std_logic_vector(77, 8),
57178 => conv_std_logic_vector(78, 8),
57179 => conv_std_logic_vector(79, 8),
57180 => conv_std_logic_vector(80, 8),
57181 => conv_std_logic_vector(81, 8),
57182 => conv_std_logic_vector(81, 8),
57183 => conv_std_logic_vector(82, 8),
57184 => conv_std_logic_vector(83, 8),
57185 => conv_std_logic_vector(84, 8),
57186 => conv_std_logic_vector(85, 8),
57187 => conv_std_logic_vector(86, 8),
57188 => conv_std_logic_vector(87, 8),
57189 => conv_std_logic_vector(87, 8),
57190 => conv_std_logic_vector(88, 8),
57191 => conv_std_logic_vector(89, 8),
57192 => conv_std_logic_vector(90, 8),
57193 => conv_std_logic_vector(91, 8),
57194 => conv_std_logic_vector(92, 8),
57195 => conv_std_logic_vector(93, 8),
57196 => conv_std_logic_vector(94, 8),
57197 => conv_std_logic_vector(94, 8),
57198 => conv_std_logic_vector(95, 8),
57199 => conv_std_logic_vector(96, 8),
57200 => conv_std_logic_vector(97, 8),
57201 => conv_std_logic_vector(98, 8),
57202 => conv_std_logic_vector(99, 8),
57203 => conv_std_logic_vector(100, 8),
57204 => conv_std_logic_vector(101, 8),
57205 => conv_std_logic_vector(101, 8),
57206 => conv_std_logic_vector(102, 8),
57207 => conv_std_logic_vector(103, 8),
57208 => conv_std_logic_vector(104, 8),
57209 => conv_std_logic_vector(105, 8),
57210 => conv_std_logic_vector(106, 8),
57211 => conv_std_logic_vector(107, 8),
57212 => conv_std_logic_vector(108, 8),
57213 => conv_std_logic_vector(108, 8),
57214 => conv_std_logic_vector(109, 8),
57215 => conv_std_logic_vector(110, 8),
57216 => conv_std_logic_vector(111, 8),
57217 => conv_std_logic_vector(112, 8),
57218 => conv_std_logic_vector(113, 8),
57219 => conv_std_logic_vector(114, 8),
57220 => conv_std_logic_vector(114, 8),
57221 => conv_std_logic_vector(115, 8),
57222 => conv_std_logic_vector(116, 8),
57223 => conv_std_logic_vector(117, 8),
57224 => conv_std_logic_vector(118, 8),
57225 => conv_std_logic_vector(119, 8),
57226 => conv_std_logic_vector(120, 8),
57227 => conv_std_logic_vector(121, 8),
57228 => conv_std_logic_vector(121, 8),
57229 => conv_std_logic_vector(122, 8),
57230 => conv_std_logic_vector(123, 8),
57231 => conv_std_logic_vector(124, 8),
57232 => conv_std_logic_vector(125, 8),
57233 => conv_std_logic_vector(126, 8),
57234 => conv_std_logic_vector(127, 8),
57235 => conv_std_logic_vector(128, 8),
57236 => conv_std_logic_vector(128, 8),
57237 => conv_std_logic_vector(129, 8),
57238 => conv_std_logic_vector(130, 8),
57239 => conv_std_logic_vector(131, 8),
57240 => conv_std_logic_vector(132, 8),
57241 => conv_std_logic_vector(133, 8),
57242 => conv_std_logic_vector(134, 8),
57243 => conv_std_logic_vector(135, 8),
57244 => conv_std_logic_vector(135, 8),
57245 => conv_std_logic_vector(136, 8),
57246 => conv_std_logic_vector(137, 8),
57247 => conv_std_logic_vector(138, 8),
57248 => conv_std_logic_vector(139, 8),
57249 => conv_std_logic_vector(140, 8),
57250 => conv_std_logic_vector(141, 8),
57251 => conv_std_logic_vector(141, 8),
57252 => conv_std_logic_vector(142, 8),
57253 => conv_std_logic_vector(143, 8),
57254 => conv_std_logic_vector(144, 8),
57255 => conv_std_logic_vector(145, 8),
57256 => conv_std_logic_vector(146, 8),
57257 => conv_std_logic_vector(147, 8),
57258 => conv_std_logic_vector(148, 8),
57259 => conv_std_logic_vector(148, 8),
57260 => conv_std_logic_vector(149, 8),
57261 => conv_std_logic_vector(150, 8),
57262 => conv_std_logic_vector(151, 8),
57263 => conv_std_logic_vector(152, 8),
57264 => conv_std_logic_vector(153, 8),
57265 => conv_std_logic_vector(154, 8),
57266 => conv_std_logic_vector(155, 8),
57267 => conv_std_logic_vector(155, 8),
57268 => conv_std_logic_vector(156, 8),
57269 => conv_std_logic_vector(157, 8),
57270 => conv_std_logic_vector(158, 8),
57271 => conv_std_logic_vector(159, 8),
57272 => conv_std_logic_vector(160, 8),
57273 => conv_std_logic_vector(161, 8),
57274 => conv_std_logic_vector(162, 8),
57275 => conv_std_logic_vector(162, 8),
57276 => conv_std_logic_vector(163, 8),
57277 => conv_std_logic_vector(164, 8),
57278 => conv_std_logic_vector(165, 8),
57279 => conv_std_logic_vector(166, 8),
57280 => conv_std_logic_vector(167, 8),
57281 => conv_std_logic_vector(168, 8),
57282 => conv_std_logic_vector(168, 8),
57283 => conv_std_logic_vector(169, 8),
57284 => conv_std_logic_vector(170, 8),
57285 => conv_std_logic_vector(171, 8),
57286 => conv_std_logic_vector(172, 8),
57287 => conv_std_logic_vector(173, 8),
57288 => conv_std_logic_vector(174, 8),
57289 => conv_std_logic_vector(175, 8),
57290 => conv_std_logic_vector(175, 8),
57291 => conv_std_logic_vector(176, 8),
57292 => conv_std_logic_vector(177, 8),
57293 => conv_std_logic_vector(178, 8),
57294 => conv_std_logic_vector(179, 8),
57295 => conv_std_logic_vector(180, 8),
57296 => conv_std_logic_vector(181, 8),
57297 => conv_std_logic_vector(182, 8),
57298 => conv_std_logic_vector(182, 8),
57299 => conv_std_logic_vector(183, 8),
57300 => conv_std_logic_vector(184, 8),
57301 => conv_std_logic_vector(185, 8),
57302 => conv_std_logic_vector(186, 8),
57303 => conv_std_logic_vector(187, 8),
57304 => conv_std_logic_vector(188, 8),
57305 => conv_std_logic_vector(189, 8),
57306 => conv_std_logic_vector(189, 8),
57307 => conv_std_logic_vector(190, 8),
57308 => conv_std_logic_vector(191, 8),
57309 => conv_std_logic_vector(192, 8),
57310 => conv_std_logic_vector(193, 8),
57311 => conv_std_logic_vector(194, 8),
57312 => conv_std_logic_vector(195, 8),
57313 => conv_std_logic_vector(195, 8),
57314 => conv_std_logic_vector(196, 8),
57315 => conv_std_logic_vector(197, 8),
57316 => conv_std_logic_vector(198, 8),
57317 => conv_std_logic_vector(199, 8),
57318 => conv_std_logic_vector(200, 8),
57319 => conv_std_logic_vector(201, 8),
57320 => conv_std_logic_vector(202, 8),
57321 => conv_std_logic_vector(202, 8),
57322 => conv_std_logic_vector(203, 8),
57323 => conv_std_logic_vector(204, 8),
57324 => conv_std_logic_vector(205, 8),
57325 => conv_std_logic_vector(206, 8),
57326 => conv_std_logic_vector(207, 8),
57327 => conv_std_logic_vector(208, 8),
57328 => conv_std_logic_vector(209, 8),
57329 => conv_std_logic_vector(209, 8),
57330 => conv_std_logic_vector(210, 8),
57331 => conv_std_logic_vector(211, 8),
57332 => conv_std_logic_vector(212, 8),
57333 => conv_std_logic_vector(213, 8),
57334 => conv_std_logic_vector(214, 8),
57335 => conv_std_logic_vector(215, 8),
57336 => conv_std_logic_vector(216, 8),
57337 => conv_std_logic_vector(216, 8),
57338 => conv_std_logic_vector(217, 8),
57339 => conv_std_logic_vector(218, 8),
57340 => conv_std_logic_vector(219, 8),
57341 => conv_std_logic_vector(220, 8),
57342 => conv_std_logic_vector(221, 8),
57343 => conv_std_logic_vector(222, 8),
57344 => conv_std_logic_vector(0, 8),
57345 => conv_std_logic_vector(0, 8),
57346 => conv_std_logic_vector(1, 8),
57347 => conv_std_logic_vector(2, 8),
57348 => conv_std_logic_vector(3, 8),
57349 => conv_std_logic_vector(4, 8),
57350 => conv_std_logic_vector(5, 8),
57351 => conv_std_logic_vector(6, 8),
57352 => conv_std_logic_vector(7, 8),
57353 => conv_std_logic_vector(7, 8),
57354 => conv_std_logic_vector(8, 8),
57355 => conv_std_logic_vector(9, 8),
57356 => conv_std_logic_vector(10, 8),
57357 => conv_std_logic_vector(11, 8),
57358 => conv_std_logic_vector(12, 8),
57359 => conv_std_logic_vector(13, 8),
57360 => conv_std_logic_vector(14, 8),
57361 => conv_std_logic_vector(14, 8),
57362 => conv_std_logic_vector(15, 8),
57363 => conv_std_logic_vector(16, 8),
57364 => conv_std_logic_vector(17, 8),
57365 => conv_std_logic_vector(18, 8),
57366 => conv_std_logic_vector(19, 8),
57367 => conv_std_logic_vector(20, 8),
57368 => conv_std_logic_vector(21, 8),
57369 => conv_std_logic_vector(21, 8),
57370 => conv_std_logic_vector(22, 8),
57371 => conv_std_logic_vector(23, 8),
57372 => conv_std_logic_vector(24, 8),
57373 => conv_std_logic_vector(25, 8),
57374 => conv_std_logic_vector(26, 8),
57375 => conv_std_logic_vector(27, 8),
57376 => conv_std_logic_vector(28, 8),
57377 => conv_std_logic_vector(28, 8),
57378 => conv_std_logic_vector(29, 8),
57379 => conv_std_logic_vector(30, 8),
57380 => conv_std_logic_vector(31, 8),
57381 => conv_std_logic_vector(32, 8),
57382 => conv_std_logic_vector(33, 8),
57383 => conv_std_logic_vector(34, 8),
57384 => conv_std_logic_vector(35, 8),
57385 => conv_std_logic_vector(35, 8),
57386 => conv_std_logic_vector(36, 8),
57387 => conv_std_logic_vector(37, 8),
57388 => conv_std_logic_vector(38, 8),
57389 => conv_std_logic_vector(39, 8),
57390 => conv_std_logic_vector(40, 8),
57391 => conv_std_logic_vector(41, 8),
57392 => conv_std_logic_vector(42, 8),
57393 => conv_std_logic_vector(42, 8),
57394 => conv_std_logic_vector(43, 8),
57395 => conv_std_logic_vector(44, 8),
57396 => conv_std_logic_vector(45, 8),
57397 => conv_std_logic_vector(46, 8),
57398 => conv_std_logic_vector(47, 8),
57399 => conv_std_logic_vector(48, 8),
57400 => conv_std_logic_vector(49, 8),
57401 => conv_std_logic_vector(49, 8),
57402 => conv_std_logic_vector(50, 8),
57403 => conv_std_logic_vector(51, 8),
57404 => conv_std_logic_vector(52, 8),
57405 => conv_std_logic_vector(53, 8),
57406 => conv_std_logic_vector(54, 8),
57407 => conv_std_logic_vector(55, 8),
57408 => conv_std_logic_vector(56, 8),
57409 => conv_std_logic_vector(56, 8),
57410 => conv_std_logic_vector(57, 8),
57411 => conv_std_logic_vector(58, 8),
57412 => conv_std_logic_vector(59, 8),
57413 => conv_std_logic_vector(60, 8),
57414 => conv_std_logic_vector(61, 8),
57415 => conv_std_logic_vector(62, 8),
57416 => conv_std_logic_vector(63, 8),
57417 => conv_std_logic_vector(63, 8),
57418 => conv_std_logic_vector(64, 8),
57419 => conv_std_logic_vector(65, 8),
57420 => conv_std_logic_vector(66, 8),
57421 => conv_std_logic_vector(67, 8),
57422 => conv_std_logic_vector(68, 8),
57423 => conv_std_logic_vector(69, 8),
57424 => conv_std_logic_vector(70, 8),
57425 => conv_std_logic_vector(70, 8),
57426 => conv_std_logic_vector(71, 8),
57427 => conv_std_logic_vector(72, 8),
57428 => conv_std_logic_vector(73, 8),
57429 => conv_std_logic_vector(74, 8),
57430 => conv_std_logic_vector(75, 8),
57431 => conv_std_logic_vector(76, 8),
57432 => conv_std_logic_vector(77, 8),
57433 => conv_std_logic_vector(77, 8),
57434 => conv_std_logic_vector(78, 8),
57435 => conv_std_logic_vector(79, 8),
57436 => conv_std_logic_vector(80, 8),
57437 => conv_std_logic_vector(81, 8),
57438 => conv_std_logic_vector(82, 8),
57439 => conv_std_logic_vector(83, 8),
57440 => conv_std_logic_vector(84, 8),
57441 => conv_std_logic_vector(84, 8),
57442 => conv_std_logic_vector(85, 8),
57443 => conv_std_logic_vector(86, 8),
57444 => conv_std_logic_vector(87, 8),
57445 => conv_std_logic_vector(88, 8),
57446 => conv_std_logic_vector(89, 8),
57447 => conv_std_logic_vector(90, 8),
57448 => conv_std_logic_vector(91, 8),
57449 => conv_std_logic_vector(91, 8),
57450 => conv_std_logic_vector(92, 8),
57451 => conv_std_logic_vector(93, 8),
57452 => conv_std_logic_vector(94, 8),
57453 => conv_std_logic_vector(95, 8),
57454 => conv_std_logic_vector(96, 8),
57455 => conv_std_logic_vector(97, 8),
57456 => conv_std_logic_vector(98, 8),
57457 => conv_std_logic_vector(98, 8),
57458 => conv_std_logic_vector(99, 8),
57459 => conv_std_logic_vector(100, 8),
57460 => conv_std_logic_vector(101, 8),
57461 => conv_std_logic_vector(102, 8),
57462 => conv_std_logic_vector(103, 8),
57463 => conv_std_logic_vector(104, 8),
57464 => conv_std_logic_vector(105, 8),
57465 => conv_std_logic_vector(105, 8),
57466 => conv_std_logic_vector(106, 8),
57467 => conv_std_logic_vector(107, 8),
57468 => conv_std_logic_vector(108, 8),
57469 => conv_std_logic_vector(109, 8),
57470 => conv_std_logic_vector(110, 8),
57471 => conv_std_logic_vector(111, 8),
57472 => conv_std_logic_vector(112, 8),
57473 => conv_std_logic_vector(112, 8),
57474 => conv_std_logic_vector(113, 8),
57475 => conv_std_logic_vector(114, 8),
57476 => conv_std_logic_vector(115, 8),
57477 => conv_std_logic_vector(116, 8),
57478 => conv_std_logic_vector(117, 8),
57479 => conv_std_logic_vector(118, 8),
57480 => conv_std_logic_vector(119, 8),
57481 => conv_std_logic_vector(119, 8),
57482 => conv_std_logic_vector(120, 8),
57483 => conv_std_logic_vector(121, 8),
57484 => conv_std_logic_vector(122, 8),
57485 => conv_std_logic_vector(123, 8),
57486 => conv_std_logic_vector(124, 8),
57487 => conv_std_logic_vector(125, 8),
57488 => conv_std_logic_vector(126, 8),
57489 => conv_std_logic_vector(126, 8),
57490 => conv_std_logic_vector(127, 8),
57491 => conv_std_logic_vector(128, 8),
57492 => conv_std_logic_vector(129, 8),
57493 => conv_std_logic_vector(130, 8),
57494 => conv_std_logic_vector(131, 8),
57495 => conv_std_logic_vector(132, 8),
57496 => conv_std_logic_vector(133, 8),
57497 => conv_std_logic_vector(133, 8),
57498 => conv_std_logic_vector(134, 8),
57499 => conv_std_logic_vector(135, 8),
57500 => conv_std_logic_vector(136, 8),
57501 => conv_std_logic_vector(137, 8),
57502 => conv_std_logic_vector(138, 8),
57503 => conv_std_logic_vector(139, 8),
57504 => conv_std_logic_vector(140, 8),
57505 => conv_std_logic_vector(140, 8),
57506 => conv_std_logic_vector(141, 8),
57507 => conv_std_logic_vector(142, 8),
57508 => conv_std_logic_vector(143, 8),
57509 => conv_std_logic_vector(144, 8),
57510 => conv_std_logic_vector(145, 8),
57511 => conv_std_logic_vector(146, 8),
57512 => conv_std_logic_vector(147, 8),
57513 => conv_std_logic_vector(147, 8),
57514 => conv_std_logic_vector(148, 8),
57515 => conv_std_logic_vector(149, 8),
57516 => conv_std_logic_vector(150, 8),
57517 => conv_std_logic_vector(151, 8),
57518 => conv_std_logic_vector(152, 8),
57519 => conv_std_logic_vector(153, 8),
57520 => conv_std_logic_vector(154, 8),
57521 => conv_std_logic_vector(154, 8),
57522 => conv_std_logic_vector(155, 8),
57523 => conv_std_logic_vector(156, 8),
57524 => conv_std_logic_vector(157, 8),
57525 => conv_std_logic_vector(158, 8),
57526 => conv_std_logic_vector(159, 8),
57527 => conv_std_logic_vector(160, 8),
57528 => conv_std_logic_vector(161, 8),
57529 => conv_std_logic_vector(161, 8),
57530 => conv_std_logic_vector(162, 8),
57531 => conv_std_logic_vector(163, 8),
57532 => conv_std_logic_vector(164, 8),
57533 => conv_std_logic_vector(165, 8),
57534 => conv_std_logic_vector(166, 8),
57535 => conv_std_logic_vector(167, 8),
57536 => conv_std_logic_vector(168, 8),
57537 => conv_std_logic_vector(168, 8),
57538 => conv_std_logic_vector(169, 8),
57539 => conv_std_logic_vector(170, 8),
57540 => conv_std_logic_vector(171, 8),
57541 => conv_std_logic_vector(172, 8),
57542 => conv_std_logic_vector(173, 8),
57543 => conv_std_logic_vector(174, 8),
57544 => conv_std_logic_vector(175, 8),
57545 => conv_std_logic_vector(175, 8),
57546 => conv_std_logic_vector(176, 8),
57547 => conv_std_logic_vector(177, 8),
57548 => conv_std_logic_vector(178, 8),
57549 => conv_std_logic_vector(179, 8),
57550 => conv_std_logic_vector(180, 8),
57551 => conv_std_logic_vector(181, 8),
57552 => conv_std_logic_vector(182, 8),
57553 => conv_std_logic_vector(182, 8),
57554 => conv_std_logic_vector(183, 8),
57555 => conv_std_logic_vector(184, 8),
57556 => conv_std_logic_vector(185, 8),
57557 => conv_std_logic_vector(186, 8),
57558 => conv_std_logic_vector(187, 8),
57559 => conv_std_logic_vector(188, 8),
57560 => conv_std_logic_vector(189, 8),
57561 => conv_std_logic_vector(189, 8),
57562 => conv_std_logic_vector(190, 8),
57563 => conv_std_logic_vector(191, 8),
57564 => conv_std_logic_vector(192, 8),
57565 => conv_std_logic_vector(193, 8),
57566 => conv_std_logic_vector(194, 8),
57567 => conv_std_logic_vector(195, 8),
57568 => conv_std_logic_vector(196, 8),
57569 => conv_std_logic_vector(196, 8),
57570 => conv_std_logic_vector(197, 8),
57571 => conv_std_logic_vector(198, 8),
57572 => conv_std_logic_vector(199, 8),
57573 => conv_std_logic_vector(200, 8),
57574 => conv_std_logic_vector(201, 8),
57575 => conv_std_logic_vector(202, 8),
57576 => conv_std_logic_vector(203, 8),
57577 => conv_std_logic_vector(203, 8),
57578 => conv_std_logic_vector(204, 8),
57579 => conv_std_logic_vector(205, 8),
57580 => conv_std_logic_vector(206, 8),
57581 => conv_std_logic_vector(207, 8),
57582 => conv_std_logic_vector(208, 8),
57583 => conv_std_logic_vector(209, 8),
57584 => conv_std_logic_vector(210, 8),
57585 => conv_std_logic_vector(210, 8),
57586 => conv_std_logic_vector(211, 8),
57587 => conv_std_logic_vector(212, 8),
57588 => conv_std_logic_vector(213, 8),
57589 => conv_std_logic_vector(214, 8),
57590 => conv_std_logic_vector(215, 8),
57591 => conv_std_logic_vector(216, 8),
57592 => conv_std_logic_vector(217, 8),
57593 => conv_std_logic_vector(217, 8),
57594 => conv_std_logic_vector(218, 8),
57595 => conv_std_logic_vector(219, 8),
57596 => conv_std_logic_vector(220, 8),
57597 => conv_std_logic_vector(221, 8),
57598 => conv_std_logic_vector(222, 8),
57599 => conv_std_logic_vector(223, 8),
57600 => conv_std_logic_vector(0, 8),
57601 => conv_std_logic_vector(0, 8),
57602 => conv_std_logic_vector(1, 8),
57603 => conv_std_logic_vector(2, 8),
57604 => conv_std_logic_vector(3, 8),
57605 => conv_std_logic_vector(4, 8),
57606 => conv_std_logic_vector(5, 8),
57607 => conv_std_logic_vector(6, 8),
57608 => conv_std_logic_vector(7, 8),
57609 => conv_std_logic_vector(7, 8),
57610 => conv_std_logic_vector(8, 8),
57611 => conv_std_logic_vector(9, 8),
57612 => conv_std_logic_vector(10, 8),
57613 => conv_std_logic_vector(11, 8),
57614 => conv_std_logic_vector(12, 8),
57615 => conv_std_logic_vector(13, 8),
57616 => conv_std_logic_vector(14, 8),
57617 => conv_std_logic_vector(14, 8),
57618 => conv_std_logic_vector(15, 8),
57619 => conv_std_logic_vector(16, 8),
57620 => conv_std_logic_vector(17, 8),
57621 => conv_std_logic_vector(18, 8),
57622 => conv_std_logic_vector(19, 8),
57623 => conv_std_logic_vector(20, 8),
57624 => conv_std_logic_vector(21, 8),
57625 => conv_std_logic_vector(21, 8),
57626 => conv_std_logic_vector(22, 8),
57627 => conv_std_logic_vector(23, 8),
57628 => conv_std_logic_vector(24, 8),
57629 => conv_std_logic_vector(25, 8),
57630 => conv_std_logic_vector(26, 8),
57631 => conv_std_logic_vector(27, 8),
57632 => conv_std_logic_vector(28, 8),
57633 => conv_std_logic_vector(29, 8),
57634 => conv_std_logic_vector(29, 8),
57635 => conv_std_logic_vector(30, 8),
57636 => conv_std_logic_vector(31, 8),
57637 => conv_std_logic_vector(32, 8),
57638 => conv_std_logic_vector(33, 8),
57639 => conv_std_logic_vector(34, 8),
57640 => conv_std_logic_vector(35, 8),
57641 => conv_std_logic_vector(36, 8),
57642 => conv_std_logic_vector(36, 8),
57643 => conv_std_logic_vector(37, 8),
57644 => conv_std_logic_vector(38, 8),
57645 => conv_std_logic_vector(39, 8),
57646 => conv_std_logic_vector(40, 8),
57647 => conv_std_logic_vector(41, 8),
57648 => conv_std_logic_vector(42, 8),
57649 => conv_std_logic_vector(43, 8),
57650 => conv_std_logic_vector(43, 8),
57651 => conv_std_logic_vector(44, 8),
57652 => conv_std_logic_vector(45, 8),
57653 => conv_std_logic_vector(46, 8),
57654 => conv_std_logic_vector(47, 8),
57655 => conv_std_logic_vector(48, 8),
57656 => conv_std_logic_vector(49, 8),
57657 => conv_std_logic_vector(50, 8),
57658 => conv_std_logic_vector(50, 8),
57659 => conv_std_logic_vector(51, 8),
57660 => conv_std_logic_vector(52, 8),
57661 => conv_std_logic_vector(53, 8),
57662 => conv_std_logic_vector(54, 8),
57663 => conv_std_logic_vector(55, 8),
57664 => conv_std_logic_vector(56, 8),
57665 => conv_std_logic_vector(57, 8),
57666 => conv_std_logic_vector(58, 8),
57667 => conv_std_logic_vector(58, 8),
57668 => conv_std_logic_vector(59, 8),
57669 => conv_std_logic_vector(60, 8),
57670 => conv_std_logic_vector(61, 8),
57671 => conv_std_logic_vector(62, 8),
57672 => conv_std_logic_vector(63, 8),
57673 => conv_std_logic_vector(64, 8),
57674 => conv_std_logic_vector(65, 8),
57675 => conv_std_logic_vector(65, 8),
57676 => conv_std_logic_vector(66, 8),
57677 => conv_std_logic_vector(67, 8),
57678 => conv_std_logic_vector(68, 8),
57679 => conv_std_logic_vector(69, 8),
57680 => conv_std_logic_vector(70, 8),
57681 => conv_std_logic_vector(71, 8),
57682 => conv_std_logic_vector(72, 8),
57683 => conv_std_logic_vector(72, 8),
57684 => conv_std_logic_vector(73, 8),
57685 => conv_std_logic_vector(74, 8),
57686 => conv_std_logic_vector(75, 8),
57687 => conv_std_logic_vector(76, 8),
57688 => conv_std_logic_vector(77, 8),
57689 => conv_std_logic_vector(78, 8),
57690 => conv_std_logic_vector(79, 8),
57691 => conv_std_logic_vector(79, 8),
57692 => conv_std_logic_vector(80, 8),
57693 => conv_std_logic_vector(81, 8),
57694 => conv_std_logic_vector(82, 8),
57695 => conv_std_logic_vector(83, 8),
57696 => conv_std_logic_vector(84, 8),
57697 => conv_std_logic_vector(85, 8),
57698 => conv_std_logic_vector(86, 8),
57699 => conv_std_logic_vector(87, 8),
57700 => conv_std_logic_vector(87, 8),
57701 => conv_std_logic_vector(88, 8),
57702 => conv_std_logic_vector(89, 8),
57703 => conv_std_logic_vector(90, 8),
57704 => conv_std_logic_vector(91, 8),
57705 => conv_std_logic_vector(92, 8),
57706 => conv_std_logic_vector(93, 8),
57707 => conv_std_logic_vector(94, 8),
57708 => conv_std_logic_vector(94, 8),
57709 => conv_std_logic_vector(95, 8),
57710 => conv_std_logic_vector(96, 8),
57711 => conv_std_logic_vector(97, 8),
57712 => conv_std_logic_vector(98, 8),
57713 => conv_std_logic_vector(99, 8),
57714 => conv_std_logic_vector(100, 8),
57715 => conv_std_logic_vector(101, 8),
57716 => conv_std_logic_vector(101, 8),
57717 => conv_std_logic_vector(102, 8),
57718 => conv_std_logic_vector(103, 8),
57719 => conv_std_logic_vector(104, 8),
57720 => conv_std_logic_vector(105, 8),
57721 => conv_std_logic_vector(106, 8),
57722 => conv_std_logic_vector(107, 8),
57723 => conv_std_logic_vector(108, 8),
57724 => conv_std_logic_vector(108, 8),
57725 => conv_std_logic_vector(109, 8),
57726 => conv_std_logic_vector(110, 8),
57727 => conv_std_logic_vector(111, 8),
57728 => conv_std_logic_vector(112, 8),
57729 => conv_std_logic_vector(113, 8),
57730 => conv_std_logic_vector(114, 8),
57731 => conv_std_logic_vector(115, 8),
57732 => conv_std_logic_vector(116, 8),
57733 => conv_std_logic_vector(116, 8),
57734 => conv_std_logic_vector(117, 8),
57735 => conv_std_logic_vector(118, 8),
57736 => conv_std_logic_vector(119, 8),
57737 => conv_std_logic_vector(120, 8),
57738 => conv_std_logic_vector(121, 8),
57739 => conv_std_logic_vector(122, 8),
57740 => conv_std_logic_vector(123, 8),
57741 => conv_std_logic_vector(123, 8),
57742 => conv_std_logic_vector(124, 8),
57743 => conv_std_logic_vector(125, 8),
57744 => conv_std_logic_vector(126, 8),
57745 => conv_std_logic_vector(127, 8),
57746 => conv_std_logic_vector(128, 8),
57747 => conv_std_logic_vector(129, 8),
57748 => conv_std_logic_vector(130, 8),
57749 => conv_std_logic_vector(130, 8),
57750 => conv_std_logic_vector(131, 8),
57751 => conv_std_logic_vector(132, 8),
57752 => conv_std_logic_vector(133, 8),
57753 => conv_std_logic_vector(134, 8),
57754 => conv_std_logic_vector(135, 8),
57755 => conv_std_logic_vector(136, 8),
57756 => conv_std_logic_vector(137, 8),
57757 => conv_std_logic_vector(137, 8),
57758 => conv_std_logic_vector(138, 8),
57759 => conv_std_logic_vector(139, 8),
57760 => conv_std_logic_vector(140, 8),
57761 => conv_std_logic_vector(141, 8),
57762 => conv_std_logic_vector(142, 8),
57763 => conv_std_logic_vector(143, 8),
57764 => conv_std_logic_vector(144, 8),
57765 => conv_std_logic_vector(145, 8),
57766 => conv_std_logic_vector(145, 8),
57767 => conv_std_logic_vector(146, 8),
57768 => conv_std_logic_vector(147, 8),
57769 => conv_std_logic_vector(148, 8),
57770 => conv_std_logic_vector(149, 8),
57771 => conv_std_logic_vector(150, 8),
57772 => conv_std_logic_vector(151, 8),
57773 => conv_std_logic_vector(152, 8),
57774 => conv_std_logic_vector(152, 8),
57775 => conv_std_logic_vector(153, 8),
57776 => conv_std_logic_vector(154, 8),
57777 => conv_std_logic_vector(155, 8),
57778 => conv_std_logic_vector(156, 8),
57779 => conv_std_logic_vector(157, 8),
57780 => conv_std_logic_vector(158, 8),
57781 => conv_std_logic_vector(159, 8),
57782 => conv_std_logic_vector(159, 8),
57783 => conv_std_logic_vector(160, 8),
57784 => conv_std_logic_vector(161, 8),
57785 => conv_std_logic_vector(162, 8),
57786 => conv_std_logic_vector(163, 8),
57787 => conv_std_logic_vector(164, 8),
57788 => conv_std_logic_vector(165, 8),
57789 => conv_std_logic_vector(166, 8),
57790 => conv_std_logic_vector(166, 8),
57791 => conv_std_logic_vector(167, 8),
57792 => conv_std_logic_vector(168, 8),
57793 => conv_std_logic_vector(169, 8),
57794 => conv_std_logic_vector(170, 8),
57795 => conv_std_logic_vector(171, 8),
57796 => conv_std_logic_vector(172, 8),
57797 => conv_std_logic_vector(173, 8),
57798 => conv_std_logic_vector(174, 8),
57799 => conv_std_logic_vector(174, 8),
57800 => conv_std_logic_vector(175, 8),
57801 => conv_std_logic_vector(176, 8),
57802 => conv_std_logic_vector(177, 8),
57803 => conv_std_logic_vector(178, 8),
57804 => conv_std_logic_vector(179, 8),
57805 => conv_std_logic_vector(180, 8),
57806 => conv_std_logic_vector(181, 8),
57807 => conv_std_logic_vector(181, 8),
57808 => conv_std_logic_vector(182, 8),
57809 => conv_std_logic_vector(183, 8),
57810 => conv_std_logic_vector(184, 8),
57811 => conv_std_logic_vector(185, 8),
57812 => conv_std_logic_vector(186, 8),
57813 => conv_std_logic_vector(187, 8),
57814 => conv_std_logic_vector(188, 8),
57815 => conv_std_logic_vector(188, 8),
57816 => conv_std_logic_vector(189, 8),
57817 => conv_std_logic_vector(190, 8),
57818 => conv_std_logic_vector(191, 8),
57819 => conv_std_logic_vector(192, 8),
57820 => conv_std_logic_vector(193, 8),
57821 => conv_std_logic_vector(194, 8),
57822 => conv_std_logic_vector(195, 8),
57823 => conv_std_logic_vector(195, 8),
57824 => conv_std_logic_vector(196, 8),
57825 => conv_std_logic_vector(197, 8),
57826 => conv_std_logic_vector(198, 8),
57827 => conv_std_logic_vector(199, 8),
57828 => conv_std_logic_vector(200, 8),
57829 => conv_std_logic_vector(201, 8),
57830 => conv_std_logic_vector(202, 8),
57831 => conv_std_logic_vector(203, 8),
57832 => conv_std_logic_vector(203, 8),
57833 => conv_std_logic_vector(204, 8),
57834 => conv_std_logic_vector(205, 8),
57835 => conv_std_logic_vector(206, 8),
57836 => conv_std_logic_vector(207, 8),
57837 => conv_std_logic_vector(208, 8),
57838 => conv_std_logic_vector(209, 8),
57839 => conv_std_logic_vector(210, 8),
57840 => conv_std_logic_vector(210, 8),
57841 => conv_std_logic_vector(211, 8),
57842 => conv_std_logic_vector(212, 8),
57843 => conv_std_logic_vector(213, 8),
57844 => conv_std_logic_vector(214, 8),
57845 => conv_std_logic_vector(215, 8),
57846 => conv_std_logic_vector(216, 8),
57847 => conv_std_logic_vector(217, 8),
57848 => conv_std_logic_vector(217, 8),
57849 => conv_std_logic_vector(218, 8),
57850 => conv_std_logic_vector(219, 8),
57851 => conv_std_logic_vector(220, 8),
57852 => conv_std_logic_vector(221, 8),
57853 => conv_std_logic_vector(222, 8),
57854 => conv_std_logic_vector(223, 8),
57855 => conv_std_logic_vector(224, 8),
57856 => conv_std_logic_vector(0, 8),
57857 => conv_std_logic_vector(0, 8),
57858 => conv_std_logic_vector(1, 8),
57859 => conv_std_logic_vector(2, 8),
57860 => conv_std_logic_vector(3, 8),
57861 => conv_std_logic_vector(4, 8),
57862 => conv_std_logic_vector(5, 8),
57863 => conv_std_logic_vector(6, 8),
57864 => conv_std_logic_vector(7, 8),
57865 => conv_std_logic_vector(7, 8),
57866 => conv_std_logic_vector(8, 8),
57867 => conv_std_logic_vector(9, 8),
57868 => conv_std_logic_vector(10, 8),
57869 => conv_std_logic_vector(11, 8),
57870 => conv_std_logic_vector(12, 8),
57871 => conv_std_logic_vector(13, 8),
57872 => conv_std_logic_vector(14, 8),
57873 => conv_std_logic_vector(15, 8),
57874 => conv_std_logic_vector(15, 8),
57875 => conv_std_logic_vector(16, 8),
57876 => conv_std_logic_vector(17, 8),
57877 => conv_std_logic_vector(18, 8),
57878 => conv_std_logic_vector(19, 8),
57879 => conv_std_logic_vector(20, 8),
57880 => conv_std_logic_vector(21, 8),
57881 => conv_std_logic_vector(22, 8),
57882 => conv_std_logic_vector(22, 8),
57883 => conv_std_logic_vector(23, 8),
57884 => conv_std_logic_vector(24, 8),
57885 => conv_std_logic_vector(25, 8),
57886 => conv_std_logic_vector(26, 8),
57887 => conv_std_logic_vector(27, 8),
57888 => conv_std_logic_vector(28, 8),
57889 => conv_std_logic_vector(29, 8),
57890 => conv_std_logic_vector(30, 8),
57891 => conv_std_logic_vector(30, 8),
57892 => conv_std_logic_vector(31, 8),
57893 => conv_std_logic_vector(32, 8),
57894 => conv_std_logic_vector(33, 8),
57895 => conv_std_logic_vector(34, 8),
57896 => conv_std_logic_vector(35, 8),
57897 => conv_std_logic_vector(36, 8),
57898 => conv_std_logic_vector(37, 8),
57899 => conv_std_logic_vector(37, 8),
57900 => conv_std_logic_vector(38, 8),
57901 => conv_std_logic_vector(39, 8),
57902 => conv_std_logic_vector(40, 8),
57903 => conv_std_logic_vector(41, 8),
57904 => conv_std_logic_vector(42, 8),
57905 => conv_std_logic_vector(43, 8),
57906 => conv_std_logic_vector(44, 8),
57907 => conv_std_logic_vector(45, 8),
57908 => conv_std_logic_vector(45, 8),
57909 => conv_std_logic_vector(46, 8),
57910 => conv_std_logic_vector(47, 8),
57911 => conv_std_logic_vector(48, 8),
57912 => conv_std_logic_vector(49, 8),
57913 => conv_std_logic_vector(50, 8),
57914 => conv_std_logic_vector(51, 8),
57915 => conv_std_logic_vector(52, 8),
57916 => conv_std_logic_vector(52, 8),
57917 => conv_std_logic_vector(53, 8),
57918 => conv_std_logic_vector(54, 8),
57919 => conv_std_logic_vector(55, 8),
57920 => conv_std_logic_vector(56, 8),
57921 => conv_std_logic_vector(57, 8),
57922 => conv_std_logic_vector(58, 8),
57923 => conv_std_logic_vector(59, 8),
57924 => conv_std_logic_vector(60, 8),
57925 => conv_std_logic_vector(60, 8),
57926 => conv_std_logic_vector(61, 8),
57927 => conv_std_logic_vector(62, 8),
57928 => conv_std_logic_vector(63, 8),
57929 => conv_std_logic_vector(64, 8),
57930 => conv_std_logic_vector(65, 8),
57931 => conv_std_logic_vector(66, 8),
57932 => conv_std_logic_vector(67, 8),
57933 => conv_std_logic_vector(67, 8),
57934 => conv_std_logic_vector(68, 8),
57935 => conv_std_logic_vector(69, 8),
57936 => conv_std_logic_vector(70, 8),
57937 => conv_std_logic_vector(71, 8),
57938 => conv_std_logic_vector(72, 8),
57939 => conv_std_logic_vector(73, 8),
57940 => conv_std_logic_vector(74, 8),
57941 => conv_std_logic_vector(75, 8),
57942 => conv_std_logic_vector(75, 8),
57943 => conv_std_logic_vector(76, 8),
57944 => conv_std_logic_vector(77, 8),
57945 => conv_std_logic_vector(78, 8),
57946 => conv_std_logic_vector(79, 8),
57947 => conv_std_logic_vector(80, 8),
57948 => conv_std_logic_vector(81, 8),
57949 => conv_std_logic_vector(82, 8),
57950 => conv_std_logic_vector(82, 8),
57951 => conv_std_logic_vector(83, 8),
57952 => conv_std_logic_vector(84, 8),
57953 => conv_std_logic_vector(85, 8),
57954 => conv_std_logic_vector(86, 8),
57955 => conv_std_logic_vector(87, 8),
57956 => conv_std_logic_vector(88, 8),
57957 => conv_std_logic_vector(89, 8),
57958 => conv_std_logic_vector(90, 8),
57959 => conv_std_logic_vector(90, 8),
57960 => conv_std_logic_vector(91, 8),
57961 => conv_std_logic_vector(92, 8),
57962 => conv_std_logic_vector(93, 8),
57963 => conv_std_logic_vector(94, 8),
57964 => conv_std_logic_vector(95, 8),
57965 => conv_std_logic_vector(96, 8),
57966 => conv_std_logic_vector(97, 8),
57967 => conv_std_logic_vector(97, 8),
57968 => conv_std_logic_vector(98, 8),
57969 => conv_std_logic_vector(99, 8),
57970 => conv_std_logic_vector(100, 8),
57971 => conv_std_logic_vector(101, 8),
57972 => conv_std_logic_vector(102, 8),
57973 => conv_std_logic_vector(103, 8),
57974 => conv_std_logic_vector(104, 8),
57975 => conv_std_logic_vector(105, 8),
57976 => conv_std_logic_vector(105, 8),
57977 => conv_std_logic_vector(106, 8),
57978 => conv_std_logic_vector(107, 8),
57979 => conv_std_logic_vector(108, 8),
57980 => conv_std_logic_vector(109, 8),
57981 => conv_std_logic_vector(110, 8),
57982 => conv_std_logic_vector(111, 8),
57983 => conv_std_logic_vector(112, 8),
57984 => conv_std_logic_vector(113, 8),
57985 => conv_std_logic_vector(113, 8),
57986 => conv_std_logic_vector(114, 8),
57987 => conv_std_logic_vector(115, 8),
57988 => conv_std_logic_vector(116, 8),
57989 => conv_std_logic_vector(117, 8),
57990 => conv_std_logic_vector(118, 8),
57991 => conv_std_logic_vector(119, 8),
57992 => conv_std_logic_vector(120, 8),
57993 => conv_std_logic_vector(120, 8),
57994 => conv_std_logic_vector(121, 8),
57995 => conv_std_logic_vector(122, 8),
57996 => conv_std_logic_vector(123, 8),
57997 => conv_std_logic_vector(124, 8),
57998 => conv_std_logic_vector(125, 8),
57999 => conv_std_logic_vector(126, 8),
58000 => conv_std_logic_vector(127, 8),
58001 => conv_std_logic_vector(128, 8),
58002 => conv_std_logic_vector(128, 8),
58003 => conv_std_logic_vector(129, 8),
58004 => conv_std_logic_vector(130, 8),
58005 => conv_std_logic_vector(131, 8),
58006 => conv_std_logic_vector(132, 8),
58007 => conv_std_logic_vector(133, 8),
58008 => conv_std_logic_vector(134, 8),
58009 => conv_std_logic_vector(135, 8),
58010 => conv_std_logic_vector(135, 8),
58011 => conv_std_logic_vector(136, 8),
58012 => conv_std_logic_vector(137, 8),
58013 => conv_std_logic_vector(138, 8),
58014 => conv_std_logic_vector(139, 8),
58015 => conv_std_logic_vector(140, 8),
58016 => conv_std_logic_vector(141, 8),
58017 => conv_std_logic_vector(142, 8),
58018 => conv_std_logic_vector(143, 8),
58019 => conv_std_logic_vector(143, 8),
58020 => conv_std_logic_vector(144, 8),
58021 => conv_std_logic_vector(145, 8),
58022 => conv_std_logic_vector(146, 8),
58023 => conv_std_logic_vector(147, 8),
58024 => conv_std_logic_vector(148, 8),
58025 => conv_std_logic_vector(149, 8),
58026 => conv_std_logic_vector(150, 8),
58027 => conv_std_logic_vector(150, 8),
58028 => conv_std_logic_vector(151, 8),
58029 => conv_std_logic_vector(152, 8),
58030 => conv_std_logic_vector(153, 8),
58031 => conv_std_logic_vector(154, 8),
58032 => conv_std_logic_vector(155, 8),
58033 => conv_std_logic_vector(156, 8),
58034 => conv_std_logic_vector(157, 8),
58035 => conv_std_logic_vector(158, 8),
58036 => conv_std_logic_vector(158, 8),
58037 => conv_std_logic_vector(159, 8),
58038 => conv_std_logic_vector(160, 8),
58039 => conv_std_logic_vector(161, 8),
58040 => conv_std_logic_vector(162, 8),
58041 => conv_std_logic_vector(163, 8),
58042 => conv_std_logic_vector(164, 8),
58043 => conv_std_logic_vector(165, 8),
58044 => conv_std_logic_vector(165, 8),
58045 => conv_std_logic_vector(166, 8),
58046 => conv_std_logic_vector(167, 8),
58047 => conv_std_logic_vector(168, 8),
58048 => conv_std_logic_vector(169, 8),
58049 => conv_std_logic_vector(170, 8),
58050 => conv_std_logic_vector(171, 8),
58051 => conv_std_logic_vector(172, 8),
58052 => conv_std_logic_vector(173, 8),
58053 => conv_std_logic_vector(173, 8),
58054 => conv_std_logic_vector(174, 8),
58055 => conv_std_logic_vector(175, 8),
58056 => conv_std_logic_vector(176, 8),
58057 => conv_std_logic_vector(177, 8),
58058 => conv_std_logic_vector(178, 8),
58059 => conv_std_logic_vector(179, 8),
58060 => conv_std_logic_vector(180, 8),
58061 => conv_std_logic_vector(180, 8),
58062 => conv_std_logic_vector(181, 8),
58063 => conv_std_logic_vector(182, 8),
58064 => conv_std_logic_vector(183, 8),
58065 => conv_std_logic_vector(184, 8),
58066 => conv_std_logic_vector(185, 8),
58067 => conv_std_logic_vector(186, 8),
58068 => conv_std_logic_vector(187, 8),
58069 => conv_std_logic_vector(188, 8),
58070 => conv_std_logic_vector(188, 8),
58071 => conv_std_logic_vector(189, 8),
58072 => conv_std_logic_vector(190, 8),
58073 => conv_std_logic_vector(191, 8),
58074 => conv_std_logic_vector(192, 8),
58075 => conv_std_logic_vector(193, 8),
58076 => conv_std_logic_vector(194, 8),
58077 => conv_std_logic_vector(195, 8),
58078 => conv_std_logic_vector(195, 8),
58079 => conv_std_logic_vector(196, 8),
58080 => conv_std_logic_vector(197, 8),
58081 => conv_std_logic_vector(198, 8),
58082 => conv_std_logic_vector(199, 8),
58083 => conv_std_logic_vector(200, 8),
58084 => conv_std_logic_vector(201, 8),
58085 => conv_std_logic_vector(202, 8),
58086 => conv_std_logic_vector(203, 8),
58087 => conv_std_logic_vector(203, 8),
58088 => conv_std_logic_vector(204, 8),
58089 => conv_std_logic_vector(205, 8),
58090 => conv_std_logic_vector(206, 8),
58091 => conv_std_logic_vector(207, 8),
58092 => conv_std_logic_vector(208, 8),
58093 => conv_std_logic_vector(209, 8),
58094 => conv_std_logic_vector(210, 8),
58095 => conv_std_logic_vector(210, 8),
58096 => conv_std_logic_vector(211, 8),
58097 => conv_std_logic_vector(212, 8),
58098 => conv_std_logic_vector(213, 8),
58099 => conv_std_logic_vector(214, 8),
58100 => conv_std_logic_vector(215, 8),
58101 => conv_std_logic_vector(216, 8),
58102 => conv_std_logic_vector(217, 8),
58103 => conv_std_logic_vector(218, 8),
58104 => conv_std_logic_vector(218, 8),
58105 => conv_std_logic_vector(219, 8),
58106 => conv_std_logic_vector(220, 8),
58107 => conv_std_logic_vector(221, 8),
58108 => conv_std_logic_vector(222, 8),
58109 => conv_std_logic_vector(223, 8),
58110 => conv_std_logic_vector(224, 8),
58111 => conv_std_logic_vector(225, 8),
58112 => conv_std_logic_vector(0, 8),
58113 => conv_std_logic_vector(0, 8),
58114 => conv_std_logic_vector(1, 8),
58115 => conv_std_logic_vector(2, 8),
58116 => conv_std_logic_vector(3, 8),
58117 => conv_std_logic_vector(4, 8),
58118 => conv_std_logic_vector(5, 8),
58119 => conv_std_logic_vector(6, 8),
58120 => conv_std_logic_vector(7, 8),
58121 => conv_std_logic_vector(7, 8),
58122 => conv_std_logic_vector(8, 8),
58123 => conv_std_logic_vector(9, 8),
58124 => conv_std_logic_vector(10, 8),
58125 => conv_std_logic_vector(11, 8),
58126 => conv_std_logic_vector(12, 8),
58127 => conv_std_logic_vector(13, 8),
58128 => conv_std_logic_vector(14, 8),
58129 => conv_std_logic_vector(15, 8),
58130 => conv_std_logic_vector(15, 8),
58131 => conv_std_logic_vector(16, 8),
58132 => conv_std_logic_vector(17, 8),
58133 => conv_std_logic_vector(18, 8),
58134 => conv_std_logic_vector(19, 8),
58135 => conv_std_logic_vector(20, 8),
58136 => conv_std_logic_vector(21, 8),
58137 => conv_std_logic_vector(22, 8),
58138 => conv_std_logic_vector(23, 8),
58139 => conv_std_logic_vector(23, 8),
58140 => conv_std_logic_vector(24, 8),
58141 => conv_std_logic_vector(25, 8),
58142 => conv_std_logic_vector(26, 8),
58143 => conv_std_logic_vector(27, 8),
58144 => conv_std_logic_vector(28, 8),
58145 => conv_std_logic_vector(29, 8),
58146 => conv_std_logic_vector(30, 8),
58147 => conv_std_logic_vector(31, 8),
58148 => conv_std_logic_vector(31, 8),
58149 => conv_std_logic_vector(32, 8),
58150 => conv_std_logic_vector(33, 8),
58151 => conv_std_logic_vector(34, 8),
58152 => conv_std_logic_vector(35, 8),
58153 => conv_std_logic_vector(36, 8),
58154 => conv_std_logic_vector(37, 8),
58155 => conv_std_logic_vector(38, 8),
58156 => conv_std_logic_vector(39, 8),
58157 => conv_std_logic_vector(39, 8),
58158 => conv_std_logic_vector(40, 8),
58159 => conv_std_logic_vector(41, 8),
58160 => conv_std_logic_vector(42, 8),
58161 => conv_std_logic_vector(43, 8),
58162 => conv_std_logic_vector(44, 8),
58163 => conv_std_logic_vector(45, 8),
58164 => conv_std_logic_vector(46, 8),
58165 => conv_std_logic_vector(46, 8),
58166 => conv_std_logic_vector(47, 8),
58167 => conv_std_logic_vector(48, 8),
58168 => conv_std_logic_vector(49, 8),
58169 => conv_std_logic_vector(50, 8),
58170 => conv_std_logic_vector(51, 8),
58171 => conv_std_logic_vector(52, 8),
58172 => conv_std_logic_vector(53, 8),
58173 => conv_std_logic_vector(54, 8),
58174 => conv_std_logic_vector(54, 8),
58175 => conv_std_logic_vector(55, 8),
58176 => conv_std_logic_vector(56, 8),
58177 => conv_std_logic_vector(57, 8),
58178 => conv_std_logic_vector(58, 8),
58179 => conv_std_logic_vector(59, 8),
58180 => conv_std_logic_vector(60, 8),
58181 => conv_std_logic_vector(61, 8),
58182 => conv_std_logic_vector(62, 8),
58183 => conv_std_logic_vector(62, 8),
58184 => conv_std_logic_vector(63, 8),
58185 => conv_std_logic_vector(64, 8),
58186 => conv_std_logic_vector(65, 8),
58187 => conv_std_logic_vector(66, 8),
58188 => conv_std_logic_vector(67, 8),
58189 => conv_std_logic_vector(68, 8),
58190 => conv_std_logic_vector(69, 8),
58191 => conv_std_logic_vector(70, 8),
58192 => conv_std_logic_vector(70, 8),
58193 => conv_std_logic_vector(71, 8),
58194 => conv_std_logic_vector(72, 8),
58195 => conv_std_logic_vector(73, 8),
58196 => conv_std_logic_vector(74, 8),
58197 => conv_std_logic_vector(75, 8),
58198 => conv_std_logic_vector(76, 8),
58199 => conv_std_logic_vector(77, 8),
58200 => conv_std_logic_vector(78, 8),
58201 => conv_std_logic_vector(78, 8),
58202 => conv_std_logic_vector(79, 8),
58203 => conv_std_logic_vector(80, 8),
58204 => conv_std_logic_vector(81, 8),
58205 => conv_std_logic_vector(82, 8),
58206 => conv_std_logic_vector(83, 8),
58207 => conv_std_logic_vector(84, 8),
58208 => conv_std_logic_vector(85, 8),
58209 => conv_std_logic_vector(86, 8),
58210 => conv_std_logic_vector(86, 8),
58211 => conv_std_logic_vector(87, 8),
58212 => conv_std_logic_vector(88, 8),
58213 => conv_std_logic_vector(89, 8),
58214 => conv_std_logic_vector(90, 8),
58215 => conv_std_logic_vector(91, 8),
58216 => conv_std_logic_vector(92, 8),
58217 => conv_std_logic_vector(93, 8),
58218 => conv_std_logic_vector(93, 8),
58219 => conv_std_logic_vector(94, 8),
58220 => conv_std_logic_vector(95, 8),
58221 => conv_std_logic_vector(96, 8),
58222 => conv_std_logic_vector(97, 8),
58223 => conv_std_logic_vector(98, 8),
58224 => conv_std_logic_vector(99, 8),
58225 => conv_std_logic_vector(100, 8),
58226 => conv_std_logic_vector(101, 8),
58227 => conv_std_logic_vector(101, 8),
58228 => conv_std_logic_vector(102, 8),
58229 => conv_std_logic_vector(103, 8),
58230 => conv_std_logic_vector(104, 8),
58231 => conv_std_logic_vector(105, 8),
58232 => conv_std_logic_vector(106, 8),
58233 => conv_std_logic_vector(107, 8),
58234 => conv_std_logic_vector(108, 8),
58235 => conv_std_logic_vector(109, 8),
58236 => conv_std_logic_vector(109, 8),
58237 => conv_std_logic_vector(110, 8),
58238 => conv_std_logic_vector(111, 8),
58239 => conv_std_logic_vector(112, 8),
58240 => conv_std_logic_vector(113, 8),
58241 => conv_std_logic_vector(114, 8),
58242 => conv_std_logic_vector(115, 8),
58243 => conv_std_logic_vector(116, 8),
58244 => conv_std_logic_vector(117, 8),
58245 => conv_std_logic_vector(117, 8),
58246 => conv_std_logic_vector(118, 8),
58247 => conv_std_logic_vector(119, 8),
58248 => conv_std_logic_vector(120, 8),
58249 => conv_std_logic_vector(121, 8),
58250 => conv_std_logic_vector(122, 8),
58251 => conv_std_logic_vector(123, 8),
58252 => conv_std_logic_vector(124, 8),
58253 => conv_std_logic_vector(125, 8),
58254 => conv_std_logic_vector(125, 8),
58255 => conv_std_logic_vector(126, 8),
58256 => conv_std_logic_vector(127, 8),
58257 => conv_std_logic_vector(128, 8),
58258 => conv_std_logic_vector(129, 8),
58259 => conv_std_logic_vector(130, 8),
58260 => conv_std_logic_vector(131, 8),
58261 => conv_std_logic_vector(132, 8),
58262 => conv_std_logic_vector(133, 8),
58263 => conv_std_logic_vector(133, 8),
58264 => conv_std_logic_vector(134, 8),
58265 => conv_std_logic_vector(135, 8),
58266 => conv_std_logic_vector(136, 8),
58267 => conv_std_logic_vector(137, 8),
58268 => conv_std_logic_vector(138, 8),
58269 => conv_std_logic_vector(139, 8),
58270 => conv_std_logic_vector(140, 8),
58271 => conv_std_logic_vector(140, 8),
58272 => conv_std_logic_vector(141, 8),
58273 => conv_std_logic_vector(142, 8),
58274 => conv_std_logic_vector(143, 8),
58275 => conv_std_logic_vector(144, 8),
58276 => conv_std_logic_vector(145, 8),
58277 => conv_std_logic_vector(146, 8),
58278 => conv_std_logic_vector(147, 8),
58279 => conv_std_logic_vector(148, 8),
58280 => conv_std_logic_vector(148, 8),
58281 => conv_std_logic_vector(149, 8),
58282 => conv_std_logic_vector(150, 8),
58283 => conv_std_logic_vector(151, 8),
58284 => conv_std_logic_vector(152, 8),
58285 => conv_std_logic_vector(153, 8),
58286 => conv_std_logic_vector(154, 8),
58287 => conv_std_logic_vector(155, 8),
58288 => conv_std_logic_vector(156, 8),
58289 => conv_std_logic_vector(156, 8),
58290 => conv_std_logic_vector(157, 8),
58291 => conv_std_logic_vector(158, 8),
58292 => conv_std_logic_vector(159, 8),
58293 => conv_std_logic_vector(160, 8),
58294 => conv_std_logic_vector(161, 8),
58295 => conv_std_logic_vector(162, 8),
58296 => conv_std_logic_vector(163, 8),
58297 => conv_std_logic_vector(164, 8),
58298 => conv_std_logic_vector(164, 8),
58299 => conv_std_logic_vector(165, 8),
58300 => conv_std_logic_vector(166, 8),
58301 => conv_std_logic_vector(167, 8),
58302 => conv_std_logic_vector(168, 8),
58303 => conv_std_logic_vector(169, 8),
58304 => conv_std_logic_vector(170, 8),
58305 => conv_std_logic_vector(171, 8),
58306 => conv_std_logic_vector(172, 8),
58307 => conv_std_logic_vector(172, 8),
58308 => conv_std_logic_vector(173, 8),
58309 => conv_std_logic_vector(174, 8),
58310 => conv_std_logic_vector(175, 8),
58311 => conv_std_logic_vector(176, 8),
58312 => conv_std_logic_vector(177, 8),
58313 => conv_std_logic_vector(178, 8),
58314 => conv_std_logic_vector(179, 8),
58315 => conv_std_logic_vector(180, 8),
58316 => conv_std_logic_vector(180, 8),
58317 => conv_std_logic_vector(181, 8),
58318 => conv_std_logic_vector(182, 8),
58319 => conv_std_logic_vector(183, 8),
58320 => conv_std_logic_vector(184, 8),
58321 => conv_std_logic_vector(185, 8),
58322 => conv_std_logic_vector(186, 8),
58323 => conv_std_logic_vector(187, 8),
58324 => conv_std_logic_vector(187, 8),
58325 => conv_std_logic_vector(188, 8),
58326 => conv_std_logic_vector(189, 8),
58327 => conv_std_logic_vector(190, 8),
58328 => conv_std_logic_vector(191, 8),
58329 => conv_std_logic_vector(192, 8),
58330 => conv_std_logic_vector(193, 8),
58331 => conv_std_logic_vector(194, 8),
58332 => conv_std_logic_vector(195, 8),
58333 => conv_std_logic_vector(195, 8),
58334 => conv_std_logic_vector(196, 8),
58335 => conv_std_logic_vector(197, 8),
58336 => conv_std_logic_vector(198, 8),
58337 => conv_std_logic_vector(199, 8),
58338 => conv_std_logic_vector(200, 8),
58339 => conv_std_logic_vector(201, 8),
58340 => conv_std_logic_vector(202, 8),
58341 => conv_std_logic_vector(203, 8),
58342 => conv_std_logic_vector(203, 8),
58343 => conv_std_logic_vector(204, 8),
58344 => conv_std_logic_vector(205, 8),
58345 => conv_std_logic_vector(206, 8),
58346 => conv_std_logic_vector(207, 8),
58347 => conv_std_logic_vector(208, 8),
58348 => conv_std_logic_vector(209, 8),
58349 => conv_std_logic_vector(210, 8),
58350 => conv_std_logic_vector(211, 8),
58351 => conv_std_logic_vector(211, 8),
58352 => conv_std_logic_vector(212, 8),
58353 => conv_std_logic_vector(213, 8),
58354 => conv_std_logic_vector(214, 8),
58355 => conv_std_logic_vector(215, 8),
58356 => conv_std_logic_vector(216, 8),
58357 => conv_std_logic_vector(217, 8),
58358 => conv_std_logic_vector(218, 8),
58359 => conv_std_logic_vector(219, 8),
58360 => conv_std_logic_vector(219, 8),
58361 => conv_std_logic_vector(220, 8),
58362 => conv_std_logic_vector(221, 8),
58363 => conv_std_logic_vector(222, 8),
58364 => conv_std_logic_vector(223, 8),
58365 => conv_std_logic_vector(224, 8),
58366 => conv_std_logic_vector(225, 8),
58367 => conv_std_logic_vector(226, 8),
58368 => conv_std_logic_vector(0, 8),
58369 => conv_std_logic_vector(0, 8),
58370 => conv_std_logic_vector(1, 8),
58371 => conv_std_logic_vector(2, 8),
58372 => conv_std_logic_vector(3, 8),
58373 => conv_std_logic_vector(4, 8),
58374 => conv_std_logic_vector(5, 8),
58375 => conv_std_logic_vector(6, 8),
58376 => conv_std_logic_vector(7, 8),
58377 => conv_std_logic_vector(8, 8),
58378 => conv_std_logic_vector(8, 8),
58379 => conv_std_logic_vector(9, 8),
58380 => conv_std_logic_vector(10, 8),
58381 => conv_std_logic_vector(11, 8),
58382 => conv_std_logic_vector(12, 8),
58383 => conv_std_logic_vector(13, 8),
58384 => conv_std_logic_vector(14, 8),
58385 => conv_std_logic_vector(15, 8),
58386 => conv_std_logic_vector(16, 8),
58387 => conv_std_logic_vector(16, 8),
58388 => conv_std_logic_vector(17, 8),
58389 => conv_std_logic_vector(18, 8),
58390 => conv_std_logic_vector(19, 8),
58391 => conv_std_logic_vector(20, 8),
58392 => conv_std_logic_vector(21, 8),
58393 => conv_std_logic_vector(22, 8),
58394 => conv_std_logic_vector(23, 8),
58395 => conv_std_logic_vector(24, 8),
58396 => conv_std_logic_vector(24, 8),
58397 => conv_std_logic_vector(25, 8),
58398 => conv_std_logic_vector(26, 8),
58399 => conv_std_logic_vector(27, 8),
58400 => conv_std_logic_vector(28, 8),
58401 => conv_std_logic_vector(29, 8),
58402 => conv_std_logic_vector(30, 8),
58403 => conv_std_logic_vector(31, 8),
58404 => conv_std_logic_vector(32, 8),
58405 => conv_std_logic_vector(32, 8),
58406 => conv_std_logic_vector(33, 8),
58407 => conv_std_logic_vector(34, 8),
58408 => conv_std_logic_vector(35, 8),
58409 => conv_std_logic_vector(36, 8),
58410 => conv_std_logic_vector(37, 8),
58411 => conv_std_logic_vector(38, 8),
58412 => conv_std_logic_vector(39, 8),
58413 => conv_std_logic_vector(40, 8),
58414 => conv_std_logic_vector(40, 8),
58415 => conv_std_logic_vector(41, 8),
58416 => conv_std_logic_vector(42, 8),
58417 => conv_std_logic_vector(43, 8),
58418 => conv_std_logic_vector(44, 8),
58419 => conv_std_logic_vector(45, 8),
58420 => conv_std_logic_vector(46, 8),
58421 => conv_std_logic_vector(47, 8),
58422 => conv_std_logic_vector(48, 8),
58423 => conv_std_logic_vector(48, 8),
58424 => conv_std_logic_vector(49, 8),
58425 => conv_std_logic_vector(50, 8),
58426 => conv_std_logic_vector(51, 8),
58427 => conv_std_logic_vector(52, 8),
58428 => conv_std_logic_vector(53, 8),
58429 => conv_std_logic_vector(54, 8),
58430 => conv_std_logic_vector(55, 8),
58431 => conv_std_logic_vector(56, 8),
58432 => conv_std_logic_vector(57, 8),
58433 => conv_std_logic_vector(57, 8),
58434 => conv_std_logic_vector(58, 8),
58435 => conv_std_logic_vector(59, 8),
58436 => conv_std_logic_vector(60, 8),
58437 => conv_std_logic_vector(61, 8),
58438 => conv_std_logic_vector(62, 8),
58439 => conv_std_logic_vector(63, 8),
58440 => conv_std_logic_vector(64, 8),
58441 => conv_std_logic_vector(65, 8),
58442 => conv_std_logic_vector(65, 8),
58443 => conv_std_logic_vector(66, 8),
58444 => conv_std_logic_vector(67, 8),
58445 => conv_std_logic_vector(68, 8),
58446 => conv_std_logic_vector(69, 8),
58447 => conv_std_logic_vector(70, 8),
58448 => conv_std_logic_vector(71, 8),
58449 => conv_std_logic_vector(72, 8),
58450 => conv_std_logic_vector(73, 8),
58451 => conv_std_logic_vector(73, 8),
58452 => conv_std_logic_vector(74, 8),
58453 => conv_std_logic_vector(75, 8),
58454 => conv_std_logic_vector(76, 8),
58455 => conv_std_logic_vector(77, 8),
58456 => conv_std_logic_vector(78, 8),
58457 => conv_std_logic_vector(79, 8),
58458 => conv_std_logic_vector(80, 8),
58459 => conv_std_logic_vector(81, 8),
58460 => conv_std_logic_vector(81, 8),
58461 => conv_std_logic_vector(82, 8),
58462 => conv_std_logic_vector(83, 8),
58463 => conv_std_logic_vector(84, 8),
58464 => conv_std_logic_vector(85, 8),
58465 => conv_std_logic_vector(86, 8),
58466 => conv_std_logic_vector(87, 8),
58467 => conv_std_logic_vector(88, 8),
58468 => conv_std_logic_vector(89, 8),
58469 => conv_std_logic_vector(89, 8),
58470 => conv_std_logic_vector(90, 8),
58471 => conv_std_logic_vector(91, 8),
58472 => conv_std_logic_vector(92, 8),
58473 => conv_std_logic_vector(93, 8),
58474 => conv_std_logic_vector(94, 8),
58475 => conv_std_logic_vector(95, 8),
58476 => conv_std_logic_vector(96, 8),
58477 => conv_std_logic_vector(97, 8),
58478 => conv_std_logic_vector(97, 8),
58479 => conv_std_logic_vector(98, 8),
58480 => conv_std_logic_vector(99, 8),
58481 => conv_std_logic_vector(100, 8),
58482 => conv_std_logic_vector(101, 8),
58483 => conv_std_logic_vector(102, 8),
58484 => conv_std_logic_vector(103, 8),
58485 => conv_std_logic_vector(104, 8),
58486 => conv_std_logic_vector(105, 8),
58487 => conv_std_logic_vector(105, 8),
58488 => conv_std_logic_vector(106, 8),
58489 => conv_std_logic_vector(107, 8),
58490 => conv_std_logic_vector(108, 8),
58491 => conv_std_logic_vector(109, 8),
58492 => conv_std_logic_vector(110, 8),
58493 => conv_std_logic_vector(111, 8),
58494 => conv_std_logic_vector(112, 8),
58495 => conv_std_logic_vector(113, 8),
58496 => conv_std_logic_vector(114, 8),
58497 => conv_std_logic_vector(114, 8),
58498 => conv_std_logic_vector(115, 8),
58499 => conv_std_logic_vector(116, 8),
58500 => conv_std_logic_vector(117, 8),
58501 => conv_std_logic_vector(118, 8),
58502 => conv_std_logic_vector(119, 8),
58503 => conv_std_logic_vector(120, 8),
58504 => conv_std_logic_vector(121, 8),
58505 => conv_std_logic_vector(122, 8),
58506 => conv_std_logic_vector(122, 8),
58507 => conv_std_logic_vector(123, 8),
58508 => conv_std_logic_vector(124, 8),
58509 => conv_std_logic_vector(125, 8),
58510 => conv_std_logic_vector(126, 8),
58511 => conv_std_logic_vector(127, 8),
58512 => conv_std_logic_vector(128, 8),
58513 => conv_std_logic_vector(129, 8),
58514 => conv_std_logic_vector(130, 8),
58515 => conv_std_logic_vector(130, 8),
58516 => conv_std_logic_vector(131, 8),
58517 => conv_std_logic_vector(132, 8),
58518 => conv_std_logic_vector(133, 8),
58519 => conv_std_logic_vector(134, 8),
58520 => conv_std_logic_vector(135, 8),
58521 => conv_std_logic_vector(136, 8),
58522 => conv_std_logic_vector(137, 8),
58523 => conv_std_logic_vector(138, 8),
58524 => conv_std_logic_vector(138, 8),
58525 => conv_std_logic_vector(139, 8),
58526 => conv_std_logic_vector(140, 8),
58527 => conv_std_logic_vector(141, 8),
58528 => conv_std_logic_vector(142, 8),
58529 => conv_std_logic_vector(143, 8),
58530 => conv_std_logic_vector(144, 8),
58531 => conv_std_logic_vector(145, 8),
58532 => conv_std_logic_vector(146, 8),
58533 => conv_std_logic_vector(146, 8),
58534 => conv_std_logic_vector(147, 8),
58535 => conv_std_logic_vector(148, 8),
58536 => conv_std_logic_vector(149, 8),
58537 => conv_std_logic_vector(150, 8),
58538 => conv_std_logic_vector(151, 8),
58539 => conv_std_logic_vector(152, 8),
58540 => conv_std_logic_vector(153, 8),
58541 => conv_std_logic_vector(154, 8),
58542 => conv_std_logic_vector(154, 8),
58543 => conv_std_logic_vector(155, 8),
58544 => conv_std_logic_vector(156, 8),
58545 => conv_std_logic_vector(157, 8),
58546 => conv_std_logic_vector(158, 8),
58547 => conv_std_logic_vector(159, 8),
58548 => conv_std_logic_vector(160, 8),
58549 => conv_std_logic_vector(161, 8),
58550 => conv_std_logic_vector(162, 8),
58551 => conv_std_logic_vector(162, 8),
58552 => conv_std_logic_vector(163, 8),
58553 => conv_std_logic_vector(164, 8),
58554 => conv_std_logic_vector(165, 8),
58555 => conv_std_logic_vector(166, 8),
58556 => conv_std_logic_vector(167, 8),
58557 => conv_std_logic_vector(168, 8),
58558 => conv_std_logic_vector(169, 8),
58559 => conv_std_logic_vector(170, 8),
58560 => conv_std_logic_vector(171, 8),
58561 => conv_std_logic_vector(171, 8),
58562 => conv_std_logic_vector(172, 8),
58563 => conv_std_logic_vector(173, 8),
58564 => conv_std_logic_vector(174, 8),
58565 => conv_std_logic_vector(175, 8),
58566 => conv_std_logic_vector(176, 8),
58567 => conv_std_logic_vector(177, 8),
58568 => conv_std_logic_vector(178, 8),
58569 => conv_std_logic_vector(179, 8),
58570 => conv_std_logic_vector(179, 8),
58571 => conv_std_logic_vector(180, 8),
58572 => conv_std_logic_vector(181, 8),
58573 => conv_std_logic_vector(182, 8),
58574 => conv_std_logic_vector(183, 8),
58575 => conv_std_logic_vector(184, 8),
58576 => conv_std_logic_vector(185, 8),
58577 => conv_std_logic_vector(186, 8),
58578 => conv_std_logic_vector(187, 8),
58579 => conv_std_logic_vector(187, 8),
58580 => conv_std_logic_vector(188, 8),
58581 => conv_std_logic_vector(189, 8),
58582 => conv_std_logic_vector(190, 8),
58583 => conv_std_logic_vector(191, 8),
58584 => conv_std_logic_vector(192, 8),
58585 => conv_std_logic_vector(193, 8),
58586 => conv_std_logic_vector(194, 8),
58587 => conv_std_logic_vector(195, 8),
58588 => conv_std_logic_vector(195, 8),
58589 => conv_std_logic_vector(196, 8),
58590 => conv_std_logic_vector(197, 8),
58591 => conv_std_logic_vector(198, 8),
58592 => conv_std_logic_vector(199, 8),
58593 => conv_std_logic_vector(200, 8),
58594 => conv_std_logic_vector(201, 8),
58595 => conv_std_logic_vector(202, 8),
58596 => conv_std_logic_vector(203, 8),
58597 => conv_std_logic_vector(203, 8),
58598 => conv_std_logic_vector(204, 8),
58599 => conv_std_logic_vector(205, 8),
58600 => conv_std_logic_vector(206, 8),
58601 => conv_std_logic_vector(207, 8),
58602 => conv_std_logic_vector(208, 8),
58603 => conv_std_logic_vector(209, 8),
58604 => conv_std_logic_vector(210, 8),
58605 => conv_std_logic_vector(211, 8),
58606 => conv_std_logic_vector(211, 8),
58607 => conv_std_logic_vector(212, 8),
58608 => conv_std_logic_vector(213, 8),
58609 => conv_std_logic_vector(214, 8),
58610 => conv_std_logic_vector(215, 8),
58611 => conv_std_logic_vector(216, 8),
58612 => conv_std_logic_vector(217, 8),
58613 => conv_std_logic_vector(218, 8),
58614 => conv_std_logic_vector(219, 8),
58615 => conv_std_logic_vector(219, 8),
58616 => conv_std_logic_vector(220, 8),
58617 => conv_std_logic_vector(221, 8),
58618 => conv_std_logic_vector(222, 8),
58619 => conv_std_logic_vector(223, 8),
58620 => conv_std_logic_vector(224, 8),
58621 => conv_std_logic_vector(225, 8),
58622 => conv_std_logic_vector(226, 8),
58623 => conv_std_logic_vector(227, 8),
58624 => conv_std_logic_vector(0, 8),
58625 => conv_std_logic_vector(0, 8),
58626 => conv_std_logic_vector(1, 8),
58627 => conv_std_logic_vector(2, 8),
58628 => conv_std_logic_vector(3, 8),
58629 => conv_std_logic_vector(4, 8),
58630 => conv_std_logic_vector(5, 8),
58631 => conv_std_logic_vector(6, 8),
58632 => conv_std_logic_vector(7, 8),
58633 => conv_std_logic_vector(8, 8),
58634 => conv_std_logic_vector(8, 8),
58635 => conv_std_logic_vector(9, 8),
58636 => conv_std_logic_vector(10, 8),
58637 => conv_std_logic_vector(11, 8),
58638 => conv_std_logic_vector(12, 8),
58639 => conv_std_logic_vector(13, 8),
58640 => conv_std_logic_vector(14, 8),
58641 => conv_std_logic_vector(15, 8),
58642 => conv_std_logic_vector(16, 8),
58643 => conv_std_logic_vector(16, 8),
58644 => conv_std_logic_vector(17, 8),
58645 => conv_std_logic_vector(18, 8),
58646 => conv_std_logic_vector(19, 8),
58647 => conv_std_logic_vector(20, 8),
58648 => conv_std_logic_vector(21, 8),
58649 => conv_std_logic_vector(22, 8),
58650 => conv_std_logic_vector(23, 8),
58651 => conv_std_logic_vector(24, 8),
58652 => conv_std_logic_vector(25, 8),
58653 => conv_std_logic_vector(25, 8),
58654 => conv_std_logic_vector(26, 8),
58655 => conv_std_logic_vector(27, 8),
58656 => conv_std_logic_vector(28, 8),
58657 => conv_std_logic_vector(29, 8),
58658 => conv_std_logic_vector(30, 8),
58659 => conv_std_logic_vector(31, 8),
58660 => conv_std_logic_vector(32, 8),
58661 => conv_std_logic_vector(33, 8),
58662 => conv_std_logic_vector(33, 8),
58663 => conv_std_logic_vector(34, 8),
58664 => conv_std_logic_vector(35, 8),
58665 => conv_std_logic_vector(36, 8),
58666 => conv_std_logic_vector(37, 8),
58667 => conv_std_logic_vector(38, 8),
58668 => conv_std_logic_vector(39, 8),
58669 => conv_std_logic_vector(40, 8),
58670 => conv_std_logic_vector(41, 8),
58671 => conv_std_logic_vector(42, 8),
58672 => conv_std_logic_vector(42, 8),
58673 => conv_std_logic_vector(43, 8),
58674 => conv_std_logic_vector(44, 8),
58675 => conv_std_logic_vector(45, 8),
58676 => conv_std_logic_vector(46, 8),
58677 => conv_std_logic_vector(47, 8),
58678 => conv_std_logic_vector(48, 8),
58679 => conv_std_logic_vector(49, 8),
58680 => conv_std_logic_vector(50, 8),
58681 => conv_std_logic_vector(50, 8),
58682 => conv_std_logic_vector(51, 8),
58683 => conv_std_logic_vector(52, 8),
58684 => conv_std_logic_vector(53, 8),
58685 => conv_std_logic_vector(54, 8),
58686 => conv_std_logic_vector(55, 8),
58687 => conv_std_logic_vector(56, 8),
58688 => conv_std_logic_vector(57, 8),
58689 => conv_std_logic_vector(58, 8),
58690 => conv_std_logic_vector(59, 8),
58691 => conv_std_logic_vector(59, 8),
58692 => conv_std_logic_vector(60, 8),
58693 => conv_std_logic_vector(61, 8),
58694 => conv_std_logic_vector(62, 8),
58695 => conv_std_logic_vector(63, 8),
58696 => conv_std_logic_vector(64, 8),
58697 => conv_std_logic_vector(65, 8),
58698 => conv_std_logic_vector(66, 8),
58699 => conv_std_logic_vector(67, 8),
58700 => conv_std_logic_vector(67, 8),
58701 => conv_std_logic_vector(68, 8),
58702 => conv_std_logic_vector(69, 8),
58703 => conv_std_logic_vector(70, 8),
58704 => conv_std_logic_vector(71, 8),
58705 => conv_std_logic_vector(72, 8),
58706 => conv_std_logic_vector(73, 8),
58707 => conv_std_logic_vector(74, 8),
58708 => conv_std_logic_vector(75, 8),
58709 => conv_std_logic_vector(76, 8),
58710 => conv_std_logic_vector(76, 8),
58711 => conv_std_logic_vector(77, 8),
58712 => conv_std_logic_vector(78, 8),
58713 => conv_std_logic_vector(79, 8),
58714 => conv_std_logic_vector(80, 8),
58715 => conv_std_logic_vector(81, 8),
58716 => conv_std_logic_vector(82, 8),
58717 => conv_std_logic_vector(83, 8),
58718 => conv_std_logic_vector(84, 8),
58719 => conv_std_logic_vector(84, 8),
58720 => conv_std_logic_vector(85, 8),
58721 => conv_std_logic_vector(86, 8),
58722 => conv_std_logic_vector(87, 8),
58723 => conv_std_logic_vector(88, 8),
58724 => conv_std_logic_vector(89, 8),
58725 => conv_std_logic_vector(90, 8),
58726 => conv_std_logic_vector(91, 8),
58727 => conv_std_logic_vector(92, 8),
58728 => conv_std_logic_vector(93, 8),
58729 => conv_std_logic_vector(93, 8),
58730 => conv_std_logic_vector(94, 8),
58731 => conv_std_logic_vector(95, 8),
58732 => conv_std_logic_vector(96, 8),
58733 => conv_std_logic_vector(97, 8),
58734 => conv_std_logic_vector(98, 8),
58735 => conv_std_logic_vector(99, 8),
58736 => conv_std_logic_vector(100, 8),
58737 => conv_std_logic_vector(101, 8),
58738 => conv_std_logic_vector(101, 8),
58739 => conv_std_logic_vector(102, 8),
58740 => conv_std_logic_vector(103, 8),
58741 => conv_std_logic_vector(104, 8),
58742 => conv_std_logic_vector(105, 8),
58743 => conv_std_logic_vector(106, 8),
58744 => conv_std_logic_vector(107, 8),
58745 => conv_std_logic_vector(108, 8),
58746 => conv_std_logic_vector(109, 8),
58747 => conv_std_logic_vector(110, 8),
58748 => conv_std_logic_vector(110, 8),
58749 => conv_std_logic_vector(111, 8),
58750 => conv_std_logic_vector(112, 8),
58751 => conv_std_logic_vector(113, 8),
58752 => conv_std_logic_vector(114, 8),
58753 => conv_std_logic_vector(115, 8),
58754 => conv_std_logic_vector(116, 8),
58755 => conv_std_logic_vector(117, 8),
58756 => conv_std_logic_vector(118, 8),
58757 => conv_std_logic_vector(118, 8),
58758 => conv_std_logic_vector(119, 8),
58759 => conv_std_logic_vector(120, 8),
58760 => conv_std_logic_vector(121, 8),
58761 => conv_std_logic_vector(122, 8),
58762 => conv_std_logic_vector(123, 8),
58763 => conv_std_logic_vector(124, 8),
58764 => conv_std_logic_vector(125, 8),
58765 => conv_std_logic_vector(126, 8),
58766 => conv_std_logic_vector(127, 8),
58767 => conv_std_logic_vector(127, 8),
58768 => conv_std_logic_vector(128, 8),
58769 => conv_std_logic_vector(129, 8),
58770 => conv_std_logic_vector(130, 8),
58771 => conv_std_logic_vector(131, 8),
58772 => conv_std_logic_vector(132, 8),
58773 => conv_std_logic_vector(133, 8),
58774 => conv_std_logic_vector(134, 8),
58775 => conv_std_logic_vector(135, 8),
58776 => conv_std_logic_vector(135, 8),
58777 => conv_std_logic_vector(136, 8),
58778 => conv_std_logic_vector(137, 8),
58779 => conv_std_logic_vector(138, 8),
58780 => conv_std_logic_vector(139, 8),
58781 => conv_std_logic_vector(140, 8),
58782 => conv_std_logic_vector(141, 8),
58783 => conv_std_logic_vector(142, 8),
58784 => conv_std_logic_vector(143, 8),
58785 => conv_std_logic_vector(144, 8),
58786 => conv_std_logic_vector(144, 8),
58787 => conv_std_logic_vector(145, 8),
58788 => conv_std_logic_vector(146, 8),
58789 => conv_std_logic_vector(147, 8),
58790 => conv_std_logic_vector(148, 8),
58791 => conv_std_logic_vector(149, 8),
58792 => conv_std_logic_vector(150, 8),
58793 => conv_std_logic_vector(151, 8),
58794 => conv_std_logic_vector(152, 8),
58795 => conv_std_logic_vector(152, 8),
58796 => conv_std_logic_vector(153, 8),
58797 => conv_std_logic_vector(154, 8),
58798 => conv_std_logic_vector(155, 8),
58799 => conv_std_logic_vector(156, 8),
58800 => conv_std_logic_vector(157, 8),
58801 => conv_std_logic_vector(158, 8),
58802 => conv_std_logic_vector(159, 8),
58803 => conv_std_logic_vector(160, 8),
58804 => conv_std_logic_vector(161, 8),
58805 => conv_std_logic_vector(161, 8),
58806 => conv_std_logic_vector(162, 8),
58807 => conv_std_logic_vector(163, 8),
58808 => conv_std_logic_vector(164, 8),
58809 => conv_std_logic_vector(165, 8),
58810 => conv_std_logic_vector(166, 8),
58811 => conv_std_logic_vector(167, 8),
58812 => conv_std_logic_vector(168, 8),
58813 => conv_std_logic_vector(169, 8),
58814 => conv_std_logic_vector(169, 8),
58815 => conv_std_logic_vector(170, 8),
58816 => conv_std_logic_vector(171, 8),
58817 => conv_std_logic_vector(172, 8),
58818 => conv_std_logic_vector(173, 8),
58819 => conv_std_logic_vector(174, 8),
58820 => conv_std_logic_vector(175, 8),
58821 => conv_std_logic_vector(176, 8),
58822 => conv_std_logic_vector(177, 8),
58823 => conv_std_logic_vector(178, 8),
58824 => conv_std_logic_vector(178, 8),
58825 => conv_std_logic_vector(179, 8),
58826 => conv_std_logic_vector(180, 8),
58827 => conv_std_logic_vector(181, 8),
58828 => conv_std_logic_vector(182, 8),
58829 => conv_std_logic_vector(183, 8),
58830 => conv_std_logic_vector(184, 8),
58831 => conv_std_logic_vector(185, 8),
58832 => conv_std_logic_vector(186, 8),
58833 => conv_std_logic_vector(186, 8),
58834 => conv_std_logic_vector(187, 8),
58835 => conv_std_logic_vector(188, 8),
58836 => conv_std_logic_vector(189, 8),
58837 => conv_std_logic_vector(190, 8),
58838 => conv_std_logic_vector(191, 8),
58839 => conv_std_logic_vector(192, 8),
58840 => conv_std_logic_vector(193, 8),
58841 => conv_std_logic_vector(194, 8),
58842 => conv_std_logic_vector(195, 8),
58843 => conv_std_logic_vector(195, 8),
58844 => conv_std_logic_vector(196, 8),
58845 => conv_std_logic_vector(197, 8),
58846 => conv_std_logic_vector(198, 8),
58847 => conv_std_logic_vector(199, 8),
58848 => conv_std_logic_vector(200, 8),
58849 => conv_std_logic_vector(201, 8),
58850 => conv_std_logic_vector(202, 8),
58851 => conv_std_logic_vector(203, 8),
58852 => conv_std_logic_vector(203, 8),
58853 => conv_std_logic_vector(204, 8),
58854 => conv_std_logic_vector(205, 8),
58855 => conv_std_logic_vector(206, 8),
58856 => conv_std_logic_vector(207, 8),
58857 => conv_std_logic_vector(208, 8),
58858 => conv_std_logic_vector(209, 8),
58859 => conv_std_logic_vector(210, 8),
58860 => conv_std_logic_vector(211, 8),
58861 => conv_std_logic_vector(212, 8),
58862 => conv_std_logic_vector(212, 8),
58863 => conv_std_logic_vector(213, 8),
58864 => conv_std_logic_vector(214, 8),
58865 => conv_std_logic_vector(215, 8),
58866 => conv_std_logic_vector(216, 8),
58867 => conv_std_logic_vector(217, 8),
58868 => conv_std_logic_vector(218, 8),
58869 => conv_std_logic_vector(219, 8),
58870 => conv_std_logic_vector(220, 8),
58871 => conv_std_logic_vector(220, 8),
58872 => conv_std_logic_vector(221, 8),
58873 => conv_std_logic_vector(222, 8),
58874 => conv_std_logic_vector(223, 8),
58875 => conv_std_logic_vector(224, 8),
58876 => conv_std_logic_vector(225, 8),
58877 => conv_std_logic_vector(226, 8),
58878 => conv_std_logic_vector(227, 8),
58879 => conv_std_logic_vector(228, 8),
58880 => conv_std_logic_vector(0, 8),
58881 => conv_std_logic_vector(0, 8),
58882 => conv_std_logic_vector(1, 8),
58883 => conv_std_logic_vector(2, 8),
58884 => conv_std_logic_vector(3, 8),
58885 => conv_std_logic_vector(4, 8),
58886 => conv_std_logic_vector(5, 8),
58887 => conv_std_logic_vector(6, 8),
58888 => conv_std_logic_vector(7, 8),
58889 => conv_std_logic_vector(8, 8),
58890 => conv_std_logic_vector(8, 8),
58891 => conv_std_logic_vector(9, 8),
58892 => conv_std_logic_vector(10, 8),
58893 => conv_std_logic_vector(11, 8),
58894 => conv_std_logic_vector(12, 8),
58895 => conv_std_logic_vector(13, 8),
58896 => conv_std_logic_vector(14, 8),
58897 => conv_std_logic_vector(15, 8),
58898 => conv_std_logic_vector(16, 8),
58899 => conv_std_logic_vector(17, 8),
58900 => conv_std_logic_vector(17, 8),
58901 => conv_std_logic_vector(18, 8),
58902 => conv_std_logic_vector(19, 8),
58903 => conv_std_logic_vector(20, 8),
58904 => conv_std_logic_vector(21, 8),
58905 => conv_std_logic_vector(22, 8),
58906 => conv_std_logic_vector(23, 8),
58907 => conv_std_logic_vector(24, 8),
58908 => conv_std_logic_vector(25, 8),
58909 => conv_std_logic_vector(26, 8),
58910 => conv_std_logic_vector(26, 8),
58911 => conv_std_logic_vector(27, 8),
58912 => conv_std_logic_vector(28, 8),
58913 => conv_std_logic_vector(29, 8),
58914 => conv_std_logic_vector(30, 8),
58915 => conv_std_logic_vector(31, 8),
58916 => conv_std_logic_vector(32, 8),
58917 => conv_std_logic_vector(33, 8),
58918 => conv_std_logic_vector(34, 8),
58919 => conv_std_logic_vector(35, 8),
58920 => conv_std_logic_vector(35, 8),
58921 => conv_std_logic_vector(36, 8),
58922 => conv_std_logic_vector(37, 8),
58923 => conv_std_logic_vector(38, 8),
58924 => conv_std_logic_vector(39, 8),
58925 => conv_std_logic_vector(40, 8),
58926 => conv_std_logic_vector(41, 8),
58927 => conv_std_logic_vector(42, 8),
58928 => conv_std_logic_vector(43, 8),
58929 => conv_std_logic_vector(44, 8),
58930 => conv_std_logic_vector(44, 8),
58931 => conv_std_logic_vector(45, 8),
58932 => conv_std_logic_vector(46, 8),
58933 => conv_std_logic_vector(47, 8),
58934 => conv_std_logic_vector(48, 8),
58935 => conv_std_logic_vector(49, 8),
58936 => conv_std_logic_vector(50, 8),
58937 => conv_std_logic_vector(51, 8),
58938 => conv_std_logic_vector(52, 8),
58939 => conv_std_logic_vector(53, 8),
58940 => conv_std_logic_vector(53, 8),
58941 => conv_std_logic_vector(54, 8),
58942 => conv_std_logic_vector(55, 8),
58943 => conv_std_logic_vector(56, 8),
58944 => conv_std_logic_vector(57, 8),
58945 => conv_std_logic_vector(58, 8),
58946 => conv_std_logic_vector(59, 8),
58947 => conv_std_logic_vector(60, 8),
58948 => conv_std_logic_vector(61, 8),
58949 => conv_std_logic_vector(61, 8),
58950 => conv_std_logic_vector(62, 8),
58951 => conv_std_logic_vector(63, 8),
58952 => conv_std_logic_vector(64, 8),
58953 => conv_std_logic_vector(65, 8),
58954 => conv_std_logic_vector(66, 8),
58955 => conv_std_logic_vector(67, 8),
58956 => conv_std_logic_vector(68, 8),
58957 => conv_std_logic_vector(69, 8),
58958 => conv_std_logic_vector(70, 8),
58959 => conv_std_logic_vector(70, 8),
58960 => conv_std_logic_vector(71, 8),
58961 => conv_std_logic_vector(72, 8),
58962 => conv_std_logic_vector(73, 8),
58963 => conv_std_logic_vector(74, 8),
58964 => conv_std_logic_vector(75, 8),
58965 => conv_std_logic_vector(76, 8),
58966 => conv_std_logic_vector(77, 8),
58967 => conv_std_logic_vector(78, 8),
58968 => conv_std_logic_vector(79, 8),
58969 => conv_std_logic_vector(79, 8),
58970 => conv_std_logic_vector(80, 8),
58971 => conv_std_logic_vector(81, 8),
58972 => conv_std_logic_vector(82, 8),
58973 => conv_std_logic_vector(83, 8),
58974 => conv_std_logic_vector(84, 8),
58975 => conv_std_logic_vector(85, 8),
58976 => conv_std_logic_vector(86, 8),
58977 => conv_std_logic_vector(87, 8),
58978 => conv_std_logic_vector(88, 8),
58979 => conv_std_logic_vector(88, 8),
58980 => conv_std_logic_vector(89, 8),
58981 => conv_std_logic_vector(90, 8),
58982 => conv_std_logic_vector(91, 8),
58983 => conv_std_logic_vector(92, 8),
58984 => conv_std_logic_vector(93, 8),
58985 => conv_std_logic_vector(94, 8),
58986 => conv_std_logic_vector(95, 8),
58987 => conv_std_logic_vector(96, 8),
58988 => conv_std_logic_vector(97, 8),
58989 => conv_std_logic_vector(97, 8),
58990 => conv_std_logic_vector(98, 8),
58991 => conv_std_logic_vector(99, 8),
58992 => conv_std_logic_vector(100, 8),
58993 => conv_std_logic_vector(101, 8),
58994 => conv_std_logic_vector(102, 8),
58995 => conv_std_logic_vector(103, 8),
58996 => conv_std_logic_vector(104, 8),
58997 => conv_std_logic_vector(105, 8),
58998 => conv_std_logic_vector(106, 8),
58999 => conv_std_logic_vector(106, 8),
59000 => conv_std_logic_vector(107, 8),
59001 => conv_std_logic_vector(108, 8),
59002 => conv_std_logic_vector(109, 8),
59003 => conv_std_logic_vector(110, 8),
59004 => conv_std_logic_vector(111, 8),
59005 => conv_std_logic_vector(112, 8),
59006 => conv_std_logic_vector(113, 8),
59007 => conv_std_logic_vector(114, 8),
59008 => conv_std_logic_vector(115, 8),
59009 => conv_std_logic_vector(115, 8),
59010 => conv_std_logic_vector(116, 8),
59011 => conv_std_logic_vector(117, 8),
59012 => conv_std_logic_vector(118, 8),
59013 => conv_std_logic_vector(119, 8),
59014 => conv_std_logic_vector(120, 8),
59015 => conv_std_logic_vector(121, 8),
59016 => conv_std_logic_vector(122, 8),
59017 => conv_std_logic_vector(123, 8),
59018 => conv_std_logic_vector(123, 8),
59019 => conv_std_logic_vector(124, 8),
59020 => conv_std_logic_vector(125, 8),
59021 => conv_std_logic_vector(126, 8),
59022 => conv_std_logic_vector(127, 8),
59023 => conv_std_logic_vector(128, 8),
59024 => conv_std_logic_vector(129, 8),
59025 => conv_std_logic_vector(130, 8),
59026 => conv_std_logic_vector(131, 8),
59027 => conv_std_logic_vector(132, 8),
59028 => conv_std_logic_vector(132, 8),
59029 => conv_std_logic_vector(133, 8),
59030 => conv_std_logic_vector(134, 8),
59031 => conv_std_logic_vector(135, 8),
59032 => conv_std_logic_vector(136, 8),
59033 => conv_std_logic_vector(137, 8),
59034 => conv_std_logic_vector(138, 8),
59035 => conv_std_logic_vector(139, 8),
59036 => conv_std_logic_vector(140, 8),
59037 => conv_std_logic_vector(141, 8),
59038 => conv_std_logic_vector(141, 8),
59039 => conv_std_logic_vector(142, 8),
59040 => conv_std_logic_vector(143, 8),
59041 => conv_std_logic_vector(144, 8),
59042 => conv_std_logic_vector(145, 8),
59043 => conv_std_logic_vector(146, 8),
59044 => conv_std_logic_vector(147, 8),
59045 => conv_std_logic_vector(148, 8),
59046 => conv_std_logic_vector(149, 8),
59047 => conv_std_logic_vector(150, 8),
59048 => conv_std_logic_vector(150, 8),
59049 => conv_std_logic_vector(151, 8),
59050 => conv_std_logic_vector(152, 8),
59051 => conv_std_logic_vector(153, 8),
59052 => conv_std_logic_vector(154, 8),
59053 => conv_std_logic_vector(155, 8),
59054 => conv_std_logic_vector(156, 8),
59055 => conv_std_logic_vector(157, 8),
59056 => conv_std_logic_vector(158, 8),
59057 => conv_std_logic_vector(159, 8),
59058 => conv_std_logic_vector(159, 8),
59059 => conv_std_logic_vector(160, 8),
59060 => conv_std_logic_vector(161, 8),
59061 => conv_std_logic_vector(162, 8),
59062 => conv_std_logic_vector(163, 8),
59063 => conv_std_logic_vector(164, 8),
59064 => conv_std_logic_vector(165, 8),
59065 => conv_std_logic_vector(166, 8),
59066 => conv_std_logic_vector(167, 8),
59067 => conv_std_logic_vector(168, 8),
59068 => conv_std_logic_vector(168, 8),
59069 => conv_std_logic_vector(169, 8),
59070 => conv_std_logic_vector(170, 8),
59071 => conv_std_logic_vector(171, 8),
59072 => conv_std_logic_vector(172, 8),
59073 => conv_std_logic_vector(173, 8),
59074 => conv_std_logic_vector(174, 8),
59075 => conv_std_logic_vector(175, 8),
59076 => conv_std_logic_vector(176, 8),
59077 => conv_std_logic_vector(176, 8),
59078 => conv_std_logic_vector(177, 8),
59079 => conv_std_logic_vector(178, 8),
59080 => conv_std_logic_vector(179, 8),
59081 => conv_std_logic_vector(180, 8),
59082 => conv_std_logic_vector(181, 8),
59083 => conv_std_logic_vector(182, 8),
59084 => conv_std_logic_vector(183, 8),
59085 => conv_std_logic_vector(184, 8),
59086 => conv_std_logic_vector(185, 8),
59087 => conv_std_logic_vector(185, 8),
59088 => conv_std_logic_vector(186, 8),
59089 => conv_std_logic_vector(187, 8),
59090 => conv_std_logic_vector(188, 8),
59091 => conv_std_logic_vector(189, 8),
59092 => conv_std_logic_vector(190, 8),
59093 => conv_std_logic_vector(191, 8),
59094 => conv_std_logic_vector(192, 8),
59095 => conv_std_logic_vector(193, 8),
59096 => conv_std_logic_vector(194, 8),
59097 => conv_std_logic_vector(194, 8),
59098 => conv_std_logic_vector(195, 8),
59099 => conv_std_logic_vector(196, 8),
59100 => conv_std_logic_vector(197, 8),
59101 => conv_std_logic_vector(198, 8),
59102 => conv_std_logic_vector(199, 8),
59103 => conv_std_logic_vector(200, 8),
59104 => conv_std_logic_vector(201, 8),
59105 => conv_std_logic_vector(202, 8),
59106 => conv_std_logic_vector(203, 8),
59107 => conv_std_logic_vector(203, 8),
59108 => conv_std_logic_vector(204, 8),
59109 => conv_std_logic_vector(205, 8),
59110 => conv_std_logic_vector(206, 8),
59111 => conv_std_logic_vector(207, 8),
59112 => conv_std_logic_vector(208, 8),
59113 => conv_std_logic_vector(209, 8),
59114 => conv_std_logic_vector(210, 8),
59115 => conv_std_logic_vector(211, 8),
59116 => conv_std_logic_vector(212, 8),
59117 => conv_std_logic_vector(212, 8),
59118 => conv_std_logic_vector(213, 8),
59119 => conv_std_logic_vector(214, 8),
59120 => conv_std_logic_vector(215, 8),
59121 => conv_std_logic_vector(216, 8),
59122 => conv_std_logic_vector(217, 8),
59123 => conv_std_logic_vector(218, 8),
59124 => conv_std_logic_vector(219, 8),
59125 => conv_std_logic_vector(220, 8),
59126 => conv_std_logic_vector(221, 8),
59127 => conv_std_logic_vector(221, 8),
59128 => conv_std_logic_vector(222, 8),
59129 => conv_std_logic_vector(223, 8),
59130 => conv_std_logic_vector(224, 8),
59131 => conv_std_logic_vector(225, 8),
59132 => conv_std_logic_vector(226, 8),
59133 => conv_std_logic_vector(227, 8),
59134 => conv_std_logic_vector(228, 8),
59135 => conv_std_logic_vector(229, 8),
59136 => conv_std_logic_vector(0, 8),
59137 => conv_std_logic_vector(0, 8),
59138 => conv_std_logic_vector(1, 8),
59139 => conv_std_logic_vector(2, 8),
59140 => conv_std_logic_vector(3, 8),
59141 => conv_std_logic_vector(4, 8),
59142 => conv_std_logic_vector(5, 8),
59143 => conv_std_logic_vector(6, 8),
59144 => conv_std_logic_vector(7, 8),
59145 => conv_std_logic_vector(8, 8),
59146 => conv_std_logic_vector(9, 8),
59147 => conv_std_logic_vector(9, 8),
59148 => conv_std_logic_vector(10, 8),
59149 => conv_std_logic_vector(11, 8),
59150 => conv_std_logic_vector(12, 8),
59151 => conv_std_logic_vector(13, 8),
59152 => conv_std_logic_vector(14, 8),
59153 => conv_std_logic_vector(15, 8),
59154 => conv_std_logic_vector(16, 8),
59155 => conv_std_logic_vector(17, 8),
59156 => conv_std_logic_vector(18, 8),
59157 => conv_std_logic_vector(18, 8),
59158 => conv_std_logic_vector(19, 8),
59159 => conv_std_logic_vector(20, 8),
59160 => conv_std_logic_vector(21, 8),
59161 => conv_std_logic_vector(22, 8),
59162 => conv_std_logic_vector(23, 8),
59163 => conv_std_logic_vector(24, 8),
59164 => conv_std_logic_vector(25, 8),
59165 => conv_std_logic_vector(26, 8),
59166 => conv_std_logic_vector(27, 8),
59167 => conv_std_logic_vector(27, 8),
59168 => conv_std_logic_vector(28, 8),
59169 => conv_std_logic_vector(29, 8),
59170 => conv_std_logic_vector(30, 8),
59171 => conv_std_logic_vector(31, 8),
59172 => conv_std_logic_vector(32, 8),
59173 => conv_std_logic_vector(33, 8),
59174 => conv_std_logic_vector(34, 8),
59175 => conv_std_logic_vector(35, 8),
59176 => conv_std_logic_vector(36, 8),
59177 => conv_std_logic_vector(36, 8),
59178 => conv_std_logic_vector(37, 8),
59179 => conv_std_logic_vector(38, 8),
59180 => conv_std_logic_vector(39, 8),
59181 => conv_std_logic_vector(40, 8),
59182 => conv_std_logic_vector(41, 8),
59183 => conv_std_logic_vector(42, 8),
59184 => conv_std_logic_vector(43, 8),
59185 => conv_std_logic_vector(44, 8),
59186 => conv_std_logic_vector(45, 8),
59187 => conv_std_logic_vector(46, 8),
59188 => conv_std_logic_vector(46, 8),
59189 => conv_std_logic_vector(47, 8),
59190 => conv_std_logic_vector(48, 8),
59191 => conv_std_logic_vector(49, 8),
59192 => conv_std_logic_vector(50, 8),
59193 => conv_std_logic_vector(51, 8),
59194 => conv_std_logic_vector(52, 8),
59195 => conv_std_logic_vector(53, 8),
59196 => conv_std_logic_vector(54, 8),
59197 => conv_std_logic_vector(55, 8),
59198 => conv_std_logic_vector(55, 8),
59199 => conv_std_logic_vector(56, 8),
59200 => conv_std_logic_vector(57, 8),
59201 => conv_std_logic_vector(58, 8),
59202 => conv_std_logic_vector(59, 8),
59203 => conv_std_logic_vector(60, 8),
59204 => conv_std_logic_vector(61, 8),
59205 => conv_std_logic_vector(62, 8),
59206 => conv_std_logic_vector(63, 8),
59207 => conv_std_logic_vector(64, 8),
59208 => conv_std_logic_vector(64, 8),
59209 => conv_std_logic_vector(65, 8),
59210 => conv_std_logic_vector(66, 8),
59211 => conv_std_logic_vector(67, 8),
59212 => conv_std_logic_vector(68, 8),
59213 => conv_std_logic_vector(69, 8),
59214 => conv_std_logic_vector(70, 8),
59215 => conv_std_logic_vector(71, 8),
59216 => conv_std_logic_vector(72, 8),
59217 => conv_std_logic_vector(73, 8),
59218 => conv_std_logic_vector(73, 8),
59219 => conv_std_logic_vector(74, 8),
59220 => conv_std_logic_vector(75, 8),
59221 => conv_std_logic_vector(76, 8),
59222 => conv_std_logic_vector(77, 8),
59223 => conv_std_logic_vector(78, 8),
59224 => conv_std_logic_vector(79, 8),
59225 => conv_std_logic_vector(80, 8),
59226 => conv_std_logic_vector(81, 8),
59227 => conv_std_logic_vector(82, 8),
59228 => conv_std_logic_vector(83, 8),
59229 => conv_std_logic_vector(83, 8),
59230 => conv_std_logic_vector(84, 8),
59231 => conv_std_logic_vector(85, 8),
59232 => conv_std_logic_vector(86, 8),
59233 => conv_std_logic_vector(87, 8),
59234 => conv_std_logic_vector(88, 8),
59235 => conv_std_logic_vector(89, 8),
59236 => conv_std_logic_vector(90, 8),
59237 => conv_std_logic_vector(91, 8),
59238 => conv_std_logic_vector(92, 8),
59239 => conv_std_logic_vector(92, 8),
59240 => conv_std_logic_vector(93, 8),
59241 => conv_std_logic_vector(94, 8),
59242 => conv_std_logic_vector(95, 8),
59243 => conv_std_logic_vector(96, 8),
59244 => conv_std_logic_vector(97, 8),
59245 => conv_std_logic_vector(98, 8),
59246 => conv_std_logic_vector(99, 8),
59247 => conv_std_logic_vector(100, 8),
59248 => conv_std_logic_vector(101, 8),
59249 => conv_std_logic_vector(101, 8),
59250 => conv_std_logic_vector(102, 8),
59251 => conv_std_logic_vector(103, 8),
59252 => conv_std_logic_vector(104, 8),
59253 => conv_std_logic_vector(105, 8),
59254 => conv_std_logic_vector(106, 8),
59255 => conv_std_logic_vector(107, 8),
59256 => conv_std_logic_vector(108, 8),
59257 => conv_std_logic_vector(109, 8),
59258 => conv_std_logic_vector(110, 8),
59259 => conv_std_logic_vector(110, 8),
59260 => conv_std_logic_vector(111, 8),
59261 => conv_std_logic_vector(112, 8),
59262 => conv_std_logic_vector(113, 8),
59263 => conv_std_logic_vector(114, 8),
59264 => conv_std_logic_vector(115, 8),
59265 => conv_std_logic_vector(116, 8),
59266 => conv_std_logic_vector(117, 8),
59267 => conv_std_logic_vector(118, 8),
59268 => conv_std_logic_vector(119, 8),
59269 => conv_std_logic_vector(120, 8),
59270 => conv_std_logic_vector(120, 8),
59271 => conv_std_logic_vector(121, 8),
59272 => conv_std_logic_vector(122, 8),
59273 => conv_std_logic_vector(123, 8),
59274 => conv_std_logic_vector(124, 8),
59275 => conv_std_logic_vector(125, 8),
59276 => conv_std_logic_vector(126, 8),
59277 => conv_std_logic_vector(127, 8),
59278 => conv_std_logic_vector(128, 8),
59279 => conv_std_logic_vector(129, 8),
59280 => conv_std_logic_vector(129, 8),
59281 => conv_std_logic_vector(130, 8),
59282 => conv_std_logic_vector(131, 8),
59283 => conv_std_logic_vector(132, 8),
59284 => conv_std_logic_vector(133, 8),
59285 => conv_std_logic_vector(134, 8),
59286 => conv_std_logic_vector(135, 8),
59287 => conv_std_logic_vector(136, 8),
59288 => conv_std_logic_vector(137, 8),
59289 => conv_std_logic_vector(138, 8),
59290 => conv_std_logic_vector(138, 8),
59291 => conv_std_logic_vector(139, 8),
59292 => conv_std_logic_vector(140, 8),
59293 => conv_std_logic_vector(141, 8),
59294 => conv_std_logic_vector(142, 8),
59295 => conv_std_logic_vector(143, 8),
59296 => conv_std_logic_vector(144, 8),
59297 => conv_std_logic_vector(145, 8),
59298 => conv_std_logic_vector(146, 8),
59299 => conv_std_logic_vector(147, 8),
59300 => conv_std_logic_vector(147, 8),
59301 => conv_std_logic_vector(148, 8),
59302 => conv_std_logic_vector(149, 8),
59303 => conv_std_logic_vector(150, 8),
59304 => conv_std_logic_vector(151, 8),
59305 => conv_std_logic_vector(152, 8),
59306 => conv_std_logic_vector(153, 8),
59307 => conv_std_logic_vector(154, 8),
59308 => conv_std_logic_vector(155, 8),
59309 => conv_std_logic_vector(156, 8),
59310 => conv_std_logic_vector(157, 8),
59311 => conv_std_logic_vector(157, 8),
59312 => conv_std_logic_vector(158, 8),
59313 => conv_std_logic_vector(159, 8),
59314 => conv_std_logic_vector(160, 8),
59315 => conv_std_logic_vector(161, 8),
59316 => conv_std_logic_vector(162, 8),
59317 => conv_std_logic_vector(163, 8),
59318 => conv_std_logic_vector(164, 8),
59319 => conv_std_logic_vector(165, 8),
59320 => conv_std_logic_vector(166, 8),
59321 => conv_std_logic_vector(166, 8),
59322 => conv_std_logic_vector(167, 8),
59323 => conv_std_logic_vector(168, 8),
59324 => conv_std_logic_vector(169, 8),
59325 => conv_std_logic_vector(170, 8),
59326 => conv_std_logic_vector(171, 8),
59327 => conv_std_logic_vector(172, 8),
59328 => conv_std_logic_vector(173, 8),
59329 => conv_std_logic_vector(174, 8),
59330 => conv_std_logic_vector(175, 8),
59331 => conv_std_logic_vector(175, 8),
59332 => conv_std_logic_vector(176, 8),
59333 => conv_std_logic_vector(177, 8),
59334 => conv_std_logic_vector(178, 8),
59335 => conv_std_logic_vector(179, 8),
59336 => conv_std_logic_vector(180, 8),
59337 => conv_std_logic_vector(181, 8),
59338 => conv_std_logic_vector(182, 8),
59339 => conv_std_logic_vector(183, 8),
59340 => conv_std_logic_vector(184, 8),
59341 => conv_std_logic_vector(184, 8),
59342 => conv_std_logic_vector(185, 8),
59343 => conv_std_logic_vector(186, 8),
59344 => conv_std_logic_vector(187, 8),
59345 => conv_std_logic_vector(188, 8),
59346 => conv_std_logic_vector(189, 8),
59347 => conv_std_logic_vector(190, 8),
59348 => conv_std_logic_vector(191, 8),
59349 => conv_std_logic_vector(192, 8),
59350 => conv_std_logic_vector(193, 8),
59351 => conv_std_logic_vector(194, 8),
59352 => conv_std_logic_vector(194, 8),
59353 => conv_std_logic_vector(195, 8),
59354 => conv_std_logic_vector(196, 8),
59355 => conv_std_logic_vector(197, 8),
59356 => conv_std_logic_vector(198, 8),
59357 => conv_std_logic_vector(199, 8),
59358 => conv_std_logic_vector(200, 8),
59359 => conv_std_logic_vector(201, 8),
59360 => conv_std_logic_vector(202, 8),
59361 => conv_std_logic_vector(203, 8),
59362 => conv_std_logic_vector(203, 8),
59363 => conv_std_logic_vector(204, 8),
59364 => conv_std_logic_vector(205, 8),
59365 => conv_std_logic_vector(206, 8),
59366 => conv_std_logic_vector(207, 8),
59367 => conv_std_logic_vector(208, 8),
59368 => conv_std_logic_vector(209, 8),
59369 => conv_std_logic_vector(210, 8),
59370 => conv_std_logic_vector(211, 8),
59371 => conv_std_logic_vector(212, 8),
59372 => conv_std_logic_vector(212, 8),
59373 => conv_std_logic_vector(213, 8),
59374 => conv_std_logic_vector(214, 8),
59375 => conv_std_logic_vector(215, 8),
59376 => conv_std_logic_vector(216, 8),
59377 => conv_std_logic_vector(217, 8),
59378 => conv_std_logic_vector(218, 8),
59379 => conv_std_logic_vector(219, 8),
59380 => conv_std_logic_vector(220, 8),
59381 => conv_std_logic_vector(221, 8),
59382 => conv_std_logic_vector(221, 8),
59383 => conv_std_logic_vector(222, 8),
59384 => conv_std_logic_vector(223, 8),
59385 => conv_std_logic_vector(224, 8),
59386 => conv_std_logic_vector(225, 8),
59387 => conv_std_logic_vector(226, 8),
59388 => conv_std_logic_vector(227, 8),
59389 => conv_std_logic_vector(228, 8),
59390 => conv_std_logic_vector(229, 8),
59391 => conv_std_logic_vector(230, 8),
59392 => conv_std_logic_vector(0, 8),
59393 => conv_std_logic_vector(0, 8),
59394 => conv_std_logic_vector(1, 8),
59395 => conv_std_logic_vector(2, 8),
59396 => conv_std_logic_vector(3, 8),
59397 => conv_std_logic_vector(4, 8),
59398 => conv_std_logic_vector(5, 8),
59399 => conv_std_logic_vector(6, 8),
59400 => conv_std_logic_vector(7, 8),
59401 => conv_std_logic_vector(8, 8),
59402 => conv_std_logic_vector(9, 8),
59403 => conv_std_logic_vector(9, 8),
59404 => conv_std_logic_vector(10, 8),
59405 => conv_std_logic_vector(11, 8),
59406 => conv_std_logic_vector(12, 8),
59407 => conv_std_logic_vector(13, 8),
59408 => conv_std_logic_vector(14, 8),
59409 => conv_std_logic_vector(15, 8),
59410 => conv_std_logic_vector(16, 8),
59411 => conv_std_logic_vector(17, 8),
59412 => conv_std_logic_vector(18, 8),
59413 => conv_std_logic_vector(19, 8),
59414 => conv_std_logic_vector(19, 8),
59415 => conv_std_logic_vector(20, 8),
59416 => conv_std_logic_vector(21, 8),
59417 => conv_std_logic_vector(22, 8),
59418 => conv_std_logic_vector(23, 8),
59419 => conv_std_logic_vector(24, 8),
59420 => conv_std_logic_vector(25, 8),
59421 => conv_std_logic_vector(26, 8),
59422 => conv_std_logic_vector(27, 8),
59423 => conv_std_logic_vector(28, 8),
59424 => conv_std_logic_vector(29, 8),
59425 => conv_std_logic_vector(29, 8),
59426 => conv_std_logic_vector(30, 8),
59427 => conv_std_logic_vector(31, 8),
59428 => conv_std_logic_vector(32, 8),
59429 => conv_std_logic_vector(33, 8),
59430 => conv_std_logic_vector(34, 8),
59431 => conv_std_logic_vector(35, 8),
59432 => conv_std_logic_vector(36, 8),
59433 => conv_std_logic_vector(37, 8),
59434 => conv_std_logic_vector(38, 8),
59435 => conv_std_logic_vector(38, 8),
59436 => conv_std_logic_vector(39, 8),
59437 => conv_std_logic_vector(40, 8),
59438 => conv_std_logic_vector(41, 8),
59439 => conv_std_logic_vector(42, 8),
59440 => conv_std_logic_vector(43, 8),
59441 => conv_std_logic_vector(44, 8),
59442 => conv_std_logic_vector(45, 8),
59443 => conv_std_logic_vector(46, 8),
59444 => conv_std_logic_vector(47, 8),
59445 => conv_std_logic_vector(48, 8),
59446 => conv_std_logic_vector(48, 8),
59447 => conv_std_logic_vector(49, 8),
59448 => conv_std_logic_vector(50, 8),
59449 => conv_std_logic_vector(51, 8),
59450 => conv_std_logic_vector(52, 8),
59451 => conv_std_logic_vector(53, 8),
59452 => conv_std_logic_vector(54, 8),
59453 => conv_std_logic_vector(55, 8),
59454 => conv_std_logic_vector(56, 8),
59455 => conv_std_logic_vector(57, 8),
59456 => conv_std_logic_vector(58, 8),
59457 => conv_std_logic_vector(58, 8),
59458 => conv_std_logic_vector(59, 8),
59459 => conv_std_logic_vector(60, 8),
59460 => conv_std_logic_vector(61, 8),
59461 => conv_std_logic_vector(62, 8),
59462 => conv_std_logic_vector(63, 8),
59463 => conv_std_logic_vector(64, 8),
59464 => conv_std_logic_vector(65, 8),
59465 => conv_std_logic_vector(66, 8),
59466 => conv_std_logic_vector(67, 8),
59467 => conv_std_logic_vector(67, 8),
59468 => conv_std_logic_vector(68, 8),
59469 => conv_std_logic_vector(69, 8),
59470 => conv_std_logic_vector(70, 8),
59471 => conv_std_logic_vector(71, 8),
59472 => conv_std_logic_vector(72, 8),
59473 => conv_std_logic_vector(73, 8),
59474 => conv_std_logic_vector(74, 8),
59475 => conv_std_logic_vector(75, 8),
59476 => conv_std_logic_vector(76, 8),
59477 => conv_std_logic_vector(77, 8),
59478 => conv_std_logic_vector(77, 8),
59479 => conv_std_logic_vector(78, 8),
59480 => conv_std_logic_vector(79, 8),
59481 => conv_std_logic_vector(80, 8),
59482 => conv_std_logic_vector(81, 8),
59483 => conv_std_logic_vector(82, 8),
59484 => conv_std_logic_vector(83, 8),
59485 => conv_std_logic_vector(84, 8),
59486 => conv_std_logic_vector(85, 8),
59487 => conv_std_logic_vector(86, 8),
59488 => conv_std_logic_vector(87, 8),
59489 => conv_std_logic_vector(87, 8),
59490 => conv_std_logic_vector(88, 8),
59491 => conv_std_logic_vector(89, 8),
59492 => conv_std_logic_vector(90, 8),
59493 => conv_std_logic_vector(91, 8),
59494 => conv_std_logic_vector(92, 8),
59495 => conv_std_logic_vector(93, 8),
59496 => conv_std_logic_vector(94, 8),
59497 => conv_std_logic_vector(95, 8),
59498 => conv_std_logic_vector(96, 8),
59499 => conv_std_logic_vector(96, 8),
59500 => conv_std_logic_vector(97, 8),
59501 => conv_std_logic_vector(98, 8),
59502 => conv_std_logic_vector(99, 8),
59503 => conv_std_logic_vector(100, 8),
59504 => conv_std_logic_vector(101, 8),
59505 => conv_std_logic_vector(102, 8),
59506 => conv_std_logic_vector(103, 8),
59507 => conv_std_logic_vector(104, 8),
59508 => conv_std_logic_vector(105, 8),
59509 => conv_std_logic_vector(106, 8),
59510 => conv_std_logic_vector(106, 8),
59511 => conv_std_logic_vector(107, 8),
59512 => conv_std_logic_vector(108, 8),
59513 => conv_std_logic_vector(109, 8),
59514 => conv_std_logic_vector(110, 8),
59515 => conv_std_logic_vector(111, 8),
59516 => conv_std_logic_vector(112, 8),
59517 => conv_std_logic_vector(113, 8),
59518 => conv_std_logic_vector(114, 8),
59519 => conv_std_logic_vector(115, 8),
59520 => conv_std_logic_vector(116, 8),
59521 => conv_std_logic_vector(116, 8),
59522 => conv_std_logic_vector(117, 8),
59523 => conv_std_logic_vector(118, 8),
59524 => conv_std_logic_vector(119, 8),
59525 => conv_std_logic_vector(120, 8),
59526 => conv_std_logic_vector(121, 8),
59527 => conv_std_logic_vector(122, 8),
59528 => conv_std_logic_vector(123, 8),
59529 => conv_std_logic_vector(124, 8),
59530 => conv_std_logic_vector(125, 8),
59531 => conv_std_logic_vector(125, 8),
59532 => conv_std_logic_vector(126, 8),
59533 => conv_std_logic_vector(127, 8),
59534 => conv_std_logic_vector(128, 8),
59535 => conv_std_logic_vector(129, 8),
59536 => conv_std_logic_vector(130, 8),
59537 => conv_std_logic_vector(131, 8),
59538 => conv_std_logic_vector(132, 8),
59539 => conv_std_logic_vector(133, 8),
59540 => conv_std_logic_vector(134, 8),
59541 => conv_std_logic_vector(135, 8),
59542 => conv_std_logic_vector(135, 8),
59543 => conv_std_logic_vector(136, 8),
59544 => conv_std_logic_vector(137, 8),
59545 => conv_std_logic_vector(138, 8),
59546 => conv_std_logic_vector(139, 8),
59547 => conv_std_logic_vector(140, 8),
59548 => conv_std_logic_vector(141, 8),
59549 => conv_std_logic_vector(142, 8),
59550 => conv_std_logic_vector(143, 8),
59551 => conv_std_logic_vector(144, 8),
59552 => conv_std_logic_vector(145, 8),
59553 => conv_std_logic_vector(145, 8),
59554 => conv_std_logic_vector(146, 8),
59555 => conv_std_logic_vector(147, 8),
59556 => conv_std_logic_vector(148, 8),
59557 => conv_std_logic_vector(149, 8),
59558 => conv_std_logic_vector(150, 8),
59559 => conv_std_logic_vector(151, 8),
59560 => conv_std_logic_vector(152, 8),
59561 => conv_std_logic_vector(153, 8),
59562 => conv_std_logic_vector(154, 8),
59563 => conv_std_logic_vector(154, 8),
59564 => conv_std_logic_vector(155, 8),
59565 => conv_std_logic_vector(156, 8),
59566 => conv_std_logic_vector(157, 8),
59567 => conv_std_logic_vector(158, 8),
59568 => conv_std_logic_vector(159, 8),
59569 => conv_std_logic_vector(160, 8),
59570 => conv_std_logic_vector(161, 8),
59571 => conv_std_logic_vector(162, 8),
59572 => conv_std_logic_vector(163, 8),
59573 => conv_std_logic_vector(164, 8),
59574 => conv_std_logic_vector(164, 8),
59575 => conv_std_logic_vector(165, 8),
59576 => conv_std_logic_vector(166, 8),
59577 => conv_std_logic_vector(167, 8),
59578 => conv_std_logic_vector(168, 8),
59579 => conv_std_logic_vector(169, 8),
59580 => conv_std_logic_vector(170, 8),
59581 => conv_std_logic_vector(171, 8),
59582 => conv_std_logic_vector(172, 8),
59583 => conv_std_logic_vector(173, 8),
59584 => conv_std_logic_vector(174, 8),
59585 => conv_std_logic_vector(174, 8),
59586 => conv_std_logic_vector(175, 8),
59587 => conv_std_logic_vector(176, 8),
59588 => conv_std_logic_vector(177, 8),
59589 => conv_std_logic_vector(178, 8),
59590 => conv_std_logic_vector(179, 8),
59591 => conv_std_logic_vector(180, 8),
59592 => conv_std_logic_vector(181, 8),
59593 => conv_std_logic_vector(182, 8),
59594 => conv_std_logic_vector(183, 8),
59595 => conv_std_logic_vector(183, 8),
59596 => conv_std_logic_vector(184, 8),
59597 => conv_std_logic_vector(185, 8),
59598 => conv_std_logic_vector(186, 8),
59599 => conv_std_logic_vector(187, 8),
59600 => conv_std_logic_vector(188, 8),
59601 => conv_std_logic_vector(189, 8),
59602 => conv_std_logic_vector(190, 8),
59603 => conv_std_logic_vector(191, 8),
59604 => conv_std_logic_vector(192, 8),
59605 => conv_std_logic_vector(193, 8),
59606 => conv_std_logic_vector(193, 8),
59607 => conv_std_logic_vector(194, 8),
59608 => conv_std_logic_vector(195, 8),
59609 => conv_std_logic_vector(196, 8),
59610 => conv_std_logic_vector(197, 8),
59611 => conv_std_logic_vector(198, 8),
59612 => conv_std_logic_vector(199, 8),
59613 => conv_std_logic_vector(200, 8),
59614 => conv_std_logic_vector(201, 8),
59615 => conv_std_logic_vector(202, 8),
59616 => conv_std_logic_vector(203, 8),
59617 => conv_std_logic_vector(203, 8),
59618 => conv_std_logic_vector(204, 8),
59619 => conv_std_logic_vector(205, 8),
59620 => conv_std_logic_vector(206, 8),
59621 => conv_std_logic_vector(207, 8),
59622 => conv_std_logic_vector(208, 8),
59623 => conv_std_logic_vector(209, 8),
59624 => conv_std_logic_vector(210, 8),
59625 => conv_std_logic_vector(211, 8),
59626 => conv_std_logic_vector(212, 8),
59627 => conv_std_logic_vector(212, 8),
59628 => conv_std_logic_vector(213, 8),
59629 => conv_std_logic_vector(214, 8),
59630 => conv_std_logic_vector(215, 8),
59631 => conv_std_logic_vector(216, 8),
59632 => conv_std_logic_vector(217, 8),
59633 => conv_std_logic_vector(218, 8),
59634 => conv_std_logic_vector(219, 8),
59635 => conv_std_logic_vector(220, 8),
59636 => conv_std_logic_vector(221, 8),
59637 => conv_std_logic_vector(222, 8),
59638 => conv_std_logic_vector(222, 8),
59639 => conv_std_logic_vector(223, 8),
59640 => conv_std_logic_vector(224, 8),
59641 => conv_std_logic_vector(225, 8),
59642 => conv_std_logic_vector(226, 8),
59643 => conv_std_logic_vector(227, 8),
59644 => conv_std_logic_vector(228, 8),
59645 => conv_std_logic_vector(229, 8),
59646 => conv_std_logic_vector(230, 8),
59647 => conv_std_logic_vector(231, 8),
59648 => conv_std_logic_vector(0, 8),
59649 => conv_std_logic_vector(0, 8),
59650 => conv_std_logic_vector(1, 8),
59651 => conv_std_logic_vector(2, 8),
59652 => conv_std_logic_vector(3, 8),
59653 => conv_std_logic_vector(4, 8),
59654 => conv_std_logic_vector(5, 8),
59655 => conv_std_logic_vector(6, 8),
59656 => conv_std_logic_vector(7, 8),
59657 => conv_std_logic_vector(8, 8),
59658 => conv_std_logic_vector(9, 8),
59659 => conv_std_logic_vector(10, 8),
59660 => conv_std_logic_vector(10, 8),
59661 => conv_std_logic_vector(11, 8),
59662 => conv_std_logic_vector(12, 8),
59663 => conv_std_logic_vector(13, 8),
59664 => conv_std_logic_vector(14, 8),
59665 => conv_std_logic_vector(15, 8),
59666 => conv_std_logic_vector(16, 8),
59667 => conv_std_logic_vector(17, 8),
59668 => conv_std_logic_vector(18, 8),
59669 => conv_std_logic_vector(19, 8),
59670 => conv_std_logic_vector(20, 8),
59671 => conv_std_logic_vector(20, 8),
59672 => conv_std_logic_vector(21, 8),
59673 => conv_std_logic_vector(22, 8),
59674 => conv_std_logic_vector(23, 8),
59675 => conv_std_logic_vector(24, 8),
59676 => conv_std_logic_vector(25, 8),
59677 => conv_std_logic_vector(26, 8),
59678 => conv_std_logic_vector(27, 8),
59679 => conv_std_logic_vector(28, 8),
59680 => conv_std_logic_vector(29, 8),
59681 => conv_std_logic_vector(30, 8),
59682 => conv_std_logic_vector(30, 8),
59683 => conv_std_logic_vector(31, 8),
59684 => conv_std_logic_vector(32, 8),
59685 => conv_std_logic_vector(33, 8),
59686 => conv_std_logic_vector(34, 8),
59687 => conv_std_logic_vector(35, 8),
59688 => conv_std_logic_vector(36, 8),
59689 => conv_std_logic_vector(37, 8),
59690 => conv_std_logic_vector(38, 8),
59691 => conv_std_logic_vector(39, 8),
59692 => conv_std_logic_vector(40, 8),
59693 => conv_std_logic_vector(40, 8),
59694 => conv_std_logic_vector(41, 8),
59695 => conv_std_logic_vector(42, 8),
59696 => conv_std_logic_vector(43, 8),
59697 => conv_std_logic_vector(44, 8),
59698 => conv_std_logic_vector(45, 8),
59699 => conv_std_logic_vector(46, 8),
59700 => conv_std_logic_vector(47, 8),
59701 => conv_std_logic_vector(48, 8),
59702 => conv_std_logic_vector(49, 8),
59703 => conv_std_logic_vector(50, 8),
59704 => conv_std_logic_vector(50, 8),
59705 => conv_std_logic_vector(51, 8),
59706 => conv_std_logic_vector(52, 8),
59707 => conv_std_logic_vector(53, 8),
59708 => conv_std_logic_vector(54, 8),
59709 => conv_std_logic_vector(55, 8),
59710 => conv_std_logic_vector(56, 8),
59711 => conv_std_logic_vector(57, 8),
59712 => conv_std_logic_vector(58, 8),
59713 => conv_std_logic_vector(59, 8),
59714 => conv_std_logic_vector(60, 8),
59715 => conv_std_logic_vector(60, 8),
59716 => conv_std_logic_vector(61, 8),
59717 => conv_std_logic_vector(62, 8),
59718 => conv_std_logic_vector(63, 8),
59719 => conv_std_logic_vector(64, 8),
59720 => conv_std_logic_vector(65, 8),
59721 => conv_std_logic_vector(66, 8),
59722 => conv_std_logic_vector(67, 8),
59723 => conv_std_logic_vector(68, 8),
59724 => conv_std_logic_vector(69, 8),
59725 => conv_std_logic_vector(70, 8),
59726 => conv_std_logic_vector(70, 8),
59727 => conv_std_logic_vector(71, 8),
59728 => conv_std_logic_vector(72, 8),
59729 => conv_std_logic_vector(73, 8),
59730 => conv_std_logic_vector(74, 8),
59731 => conv_std_logic_vector(75, 8),
59732 => conv_std_logic_vector(76, 8),
59733 => conv_std_logic_vector(77, 8),
59734 => conv_std_logic_vector(78, 8),
59735 => conv_std_logic_vector(79, 8),
59736 => conv_std_logic_vector(80, 8),
59737 => conv_std_logic_vector(81, 8),
59738 => conv_std_logic_vector(81, 8),
59739 => conv_std_logic_vector(82, 8),
59740 => conv_std_logic_vector(83, 8),
59741 => conv_std_logic_vector(84, 8),
59742 => conv_std_logic_vector(85, 8),
59743 => conv_std_logic_vector(86, 8),
59744 => conv_std_logic_vector(87, 8),
59745 => conv_std_logic_vector(88, 8),
59746 => conv_std_logic_vector(89, 8),
59747 => conv_std_logic_vector(90, 8),
59748 => conv_std_logic_vector(91, 8),
59749 => conv_std_logic_vector(91, 8),
59750 => conv_std_logic_vector(92, 8),
59751 => conv_std_logic_vector(93, 8),
59752 => conv_std_logic_vector(94, 8),
59753 => conv_std_logic_vector(95, 8),
59754 => conv_std_logic_vector(96, 8),
59755 => conv_std_logic_vector(97, 8),
59756 => conv_std_logic_vector(98, 8),
59757 => conv_std_logic_vector(99, 8),
59758 => conv_std_logic_vector(100, 8),
59759 => conv_std_logic_vector(101, 8),
59760 => conv_std_logic_vector(101, 8),
59761 => conv_std_logic_vector(102, 8),
59762 => conv_std_logic_vector(103, 8),
59763 => conv_std_logic_vector(104, 8),
59764 => conv_std_logic_vector(105, 8),
59765 => conv_std_logic_vector(106, 8),
59766 => conv_std_logic_vector(107, 8),
59767 => conv_std_logic_vector(108, 8),
59768 => conv_std_logic_vector(109, 8),
59769 => conv_std_logic_vector(110, 8),
59770 => conv_std_logic_vector(111, 8),
59771 => conv_std_logic_vector(111, 8),
59772 => conv_std_logic_vector(112, 8),
59773 => conv_std_logic_vector(113, 8),
59774 => conv_std_logic_vector(114, 8),
59775 => conv_std_logic_vector(115, 8),
59776 => conv_std_logic_vector(116, 8),
59777 => conv_std_logic_vector(117, 8),
59778 => conv_std_logic_vector(118, 8),
59779 => conv_std_logic_vector(119, 8),
59780 => conv_std_logic_vector(120, 8),
59781 => conv_std_logic_vector(121, 8),
59782 => conv_std_logic_vector(121, 8),
59783 => conv_std_logic_vector(122, 8),
59784 => conv_std_logic_vector(123, 8),
59785 => conv_std_logic_vector(124, 8),
59786 => conv_std_logic_vector(125, 8),
59787 => conv_std_logic_vector(126, 8),
59788 => conv_std_logic_vector(127, 8),
59789 => conv_std_logic_vector(128, 8),
59790 => conv_std_logic_vector(129, 8),
59791 => conv_std_logic_vector(130, 8),
59792 => conv_std_logic_vector(131, 8),
59793 => conv_std_logic_vector(131, 8),
59794 => conv_std_logic_vector(132, 8),
59795 => conv_std_logic_vector(133, 8),
59796 => conv_std_logic_vector(134, 8),
59797 => conv_std_logic_vector(135, 8),
59798 => conv_std_logic_vector(136, 8),
59799 => conv_std_logic_vector(137, 8),
59800 => conv_std_logic_vector(138, 8),
59801 => conv_std_logic_vector(139, 8),
59802 => conv_std_logic_vector(140, 8),
59803 => conv_std_logic_vector(141, 8),
59804 => conv_std_logic_vector(141, 8),
59805 => conv_std_logic_vector(142, 8),
59806 => conv_std_logic_vector(143, 8),
59807 => conv_std_logic_vector(144, 8),
59808 => conv_std_logic_vector(145, 8),
59809 => conv_std_logic_vector(146, 8),
59810 => conv_std_logic_vector(147, 8),
59811 => conv_std_logic_vector(148, 8),
59812 => conv_std_logic_vector(149, 8),
59813 => conv_std_logic_vector(150, 8),
59814 => conv_std_logic_vector(151, 8),
59815 => conv_std_logic_vector(151, 8),
59816 => conv_std_logic_vector(152, 8),
59817 => conv_std_logic_vector(153, 8),
59818 => conv_std_logic_vector(154, 8),
59819 => conv_std_logic_vector(155, 8),
59820 => conv_std_logic_vector(156, 8),
59821 => conv_std_logic_vector(157, 8),
59822 => conv_std_logic_vector(158, 8),
59823 => conv_std_logic_vector(159, 8),
59824 => conv_std_logic_vector(160, 8),
59825 => conv_std_logic_vector(161, 8),
59826 => conv_std_logic_vector(162, 8),
59827 => conv_std_logic_vector(162, 8),
59828 => conv_std_logic_vector(163, 8),
59829 => conv_std_logic_vector(164, 8),
59830 => conv_std_logic_vector(165, 8),
59831 => conv_std_logic_vector(166, 8),
59832 => conv_std_logic_vector(167, 8),
59833 => conv_std_logic_vector(168, 8),
59834 => conv_std_logic_vector(169, 8),
59835 => conv_std_logic_vector(170, 8),
59836 => conv_std_logic_vector(171, 8),
59837 => conv_std_logic_vector(172, 8),
59838 => conv_std_logic_vector(172, 8),
59839 => conv_std_logic_vector(173, 8),
59840 => conv_std_logic_vector(174, 8),
59841 => conv_std_logic_vector(175, 8),
59842 => conv_std_logic_vector(176, 8),
59843 => conv_std_logic_vector(177, 8),
59844 => conv_std_logic_vector(178, 8),
59845 => conv_std_logic_vector(179, 8),
59846 => conv_std_logic_vector(180, 8),
59847 => conv_std_logic_vector(181, 8),
59848 => conv_std_logic_vector(182, 8),
59849 => conv_std_logic_vector(182, 8),
59850 => conv_std_logic_vector(183, 8),
59851 => conv_std_logic_vector(184, 8),
59852 => conv_std_logic_vector(185, 8),
59853 => conv_std_logic_vector(186, 8),
59854 => conv_std_logic_vector(187, 8),
59855 => conv_std_logic_vector(188, 8),
59856 => conv_std_logic_vector(189, 8),
59857 => conv_std_logic_vector(190, 8),
59858 => conv_std_logic_vector(191, 8),
59859 => conv_std_logic_vector(192, 8),
59860 => conv_std_logic_vector(192, 8),
59861 => conv_std_logic_vector(193, 8),
59862 => conv_std_logic_vector(194, 8),
59863 => conv_std_logic_vector(195, 8),
59864 => conv_std_logic_vector(196, 8),
59865 => conv_std_logic_vector(197, 8),
59866 => conv_std_logic_vector(198, 8),
59867 => conv_std_logic_vector(199, 8),
59868 => conv_std_logic_vector(200, 8),
59869 => conv_std_logic_vector(201, 8),
59870 => conv_std_logic_vector(202, 8),
59871 => conv_std_logic_vector(202, 8),
59872 => conv_std_logic_vector(203, 8),
59873 => conv_std_logic_vector(204, 8),
59874 => conv_std_logic_vector(205, 8),
59875 => conv_std_logic_vector(206, 8),
59876 => conv_std_logic_vector(207, 8),
59877 => conv_std_logic_vector(208, 8),
59878 => conv_std_logic_vector(209, 8),
59879 => conv_std_logic_vector(210, 8),
59880 => conv_std_logic_vector(211, 8),
59881 => conv_std_logic_vector(212, 8),
59882 => conv_std_logic_vector(212, 8),
59883 => conv_std_logic_vector(213, 8),
59884 => conv_std_logic_vector(214, 8),
59885 => conv_std_logic_vector(215, 8),
59886 => conv_std_logic_vector(216, 8),
59887 => conv_std_logic_vector(217, 8),
59888 => conv_std_logic_vector(218, 8),
59889 => conv_std_logic_vector(219, 8),
59890 => conv_std_logic_vector(220, 8),
59891 => conv_std_logic_vector(221, 8),
59892 => conv_std_logic_vector(222, 8),
59893 => conv_std_logic_vector(222, 8),
59894 => conv_std_logic_vector(223, 8),
59895 => conv_std_logic_vector(224, 8),
59896 => conv_std_logic_vector(225, 8),
59897 => conv_std_logic_vector(226, 8),
59898 => conv_std_logic_vector(227, 8),
59899 => conv_std_logic_vector(228, 8),
59900 => conv_std_logic_vector(229, 8),
59901 => conv_std_logic_vector(230, 8),
59902 => conv_std_logic_vector(231, 8),
59903 => conv_std_logic_vector(232, 8),
59904 => conv_std_logic_vector(0, 8),
59905 => conv_std_logic_vector(0, 8),
59906 => conv_std_logic_vector(1, 8),
59907 => conv_std_logic_vector(2, 8),
59908 => conv_std_logic_vector(3, 8),
59909 => conv_std_logic_vector(4, 8),
59910 => conv_std_logic_vector(5, 8),
59911 => conv_std_logic_vector(6, 8),
59912 => conv_std_logic_vector(7, 8),
59913 => conv_std_logic_vector(8, 8),
59914 => conv_std_logic_vector(9, 8),
59915 => conv_std_logic_vector(10, 8),
59916 => conv_std_logic_vector(10, 8),
59917 => conv_std_logic_vector(11, 8),
59918 => conv_std_logic_vector(12, 8),
59919 => conv_std_logic_vector(13, 8),
59920 => conv_std_logic_vector(14, 8),
59921 => conv_std_logic_vector(15, 8),
59922 => conv_std_logic_vector(16, 8),
59923 => conv_std_logic_vector(17, 8),
59924 => conv_std_logic_vector(18, 8),
59925 => conv_std_logic_vector(19, 8),
59926 => conv_std_logic_vector(20, 8),
59927 => conv_std_logic_vector(21, 8),
59928 => conv_std_logic_vector(21, 8),
59929 => conv_std_logic_vector(22, 8),
59930 => conv_std_logic_vector(23, 8),
59931 => conv_std_logic_vector(24, 8),
59932 => conv_std_logic_vector(25, 8),
59933 => conv_std_logic_vector(26, 8),
59934 => conv_std_logic_vector(27, 8),
59935 => conv_std_logic_vector(28, 8),
59936 => conv_std_logic_vector(29, 8),
59937 => conv_std_logic_vector(30, 8),
59938 => conv_std_logic_vector(31, 8),
59939 => conv_std_logic_vector(31, 8),
59940 => conv_std_logic_vector(32, 8),
59941 => conv_std_logic_vector(33, 8),
59942 => conv_std_logic_vector(34, 8),
59943 => conv_std_logic_vector(35, 8),
59944 => conv_std_logic_vector(36, 8),
59945 => conv_std_logic_vector(37, 8),
59946 => conv_std_logic_vector(38, 8),
59947 => conv_std_logic_vector(39, 8),
59948 => conv_std_logic_vector(40, 8),
59949 => conv_std_logic_vector(41, 8),
59950 => conv_std_logic_vector(42, 8),
59951 => conv_std_logic_vector(42, 8),
59952 => conv_std_logic_vector(43, 8),
59953 => conv_std_logic_vector(44, 8),
59954 => conv_std_logic_vector(45, 8),
59955 => conv_std_logic_vector(46, 8),
59956 => conv_std_logic_vector(47, 8),
59957 => conv_std_logic_vector(48, 8),
59958 => conv_std_logic_vector(49, 8),
59959 => conv_std_logic_vector(50, 8),
59960 => conv_std_logic_vector(51, 8),
59961 => conv_std_logic_vector(52, 8),
59962 => conv_std_logic_vector(53, 8),
59963 => conv_std_logic_vector(53, 8),
59964 => conv_std_logic_vector(54, 8),
59965 => conv_std_logic_vector(55, 8),
59966 => conv_std_logic_vector(56, 8),
59967 => conv_std_logic_vector(57, 8),
59968 => conv_std_logic_vector(58, 8),
59969 => conv_std_logic_vector(59, 8),
59970 => conv_std_logic_vector(60, 8),
59971 => conv_std_logic_vector(61, 8),
59972 => conv_std_logic_vector(62, 8),
59973 => conv_std_logic_vector(63, 8),
59974 => conv_std_logic_vector(63, 8),
59975 => conv_std_logic_vector(64, 8),
59976 => conv_std_logic_vector(65, 8),
59977 => conv_std_logic_vector(66, 8),
59978 => conv_std_logic_vector(67, 8),
59979 => conv_std_logic_vector(68, 8),
59980 => conv_std_logic_vector(69, 8),
59981 => conv_std_logic_vector(70, 8),
59982 => conv_std_logic_vector(71, 8),
59983 => conv_std_logic_vector(72, 8),
59984 => conv_std_logic_vector(73, 8),
59985 => conv_std_logic_vector(74, 8),
59986 => conv_std_logic_vector(74, 8),
59987 => conv_std_logic_vector(75, 8),
59988 => conv_std_logic_vector(76, 8),
59989 => conv_std_logic_vector(77, 8),
59990 => conv_std_logic_vector(78, 8),
59991 => conv_std_logic_vector(79, 8),
59992 => conv_std_logic_vector(80, 8),
59993 => conv_std_logic_vector(81, 8),
59994 => conv_std_logic_vector(82, 8),
59995 => conv_std_logic_vector(83, 8),
59996 => conv_std_logic_vector(84, 8),
59997 => conv_std_logic_vector(85, 8),
59998 => conv_std_logic_vector(85, 8),
59999 => conv_std_logic_vector(86, 8),
60000 => conv_std_logic_vector(87, 8),
60001 => conv_std_logic_vector(88, 8),
60002 => conv_std_logic_vector(89, 8),
60003 => conv_std_logic_vector(90, 8),
60004 => conv_std_logic_vector(91, 8),
60005 => conv_std_logic_vector(92, 8),
60006 => conv_std_logic_vector(93, 8),
60007 => conv_std_logic_vector(94, 8),
60008 => conv_std_logic_vector(95, 8),
60009 => conv_std_logic_vector(95, 8),
60010 => conv_std_logic_vector(96, 8),
60011 => conv_std_logic_vector(97, 8),
60012 => conv_std_logic_vector(98, 8),
60013 => conv_std_logic_vector(99, 8),
60014 => conv_std_logic_vector(100, 8),
60015 => conv_std_logic_vector(101, 8),
60016 => conv_std_logic_vector(102, 8),
60017 => conv_std_logic_vector(103, 8),
60018 => conv_std_logic_vector(104, 8),
60019 => conv_std_logic_vector(105, 8),
60020 => conv_std_logic_vector(106, 8),
60021 => conv_std_logic_vector(106, 8),
60022 => conv_std_logic_vector(107, 8),
60023 => conv_std_logic_vector(108, 8),
60024 => conv_std_logic_vector(109, 8),
60025 => conv_std_logic_vector(110, 8),
60026 => conv_std_logic_vector(111, 8),
60027 => conv_std_logic_vector(112, 8),
60028 => conv_std_logic_vector(113, 8),
60029 => conv_std_logic_vector(114, 8),
60030 => conv_std_logic_vector(115, 8),
60031 => conv_std_logic_vector(116, 8),
60032 => conv_std_logic_vector(117, 8),
60033 => conv_std_logic_vector(117, 8),
60034 => conv_std_logic_vector(118, 8),
60035 => conv_std_logic_vector(119, 8),
60036 => conv_std_logic_vector(120, 8),
60037 => conv_std_logic_vector(121, 8),
60038 => conv_std_logic_vector(122, 8),
60039 => conv_std_logic_vector(123, 8),
60040 => conv_std_logic_vector(124, 8),
60041 => conv_std_logic_vector(125, 8),
60042 => conv_std_logic_vector(126, 8),
60043 => conv_std_logic_vector(127, 8),
60044 => conv_std_logic_vector(127, 8),
60045 => conv_std_logic_vector(128, 8),
60046 => conv_std_logic_vector(129, 8),
60047 => conv_std_logic_vector(130, 8),
60048 => conv_std_logic_vector(131, 8),
60049 => conv_std_logic_vector(132, 8),
60050 => conv_std_logic_vector(133, 8),
60051 => conv_std_logic_vector(134, 8),
60052 => conv_std_logic_vector(135, 8),
60053 => conv_std_logic_vector(136, 8),
60054 => conv_std_logic_vector(137, 8),
60055 => conv_std_logic_vector(138, 8),
60056 => conv_std_logic_vector(138, 8),
60057 => conv_std_logic_vector(139, 8),
60058 => conv_std_logic_vector(140, 8),
60059 => conv_std_logic_vector(141, 8),
60060 => conv_std_logic_vector(142, 8),
60061 => conv_std_logic_vector(143, 8),
60062 => conv_std_logic_vector(144, 8),
60063 => conv_std_logic_vector(145, 8),
60064 => conv_std_logic_vector(146, 8),
60065 => conv_std_logic_vector(147, 8),
60066 => conv_std_logic_vector(148, 8),
60067 => conv_std_logic_vector(148, 8),
60068 => conv_std_logic_vector(149, 8),
60069 => conv_std_logic_vector(150, 8),
60070 => conv_std_logic_vector(151, 8),
60071 => conv_std_logic_vector(152, 8),
60072 => conv_std_logic_vector(153, 8),
60073 => conv_std_logic_vector(154, 8),
60074 => conv_std_logic_vector(155, 8),
60075 => conv_std_logic_vector(156, 8),
60076 => conv_std_logic_vector(157, 8),
60077 => conv_std_logic_vector(158, 8),
60078 => conv_std_logic_vector(159, 8),
60079 => conv_std_logic_vector(159, 8),
60080 => conv_std_logic_vector(160, 8),
60081 => conv_std_logic_vector(161, 8),
60082 => conv_std_logic_vector(162, 8),
60083 => conv_std_logic_vector(163, 8),
60084 => conv_std_logic_vector(164, 8),
60085 => conv_std_logic_vector(165, 8),
60086 => conv_std_logic_vector(166, 8),
60087 => conv_std_logic_vector(167, 8),
60088 => conv_std_logic_vector(168, 8),
60089 => conv_std_logic_vector(169, 8),
60090 => conv_std_logic_vector(170, 8),
60091 => conv_std_logic_vector(170, 8),
60092 => conv_std_logic_vector(171, 8),
60093 => conv_std_logic_vector(172, 8),
60094 => conv_std_logic_vector(173, 8),
60095 => conv_std_logic_vector(174, 8),
60096 => conv_std_logic_vector(175, 8),
60097 => conv_std_logic_vector(176, 8),
60098 => conv_std_logic_vector(177, 8),
60099 => conv_std_logic_vector(178, 8),
60100 => conv_std_logic_vector(179, 8),
60101 => conv_std_logic_vector(180, 8),
60102 => conv_std_logic_vector(180, 8),
60103 => conv_std_logic_vector(181, 8),
60104 => conv_std_logic_vector(182, 8),
60105 => conv_std_logic_vector(183, 8),
60106 => conv_std_logic_vector(184, 8),
60107 => conv_std_logic_vector(185, 8),
60108 => conv_std_logic_vector(186, 8),
60109 => conv_std_logic_vector(187, 8),
60110 => conv_std_logic_vector(188, 8),
60111 => conv_std_logic_vector(189, 8),
60112 => conv_std_logic_vector(190, 8),
60113 => conv_std_logic_vector(191, 8),
60114 => conv_std_logic_vector(191, 8),
60115 => conv_std_logic_vector(192, 8),
60116 => conv_std_logic_vector(193, 8),
60117 => conv_std_logic_vector(194, 8),
60118 => conv_std_logic_vector(195, 8),
60119 => conv_std_logic_vector(196, 8),
60120 => conv_std_logic_vector(197, 8),
60121 => conv_std_logic_vector(198, 8),
60122 => conv_std_logic_vector(199, 8),
60123 => conv_std_logic_vector(200, 8),
60124 => conv_std_logic_vector(201, 8),
60125 => conv_std_logic_vector(202, 8),
60126 => conv_std_logic_vector(202, 8),
60127 => conv_std_logic_vector(203, 8),
60128 => conv_std_logic_vector(204, 8),
60129 => conv_std_logic_vector(205, 8),
60130 => conv_std_logic_vector(206, 8),
60131 => conv_std_logic_vector(207, 8),
60132 => conv_std_logic_vector(208, 8),
60133 => conv_std_logic_vector(209, 8),
60134 => conv_std_logic_vector(210, 8),
60135 => conv_std_logic_vector(211, 8),
60136 => conv_std_logic_vector(212, 8),
60137 => conv_std_logic_vector(212, 8),
60138 => conv_std_logic_vector(213, 8),
60139 => conv_std_logic_vector(214, 8),
60140 => conv_std_logic_vector(215, 8),
60141 => conv_std_logic_vector(216, 8),
60142 => conv_std_logic_vector(217, 8),
60143 => conv_std_logic_vector(218, 8),
60144 => conv_std_logic_vector(219, 8),
60145 => conv_std_logic_vector(220, 8),
60146 => conv_std_logic_vector(221, 8),
60147 => conv_std_logic_vector(222, 8),
60148 => conv_std_logic_vector(223, 8),
60149 => conv_std_logic_vector(223, 8),
60150 => conv_std_logic_vector(224, 8),
60151 => conv_std_logic_vector(225, 8),
60152 => conv_std_logic_vector(226, 8),
60153 => conv_std_logic_vector(227, 8),
60154 => conv_std_logic_vector(228, 8),
60155 => conv_std_logic_vector(229, 8),
60156 => conv_std_logic_vector(230, 8),
60157 => conv_std_logic_vector(231, 8),
60158 => conv_std_logic_vector(232, 8),
60159 => conv_std_logic_vector(233, 8),
60160 => conv_std_logic_vector(0, 8),
60161 => conv_std_logic_vector(0, 8),
60162 => conv_std_logic_vector(1, 8),
60163 => conv_std_logic_vector(2, 8),
60164 => conv_std_logic_vector(3, 8),
60165 => conv_std_logic_vector(4, 8),
60166 => conv_std_logic_vector(5, 8),
60167 => conv_std_logic_vector(6, 8),
60168 => conv_std_logic_vector(7, 8),
60169 => conv_std_logic_vector(8, 8),
60170 => conv_std_logic_vector(9, 8),
60171 => conv_std_logic_vector(10, 8),
60172 => conv_std_logic_vector(11, 8),
60173 => conv_std_logic_vector(11, 8),
60174 => conv_std_logic_vector(12, 8),
60175 => conv_std_logic_vector(13, 8),
60176 => conv_std_logic_vector(14, 8),
60177 => conv_std_logic_vector(15, 8),
60178 => conv_std_logic_vector(16, 8),
60179 => conv_std_logic_vector(17, 8),
60180 => conv_std_logic_vector(18, 8),
60181 => conv_std_logic_vector(19, 8),
60182 => conv_std_logic_vector(20, 8),
60183 => conv_std_logic_vector(21, 8),
60184 => conv_std_logic_vector(22, 8),
60185 => conv_std_logic_vector(22, 8),
60186 => conv_std_logic_vector(23, 8),
60187 => conv_std_logic_vector(24, 8),
60188 => conv_std_logic_vector(25, 8),
60189 => conv_std_logic_vector(26, 8),
60190 => conv_std_logic_vector(27, 8),
60191 => conv_std_logic_vector(28, 8),
60192 => conv_std_logic_vector(29, 8),
60193 => conv_std_logic_vector(30, 8),
60194 => conv_std_logic_vector(31, 8),
60195 => conv_std_logic_vector(32, 8),
60196 => conv_std_logic_vector(33, 8),
60197 => conv_std_logic_vector(33, 8),
60198 => conv_std_logic_vector(34, 8),
60199 => conv_std_logic_vector(35, 8),
60200 => conv_std_logic_vector(36, 8),
60201 => conv_std_logic_vector(37, 8),
60202 => conv_std_logic_vector(38, 8),
60203 => conv_std_logic_vector(39, 8),
60204 => conv_std_logic_vector(40, 8),
60205 => conv_std_logic_vector(41, 8),
60206 => conv_std_logic_vector(42, 8),
60207 => conv_std_logic_vector(43, 8),
60208 => conv_std_logic_vector(44, 8),
60209 => conv_std_logic_vector(44, 8),
60210 => conv_std_logic_vector(45, 8),
60211 => conv_std_logic_vector(46, 8),
60212 => conv_std_logic_vector(47, 8),
60213 => conv_std_logic_vector(48, 8),
60214 => conv_std_logic_vector(49, 8),
60215 => conv_std_logic_vector(50, 8),
60216 => conv_std_logic_vector(51, 8),
60217 => conv_std_logic_vector(52, 8),
60218 => conv_std_logic_vector(53, 8),
60219 => conv_std_logic_vector(54, 8),
60220 => conv_std_logic_vector(55, 8),
60221 => conv_std_logic_vector(55, 8),
60222 => conv_std_logic_vector(56, 8),
60223 => conv_std_logic_vector(57, 8),
60224 => conv_std_logic_vector(58, 8),
60225 => conv_std_logic_vector(59, 8),
60226 => conv_std_logic_vector(60, 8),
60227 => conv_std_logic_vector(61, 8),
60228 => conv_std_logic_vector(62, 8),
60229 => conv_std_logic_vector(63, 8),
60230 => conv_std_logic_vector(64, 8),
60231 => conv_std_logic_vector(65, 8),
60232 => conv_std_logic_vector(66, 8),
60233 => conv_std_logic_vector(67, 8),
60234 => conv_std_logic_vector(67, 8),
60235 => conv_std_logic_vector(68, 8),
60236 => conv_std_logic_vector(69, 8),
60237 => conv_std_logic_vector(70, 8),
60238 => conv_std_logic_vector(71, 8),
60239 => conv_std_logic_vector(72, 8),
60240 => conv_std_logic_vector(73, 8),
60241 => conv_std_logic_vector(74, 8),
60242 => conv_std_logic_vector(75, 8),
60243 => conv_std_logic_vector(76, 8),
60244 => conv_std_logic_vector(77, 8),
60245 => conv_std_logic_vector(78, 8),
60246 => conv_std_logic_vector(78, 8),
60247 => conv_std_logic_vector(79, 8),
60248 => conv_std_logic_vector(80, 8),
60249 => conv_std_logic_vector(81, 8),
60250 => conv_std_logic_vector(82, 8),
60251 => conv_std_logic_vector(83, 8),
60252 => conv_std_logic_vector(84, 8),
60253 => conv_std_logic_vector(85, 8),
60254 => conv_std_logic_vector(86, 8),
60255 => conv_std_logic_vector(87, 8),
60256 => conv_std_logic_vector(88, 8),
60257 => conv_std_logic_vector(89, 8),
60258 => conv_std_logic_vector(89, 8),
60259 => conv_std_logic_vector(90, 8),
60260 => conv_std_logic_vector(91, 8),
60261 => conv_std_logic_vector(92, 8),
60262 => conv_std_logic_vector(93, 8),
60263 => conv_std_logic_vector(94, 8),
60264 => conv_std_logic_vector(95, 8),
60265 => conv_std_logic_vector(96, 8),
60266 => conv_std_logic_vector(97, 8),
60267 => conv_std_logic_vector(98, 8),
60268 => conv_std_logic_vector(99, 8),
60269 => conv_std_logic_vector(100, 8),
60270 => conv_std_logic_vector(100, 8),
60271 => conv_std_logic_vector(101, 8),
60272 => conv_std_logic_vector(102, 8),
60273 => conv_std_logic_vector(103, 8),
60274 => conv_std_logic_vector(104, 8),
60275 => conv_std_logic_vector(105, 8),
60276 => conv_std_logic_vector(106, 8),
60277 => conv_std_logic_vector(107, 8),
60278 => conv_std_logic_vector(108, 8),
60279 => conv_std_logic_vector(109, 8),
60280 => conv_std_logic_vector(110, 8),
60281 => conv_std_logic_vector(111, 8),
60282 => conv_std_logic_vector(111, 8),
60283 => conv_std_logic_vector(112, 8),
60284 => conv_std_logic_vector(113, 8),
60285 => conv_std_logic_vector(114, 8),
60286 => conv_std_logic_vector(115, 8),
60287 => conv_std_logic_vector(116, 8),
60288 => conv_std_logic_vector(117, 8),
60289 => conv_std_logic_vector(118, 8),
60290 => conv_std_logic_vector(119, 8),
60291 => conv_std_logic_vector(120, 8),
60292 => conv_std_logic_vector(121, 8),
60293 => conv_std_logic_vector(122, 8),
60294 => conv_std_logic_vector(123, 8),
60295 => conv_std_logic_vector(123, 8),
60296 => conv_std_logic_vector(124, 8),
60297 => conv_std_logic_vector(125, 8),
60298 => conv_std_logic_vector(126, 8),
60299 => conv_std_logic_vector(127, 8),
60300 => conv_std_logic_vector(128, 8),
60301 => conv_std_logic_vector(129, 8),
60302 => conv_std_logic_vector(130, 8),
60303 => conv_std_logic_vector(131, 8),
60304 => conv_std_logic_vector(132, 8),
60305 => conv_std_logic_vector(133, 8),
60306 => conv_std_logic_vector(134, 8),
60307 => conv_std_logic_vector(134, 8),
60308 => conv_std_logic_vector(135, 8),
60309 => conv_std_logic_vector(136, 8),
60310 => conv_std_logic_vector(137, 8),
60311 => conv_std_logic_vector(138, 8),
60312 => conv_std_logic_vector(139, 8),
60313 => conv_std_logic_vector(140, 8),
60314 => conv_std_logic_vector(141, 8),
60315 => conv_std_logic_vector(142, 8),
60316 => conv_std_logic_vector(143, 8),
60317 => conv_std_logic_vector(144, 8),
60318 => conv_std_logic_vector(145, 8),
60319 => conv_std_logic_vector(145, 8),
60320 => conv_std_logic_vector(146, 8),
60321 => conv_std_logic_vector(147, 8),
60322 => conv_std_logic_vector(148, 8),
60323 => conv_std_logic_vector(149, 8),
60324 => conv_std_logic_vector(150, 8),
60325 => conv_std_logic_vector(151, 8),
60326 => conv_std_logic_vector(152, 8),
60327 => conv_std_logic_vector(153, 8),
60328 => conv_std_logic_vector(154, 8),
60329 => conv_std_logic_vector(155, 8),
60330 => conv_std_logic_vector(156, 8),
60331 => conv_std_logic_vector(156, 8),
60332 => conv_std_logic_vector(157, 8),
60333 => conv_std_logic_vector(158, 8),
60334 => conv_std_logic_vector(159, 8),
60335 => conv_std_logic_vector(160, 8),
60336 => conv_std_logic_vector(161, 8),
60337 => conv_std_logic_vector(162, 8),
60338 => conv_std_logic_vector(163, 8),
60339 => conv_std_logic_vector(164, 8),
60340 => conv_std_logic_vector(165, 8),
60341 => conv_std_logic_vector(166, 8),
60342 => conv_std_logic_vector(167, 8),
60343 => conv_std_logic_vector(167, 8),
60344 => conv_std_logic_vector(168, 8),
60345 => conv_std_logic_vector(169, 8),
60346 => conv_std_logic_vector(170, 8),
60347 => conv_std_logic_vector(171, 8),
60348 => conv_std_logic_vector(172, 8),
60349 => conv_std_logic_vector(173, 8),
60350 => conv_std_logic_vector(174, 8),
60351 => conv_std_logic_vector(175, 8),
60352 => conv_std_logic_vector(176, 8),
60353 => conv_std_logic_vector(177, 8),
60354 => conv_std_logic_vector(178, 8),
60355 => conv_std_logic_vector(179, 8),
60356 => conv_std_logic_vector(179, 8),
60357 => conv_std_logic_vector(180, 8),
60358 => conv_std_logic_vector(181, 8),
60359 => conv_std_logic_vector(182, 8),
60360 => conv_std_logic_vector(183, 8),
60361 => conv_std_logic_vector(184, 8),
60362 => conv_std_logic_vector(185, 8),
60363 => conv_std_logic_vector(186, 8),
60364 => conv_std_logic_vector(187, 8),
60365 => conv_std_logic_vector(188, 8),
60366 => conv_std_logic_vector(189, 8),
60367 => conv_std_logic_vector(190, 8),
60368 => conv_std_logic_vector(190, 8),
60369 => conv_std_logic_vector(191, 8),
60370 => conv_std_logic_vector(192, 8),
60371 => conv_std_logic_vector(193, 8),
60372 => conv_std_logic_vector(194, 8),
60373 => conv_std_logic_vector(195, 8),
60374 => conv_std_logic_vector(196, 8),
60375 => conv_std_logic_vector(197, 8),
60376 => conv_std_logic_vector(198, 8),
60377 => conv_std_logic_vector(199, 8),
60378 => conv_std_logic_vector(200, 8),
60379 => conv_std_logic_vector(201, 8),
60380 => conv_std_logic_vector(201, 8),
60381 => conv_std_logic_vector(202, 8),
60382 => conv_std_logic_vector(203, 8),
60383 => conv_std_logic_vector(204, 8),
60384 => conv_std_logic_vector(205, 8),
60385 => conv_std_logic_vector(206, 8),
60386 => conv_std_logic_vector(207, 8),
60387 => conv_std_logic_vector(208, 8),
60388 => conv_std_logic_vector(209, 8),
60389 => conv_std_logic_vector(210, 8),
60390 => conv_std_logic_vector(211, 8),
60391 => conv_std_logic_vector(212, 8),
60392 => conv_std_logic_vector(212, 8),
60393 => conv_std_logic_vector(213, 8),
60394 => conv_std_logic_vector(214, 8),
60395 => conv_std_logic_vector(215, 8),
60396 => conv_std_logic_vector(216, 8),
60397 => conv_std_logic_vector(217, 8),
60398 => conv_std_logic_vector(218, 8),
60399 => conv_std_logic_vector(219, 8),
60400 => conv_std_logic_vector(220, 8),
60401 => conv_std_logic_vector(221, 8),
60402 => conv_std_logic_vector(222, 8),
60403 => conv_std_logic_vector(223, 8),
60404 => conv_std_logic_vector(223, 8),
60405 => conv_std_logic_vector(224, 8),
60406 => conv_std_logic_vector(225, 8),
60407 => conv_std_logic_vector(226, 8),
60408 => conv_std_logic_vector(227, 8),
60409 => conv_std_logic_vector(228, 8),
60410 => conv_std_logic_vector(229, 8),
60411 => conv_std_logic_vector(230, 8),
60412 => conv_std_logic_vector(231, 8),
60413 => conv_std_logic_vector(232, 8),
60414 => conv_std_logic_vector(233, 8),
60415 => conv_std_logic_vector(234, 8),
60416 => conv_std_logic_vector(0, 8),
60417 => conv_std_logic_vector(0, 8),
60418 => conv_std_logic_vector(1, 8),
60419 => conv_std_logic_vector(2, 8),
60420 => conv_std_logic_vector(3, 8),
60421 => conv_std_logic_vector(4, 8),
60422 => conv_std_logic_vector(5, 8),
60423 => conv_std_logic_vector(6, 8),
60424 => conv_std_logic_vector(7, 8),
60425 => conv_std_logic_vector(8, 8),
60426 => conv_std_logic_vector(9, 8),
60427 => conv_std_logic_vector(10, 8),
60428 => conv_std_logic_vector(11, 8),
60429 => conv_std_logic_vector(11, 8),
60430 => conv_std_logic_vector(12, 8),
60431 => conv_std_logic_vector(13, 8),
60432 => conv_std_logic_vector(14, 8),
60433 => conv_std_logic_vector(15, 8),
60434 => conv_std_logic_vector(16, 8),
60435 => conv_std_logic_vector(17, 8),
60436 => conv_std_logic_vector(18, 8),
60437 => conv_std_logic_vector(19, 8),
60438 => conv_std_logic_vector(20, 8),
60439 => conv_std_logic_vector(21, 8),
60440 => conv_std_logic_vector(22, 8),
60441 => conv_std_logic_vector(23, 8),
60442 => conv_std_logic_vector(23, 8),
60443 => conv_std_logic_vector(24, 8),
60444 => conv_std_logic_vector(25, 8),
60445 => conv_std_logic_vector(26, 8),
60446 => conv_std_logic_vector(27, 8),
60447 => conv_std_logic_vector(28, 8),
60448 => conv_std_logic_vector(29, 8),
60449 => conv_std_logic_vector(30, 8),
60450 => conv_std_logic_vector(31, 8),
60451 => conv_std_logic_vector(32, 8),
60452 => conv_std_logic_vector(33, 8),
60453 => conv_std_logic_vector(34, 8),
60454 => conv_std_logic_vector(35, 8),
60455 => conv_std_logic_vector(35, 8),
60456 => conv_std_logic_vector(36, 8),
60457 => conv_std_logic_vector(37, 8),
60458 => conv_std_logic_vector(38, 8),
60459 => conv_std_logic_vector(39, 8),
60460 => conv_std_logic_vector(40, 8),
60461 => conv_std_logic_vector(41, 8),
60462 => conv_std_logic_vector(42, 8),
60463 => conv_std_logic_vector(43, 8),
60464 => conv_std_logic_vector(44, 8),
60465 => conv_std_logic_vector(45, 8),
60466 => conv_std_logic_vector(46, 8),
60467 => conv_std_logic_vector(47, 8),
60468 => conv_std_logic_vector(47, 8),
60469 => conv_std_logic_vector(48, 8),
60470 => conv_std_logic_vector(49, 8),
60471 => conv_std_logic_vector(50, 8),
60472 => conv_std_logic_vector(51, 8),
60473 => conv_std_logic_vector(52, 8),
60474 => conv_std_logic_vector(53, 8),
60475 => conv_std_logic_vector(54, 8),
60476 => conv_std_logic_vector(55, 8),
60477 => conv_std_logic_vector(56, 8),
60478 => conv_std_logic_vector(57, 8),
60479 => conv_std_logic_vector(58, 8),
60480 => conv_std_logic_vector(59, 8),
60481 => conv_std_logic_vector(59, 8),
60482 => conv_std_logic_vector(60, 8),
60483 => conv_std_logic_vector(61, 8),
60484 => conv_std_logic_vector(62, 8),
60485 => conv_std_logic_vector(63, 8),
60486 => conv_std_logic_vector(64, 8),
60487 => conv_std_logic_vector(65, 8),
60488 => conv_std_logic_vector(66, 8),
60489 => conv_std_logic_vector(67, 8),
60490 => conv_std_logic_vector(68, 8),
60491 => conv_std_logic_vector(69, 8),
60492 => conv_std_logic_vector(70, 8),
60493 => conv_std_logic_vector(70, 8),
60494 => conv_std_logic_vector(71, 8),
60495 => conv_std_logic_vector(72, 8),
60496 => conv_std_logic_vector(73, 8),
60497 => conv_std_logic_vector(74, 8),
60498 => conv_std_logic_vector(75, 8),
60499 => conv_std_logic_vector(76, 8),
60500 => conv_std_logic_vector(77, 8),
60501 => conv_std_logic_vector(78, 8),
60502 => conv_std_logic_vector(79, 8),
60503 => conv_std_logic_vector(80, 8),
60504 => conv_std_logic_vector(81, 8),
60505 => conv_std_logic_vector(82, 8),
60506 => conv_std_logic_vector(82, 8),
60507 => conv_std_logic_vector(83, 8),
60508 => conv_std_logic_vector(84, 8),
60509 => conv_std_logic_vector(85, 8),
60510 => conv_std_logic_vector(86, 8),
60511 => conv_std_logic_vector(87, 8),
60512 => conv_std_logic_vector(88, 8),
60513 => conv_std_logic_vector(89, 8),
60514 => conv_std_logic_vector(90, 8),
60515 => conv_std_logic_vector(91, 8),
60516 => conv_std_logic_vector(92, 8),
60517 => conv_std_logic_vector(93, 8),
60518 => conv_std_logic_vector(94, 8),
60519 => conv_std_logic_vector(94, 8),
60520 => conv_std_logic_vector(95, 8),
60521 => conv_std_logic_vector(96, 8),
60522 => conv_std_logic_vector(97, 8),
60523 => conv_std_logic_vector(98, 8),
60524 => conv_std_logic_vector(99, 8),
60525 => conv_std_logic_vector(100, 8),
60526 => conv_std_logic_vector(101, 8),
60527 => conv_std_logic_vector(102, 8),
60528 => conv_std_logic_vector(103, 8),
60529 => conv_std_logic_vector(104, 8),
60530 => conv_std_logic_vector(105, 8),
60531 => conv_std_logic_vector(106, 8),
60532 => conv_std_logic_vector(106, 8),
60533 => conv_std_logic_vector(107, 8),
60534 => conv_std_logic_vector(108, 8),
60535 => conv_std_logic_vector(109, 8),
60536 => conv_std_logic_vector(110, 8),
60537 => conv_std_logic_vector(111, 8),
60538 => conv_std_logic_vector(112, 8),
60539 => conv_std_logic_vector(113, 8),
60540 => conv_std_logic_vector(114, 8),
60541 => conv_std_logic_vector(115, 8),
60542 => conv_std_logic_vector(116, 8),
60543 => conv_std_logic_vector(117, 8),
60544 => conv_std_logic_vector(118, 8),
60545 => conv_std_logic_vector(118, 8),
60546 => conv_std_logic_vector(119, 8),
60547 => conv_std_logic_vector(120, 8),
60548 => conv_std_logic_vector(121, 8),
60549 => conv_std_logic_vector(122, 8),
60550 => conv_std_logic_vector(123, 8),
60551 => conv_std_logic_vector(124, 8),
60552 => conv_std_logic_vector(125, 8),
60553 => conv_std_logic_vector(126, 8),
60554 => conv_std_logic_vector(127, 8),
60555 => conv_std_logic_vector(128, 8),
60556 => conv_std_logic_vector(129, 8),
60557 => conv_std_logic_vector(129, 8),
60558 => conv_std_logic_vector(130, 8),
60559 => conv_std_logic_vector(131, 8),
60560 => conv_std_logic_vector(132, 8),
60561 => conv_std_logic_vector(133, 8),
60562 => conv_std_logic_vector(134, 8),
60563 => conv_std_logic_vector(135, 8),
60564 => conv_std_logic_vector(136, 8),
60565 => conv_std_logic_vector(137, 8),
60566 => conv_std_logic_vector(138, 8),
60567 => conv_std_logic_vector(139, 8),
60568 => conv_std_logic_vector(140, 8),
60569 => conv_std_logic_vector(141, 8),
60570 => conv_std_logic_vector(141, 8),
60571 => conv_std_logic_vector(142, 8),
60572 => conv_std_logic_vector(143, 8),
60573 => conv_std_logic_vector(144, 8),
60574 => conv_std_logic_vector(145, 8),
60575 => conv_std_logic_vector(146, 8),
60576 => conv_std_logic_vector(147, 8),
60577 => conv_std_logic_vector(148, 8),
60578 => conv_std_logic_vector(149, 8),
60579 => conv_std_logic_vector(150, 8),
60580 => conv_std_logic_vector(151, 8),
60581 => conv_std_logic_vector(152, 8),
60582 => conv_std_logic_vector(153, 8),
60583 => conv_std_logic_vector(153, 8),
60584 => conv_std_logic_vector(154, 8),
60585 => conv_std_logic_vector(155, 8),
60586 => conv_std_logic_vector(156, 8),
60587 => conv_std_logic_vector(157, 8),
60588 => conv_std_logic_vector(158, 8),
60589 => conv_std_logic_vector(159, 8),
60590 => conv_std_logic_vector(160, 8),
60591 => conv_std_logic_vector(161, 8),
60592 => conv_std_logic_vector(162, 8),
60593 => conv_std_logic_vector(163, 8),
60594 => conv_std_logic_vector(164, 8),
60595 => conv_std_logic_vector(165, 8),
60596 => conv_std_logic_vector(165, 8),
60597 => conv_std_logic_vector(166, 8),
60598 => conv_std_logic_vector(167, 8),
60599 => conv_std_logic_vector(168, 8),
60600 => conv_std_logic_vector(169, 8),
60601 => conv_std_logic_vector(170, 8),
60602 => conv_std_logic_vector(171, 8),
60603 => conv_std_logic_vector(172, 8),
60604 => conv_std_logic_vector(173, 8),
60605 => conv_std_logic_vector(174, 8),
60606 => conv_std_logic_vector(175, 8),
60607 => conv_std_logic_vector(176, 8),
60608 => conv_std_logic_vector(177, 8),
60609 => conv_std_logic_vector(177, 8),
60610 => conv_std_logic_vector(178, 8),
60611 => conv_std_logic_vector(179, 8),
60612 => conv_std_logic_vector(180, 8),
60613 => conv_std_logic_vector(181, 8),
60614 => conv_std_logic_vector(182, 8),
60615 => conv_std_logic_vector(183, 8),
60616 => conv_std_logic_vector(184, 8),
60617 => conv_std_logic_vector(185, 8),
60618 => conv_std_logic_vector(186, 8),
60619 => conv_std_logic_vector(187, 8),
60620 => conv_std_logic_vector(188, 8),
60621 => conv_std_logic_vector(188, 8),
60622 => conv_std_logic_vector(189, 8),
60623 => conv_std_logic_vector(190, 8),
60624 => conv_std_logic_vector(191, 8),
60625 => conv_std_logic_vector(192, 8),
60626 => conv_std_logic_vector(193, 8),
60627 => conv_std_logic_vector(194, 8),
60628 => conv_std_logic_vector(195, 8),
60629 => conv_std_logic_vector(196, 8),
60630 => conv_std_logic_vector(197, 8),
60631 => conv_std_logic_vector(198, 8),
60632 => conv_std_logic_vector(199, 8),
60633 => conv_std_logic_vector(200, 8),
60634 => conv_std_logic_vector(200, 8),
60635 => conv_std_logic_vector(201, 8),
60636 => conv_std_logic_vector(202, 8),
60637 => conv_std_logic_vector(203, 8),
60638 => conv_std_logic_vector(204, 8),
60639 => conv_std_logic_vector(205, 8),
60640 => conv_std_logic_vector(206, 8),
60641 => conv_std_logic_vector(207, 8),
60642 => conv_std_logic_vector(208, 8),
60643 => conv_std_logic_vector(209, 8),
60644 => conv_std_logic_vector(210, 8),
60645 => conv_std_logic_vector(211, 8),
60646 => conv_std_logic_vector(212, 8),
60647 => conv_std_logic_vector(212, 8),
60648 => conv_std_logic_vector(213, 8),
60649 => conv_std_logic_vector(214, 8),
60650 => conv_std_logic_vector(215, 8),
60651 => conv_std_logic_vector(216, 8),
60652 => conv_std_logic_vector(217, 8),
60653 => conv_std_logic_vector(218, 8),
60654 => conv_std_logic_vector(219, 8),
60655 => conv_std_logic_vector(220, 8),
60656 => conv_std_logic_vector(221, 8),
60657 => conv_std_logic_vector(222, 8),
60658 => conv_std_logic_vector(223, 8),
60659 => conv_std_logic_vector(224, 8),
60660 => conv_std_logic_vector(224, 8),
60661 => conv_std_logic_vector(225, 8),
60662 => conv_std_logic_vector(226, 8),
60663 => conv_std_logic_vector(227, 8),
60664 => conv_std_logic_vector(228, 8),
60665 => conv_std_logic_vector(229, 8),
60666 => conv_std_logic_vector(230, 8),
60667 => conv_std_logic_vector(231, 8),
60668 => conv_std_logic_vector(232, 8),
60669 => conv_std_logic_vector(233, 8),
60670 => conv_std_logic_vector(234, 8),
60671 => conv_std_logic_vector(235, 8),
60672 => conv_std_logic_vector(0, 8),
60673 => conv_std_logic_vector(0, 8),
60674 => conv_std_logic_vector(1, 8),
60675 => conv_std_logic_vector(2, 8),
60676 => conv_std_logic_vector(3, 8),
60677 => conv_std_logic_vector(4, 8),
60678 => conv_std_logic_vector(5, 8),
60679 => conv_std_logic_vector(6, 8),
60680 => conv_std_logic_vector(7, 8),
60681 => conv_std_logic_vector(8, 8),
60682 => conv_std_logic_vector(9, 8),
60683 => conv_std_logic_vector(10, 8),
60684 => conv_std_logic_vector(11, 8),
60685 => conv_std_logic_vector(12, 8),
60686 => conv_std_logic_vector(12, 8),
60687 => conv_std_logic_vector(13, 8),
60688 => conv_std_logic_vector(14, 8),
60689 => conv_std_logic_vector(15, 8),
60690 => conv_std_logic_vector(16, 8),
60691 => conv_std_logic_vector(17, 8),
60692 => conv_std_logic_vector(18, 8),
60693 => conv_std_logic_vector(19, 8),
60694 => conv_std_logic_vector(20, 8),
60695 => conv_std_logic_vector(21, 8),
60696 => conv_std_logic_vector(22, 8),
60697 => conv_std_logic_vector(23, 8),
60698 => conv_std_logic_vector(24, 8),
60699 => conv_std_logic_vector(24, 8),
60700 => conv_std_logic_vector(25, 8),
60701 => conv_std_logic_vector(26, 8),
60702 => conv_std_logic_vector(27, 8),
60703 => conv_std_logic_vector(28, 8),
60704 => conv_std_logic_vector(29, 8),
60705 => conv_std_logic_vector(30, 8),
60706 => conv_std_logic_vector(31, 8),
60707 => conv_std_logic_vector(32, 8),
60708 => conv_std_logic_vector(33, 8),
60709 => conv_std_logic_vector(34, 8),
60710 => conv_std_logic_vector(35, 8),
60711 => conv_std_logic_vector(36, 8),
60712 => conv_std_logic_vector(37, 8),
60713 => conv_std_logic_vector(37, 8),
60714 => conv_std_logic_vector(38, 8),
60715 => conv_std_logic_vector(39, 8),
60716 => conv_std_logic_vector(40, 8),
60717 => conv_std_logic_vector(41, 8),
60718 => conv_std_logic_vector(42, 8),
60719 => conv_std_logic_vector(43, 8),
60720 => conv_std_logic_vector(44, 8),
60721 => conv_std_logic_vector(45, 8),
60722 => conv_std_logic_vector(46, 8),
60723 => conv_std_logic_vector(47, 8),
60724 => conv_std_logic_vector(48, 8),
60725 => conv_std_logic_vector(49, 8),
60726 => conv_std_logic_vector(49, 8),
60727 => conv_std_logic_vector(50, 8),
60728 => conv_std_logic_vector(51, 8),
60729 => conv_std_logic_vector(52, 8),
60730 => conv_std_logic_vector(53, 8),
60731 => conv_std_logic_vector(54, 8),
60732 => conv_std_logic_vector(55, 8),
60733 => conv_std_logic_vector(56, 8),
60734 => conv_std_logic_vector(57, 8),
60735 => conv_std_logic_vector(58, 8),
60736 => conv_std_logic_vector(59, 8),
60737 => conv_std_logic_vector(60, 8),
60738 => conv_std_logic_vector(61, 8),
60739 => conv_std_logic_vector(62, 8),
60740 => conv_std_logic_vector(62, 8),
60741 => conv_std_logic_vector(63, 8),
60742 => conv_std_logic_vector(64, 8),
60743 => conv_std_logic_vector(65, 8),
60744 => conv_std_logic_vector(66, 8),
60745 => conv_std_logic_vector(67, 8),
60746 => conv_std_logic_vector(68, 8),
60747 => conv_std_logic_vector(69, 8),
60748 => conv_std_logic_vector(70, 8),
60749 => conv_std_logic_vector(71, 8),
60750 => conv_std_logic_vector(72, 8),
60751 => conv_std_logic_vector(73, 8),
60752 => conv_std_logic_vector(74, 8),
60753 => conv_std_logic_vector(74, 8),
60754 => conv_std_logic_vector(75, 8),
60755 => conv_std_logic_vector(76, 8),
60756 => conv_std_logic_vector(77, 8),
60757 => conv_std_logic_vector(78, 8),
60758 => conv_std_logic_vector(79, 8),
60759 => conv_std_logic_vector(80, 8),
60760 => conv_std_logic_vector(81, 8),
60761 => conv_std_logic_vector(82, 8),
60762 => conv_std_logic_vector(83, 8),
60763 => conv_std_logic_vector(84, 8),
60764 => conv_std_logic_vector(85, 8),
60765 => conv_std_logic_vector(86, 8),
60766 => conv_std_logic_vector(87, 8),
60767 => conv_std_logic_vector(87, 8),
60768 => conv_std_logic_vector(88, 8),
60769 => conv_std_logic_vector(89, 8),
60770 => conv_std_logic_vector(90, 8),
60771 => conv_std_logic_vector(91, 8),
60772 => conv_std_logic_vector(92, 8),
60773 => conv_std_logic_vector(93, 8),
60774 => conv_std_logic_vector(94, 8),
60775 => conv_std_logic_vector(95, 8),
60776 => conv_std_logic_vector(96, 8),
60777 => conv_std_logic_vector(97, 8),
60778 => conv_std_logic_vector(98, 8),
60779 => conv_std_logic_vector(99, 8),
60780 => conv_std_logic_vector(99, 8),
60781 => conv_std_logic_vector(100, 8),
60782 => conv_std_logic_vector(101, 8),
60783 => conv_std_logic_vector(102, 8),
60784 => conv_std_logic_vector(103, 8),
60785 => conv_std_logic_vector(104, 8),
60786 => conv_std_logic_vector(105, 8),
60787 => conv_std_logic_vector(106, 8),
60788 => conv_std_logic_vector(107, 8),
60789 => conv_std_logic_vector(108, 8),
60790 => conv_std_logic_vector(109, 8),
60791 => conv_std_logic_vector(110, 8),
60792 => conv_std_logic_vector(111, 8),
60793 => conv_std_logic_vector(112, 8),
60794 => conv_std_logic_vector(112, 8),
60795 => conv_std_logic_vector(113, 8),
60796 => conv_std_logic_vector(114, 8),
60797 => conv_std_logic_vector(115, 8),
60798 => conv_std_logic_vector(116, 8),
60799 => conv_std_logic_vector(117, 8),
60800 => conv_std_logic_vector(118, 8),
60801 => conv_std_logic_vector(119, 8),
60802 => conv_std_logic_vector(120, 8),
60803 => conv_std_logic_vector(121, 8),
60804 => conv_std_logic_vector(122, 8),
60805 => conv_std_logic_vector(123, 8),
60806 => conv_std_logic_vector(124, 8),
60807 => conv_std_logic_vector(124, 8),
60808 => conv_std_logic_vector(125, 8),
60809 => conv_std_logic_vector(126, 8),
60810 => conv_std_logic_vector(127, 8),
60811 => conv_std_logic_vector(128, 8),
60812 => conv_std_logic_vector(129, 8),
60813 => conv_std_logic_vector(130, 8),
60814 => conv_std_logic_vector(131, 8),
60815 => conv_std_logic_vector(132, 8),
60816 => conv_std_logic_vector(133, 8),
60817 => conv_std_logic_vector(134, 8),
60818 => conv_std_logic_vector(135, 8),
60819 => conv_std_logic_vector(136, 8),
60820 => conv_std_logic_vector(137, 8),
60821 => conv_std_logic_vector(137, 8),
60822 => conv_std_logic_vector(138, 8),
60823 => conv_std_logic_vector(139, 8),
60824 => conv_std_logic_vector(140, 8),
60825 => conv_std_logic_vector(141, 8),
60826 => conv_std_logic_vector(142, 8),
60827 => conv_std_logic_vector(143, 8),
60828 => conv_std_logic_vector(144, 8),
60829 => conv_std_logic_vector(145, 8),
60830 => conv_std_logic_vector(146, 8),
60831 => conv_std_logic_vector(147, 8),
60832 => conv_std_logic_vector(148, 8),
60833 => conv_std_logic_vector(149, 8),
60834 => conv_std_logic_vector(149, 8),
60835 => conv_std_logic_vector(150, 8),
60836 => conv_std_logic_vector(151, 8),
60837 => conv_std_logic_vector(152, 8),
60838 => conv_std_logic_vector(153, 8),
60839 => conv_std_logic_vector(154, 8),
60840 => conv_std_logic_vector(155, 8),
60841 => conv_std_logic_vector(156, 8),
60842 => conv_std_logic_vector(157, 8),
60843 => conv_std_logic_vector(158, 8),
60844 => conv_std_logic_vector(159, 8),
60845 => conv_std_logic_vector(160, 8),
60846 => conv_std_logic_vector(161, 8),
60847 => conv_std_logic_vector(162, 8),
60848 => conv_std_logic_vector(162, 8),
60849 => conv_std_logic_vector(163, 8),
60850 => conv_std_logic_vector(164, 8),
60851 => conv_std_logic_vector(165, 8),
60852 => conv_std_logic_vector(166, 8),
60853 => conv_std_logic_vector(167, 8),
60854 => conv_std_logic_vector(168, 8),
60855 => conv_std_logic_vector(169, 8),
60856 => conv_std_logic_vector(170, 8),
60857 => conv_std_logic_vector(171, 8),
60858 => conv_std_logic_vector(172, 8),
60859 => conv_std_logic_vector(173, 8),
60860 => conv_std_logic_vector(174, 8),
60861 => conv_std_logic_vector(174, 8),
60862 => conv_std_logic_vector(175, 8),
60863 => conv_std_logic_vector(176, 8),
60864 => conv_std_logic_vector(177, 8),
60865 => conv_std_logic_vector(178, 8),
60866 => conv_std_logic_vector(179, 8),
60867 => conv_std_logic_vector(180, 8),
60868 => conv_std_logic_vector(181, 8),
60869 => conv_std_logic_vector(182, 8),
60870 => conv_std_logic_vector(183, 8),
60871 => conv_std_logic_vector(184, 8),
60872 => conv_std_logic_vector(185, 8),
60873 => conv_std_logic_vector(186, 8),
60874 => conv_std_logic_vector(187, 8),
60875 => conv_std_logic_vector(187, 8),
60876 => conv_std_logic_vector(188, 8),
60877 => conv_std_logic_vector(189, 8),
60878 => conv_std_logic_vector(190, 8),
60879 => conv_std_logic_vector(191, 8),
60880 => conv_std_logic_vector(192, 8),
60881 => conv_std_logic_vector(193, 8),
60882 => conv_std_logic_vector(194, 8),
60883 => conv_std_logic_vector(195, 8),
60884 => conv_std_logic_vector(196, 8),
60885 => conv_std_logic_vector(197, 8),
60886 => conv_std_logic_vector(198, 8),
60887 => conv_std_logic_vector(199, 8),
60888 => conv_std_logic_vector(199, 8),
60889 => conv_std_logic_vector(200, 8),
60890 => conv_std_logic_vector(201, 8),
60891 => conv_std_logic_vector(202, 8),
60892 => conv_std_logic_vector(203, 8),
60893 => conv_std_logic_vector(204, 8),
60894 => conv_std_logic_vector(205, 8),
60895 => conv_std_logic_vector(206, 8),
60896 => conv_std_logic_vector(207, 8),
60897 => conv_std_logic_vector(208, 8),
60898 => conv_std_logic_vector(209, 8),
60899 => conv_std_logic_vector(210, 8),
60900 => conv_std_logic_vector(211, 8),
60901 => conv_std_logic_vector(212, 8),
60902 => conv_std_logic_vector(212, 8),
60903 => conv_std_logic_vector(213, 8),
60904 => conv_std_logic_vector(214, 8),
60905 => conv_std_logic_vector(215, 8),
60906 => conv_std_logic_vector(216, 8),
60907 => conv_std_logic_vector(217, 8),
60908 => conv_std_logic_vector(218, 8),
60909 => conv_std_logic_vector(219, 8),
60910 => conv_std_logic_vector(220, 8),
60911 => conv_std_logic_vector(221, 8),
60912 => conv_std_logic_vector(222, 8),
60913 => conv_std_logic_vector(223, 8),
60914 => conv_std_logic_vector(224, 8),
60915 => conv_std_logic_vector(224, 8),
60916 => conv_std_logic_vector(225, 8),
60917 => conv_std_logic_vector(226, 8),
60918 => conv_std_logic_vector(227, 8),
60919 => conv_std_logic_vector(228, 8),
60920 => conv_std_logic_vector(229, 8),
60921 => conv_std_logic_vector(230, 8),
60922 => conv_std_logic_vector(231, 8),
60923 => conv_std_logic_vector(232, 8),
60924 => conv_std_logic_vector(233, 8),
60925 => conv_std_logic_vector(234, 8),
60926 => conv_std_logic_vector(235, 8),
60927 => conv_std_logic_vector(236, 8),
60928 => conv_std_logic_vector(0, 8),
60929 => conv_std_logic_vector(0, 8),
60930 => conv_std_logic_vector(1, 8),
60931 => conv_std_logic_vector(2, 8),
60932 => conv_std_logic_vector(3, 8),
60933 => conv_std_logic_vector(4, 8),
60934 => conv_std_logic_vector(5, 8),
60935 => conv_std_logic_vector(6, 8),
60936 => conv_std_logic_vector(7, 8),
60937 => conv_std_logic_vector(8, 8),
60938 => conv_std_logic_vector(9, 8),
60939 => conv_std_logic_vector(10, 8),
60940 => conv_std_logic_vector(11, 8),
60941 => conv_std_logic_vector(12, 8),
60942 => conv_std_logic_vector(13, 8),
60943 => conv_std_logic_vector(13, 8),
60944 => conv_std_logic_vector(14, 8),
60945 => conv_std_logic_vector(15, 8),
60946 => conv_std_logic_vector(16, 8),
60947 => conv_std_logic_vector(17, 8),
60948 => conv_std_logic_vector(18, 8),
60949 => conv_std_logic_vector(19, 8),
60950 => conv_std_logic_vector(20, 8),
60951 => conv_std_logic_vector(21, 8),
60952 => conv_std_logic_vector(22, 8),
60953 => conv_std_logic_vector(23, 8),
60954 => conv_std_logic_vector(24, 8),
60955 => conv_std_logic_vector(25, 8),
60956 => conv_std_logic_vector(26, 8),
60957 => conv_std_logic_vector(26, 8),
60958 => conv_std_logic_vector(27, 8),
60959 => conv_std_logic_vector(28, 8),
60960 => conv_std_logic_vector(29, 8),
60961 => conv_std_logic_vector(30, 8),
60962 => conv_std_logic_vector(31, 8),
60963 => conv_std_logic_vector(32, 8),
60964 => conv_std_logic_vector(33, 8),
60965 => conv_std_logic_vector(34, 8),
60966 => conv_std_logic_vector(35, 8),
60967 => conv_std_logic_vector(36, 8),
60968 => conv_std_logic_vector(37, 8),
60969 => conv_std_logic_vector(38, 8),
60970 => conv_std_logic_vector(39, 8),
60971 => conv_std_logic_vector(39, 8),
60972 => conv_std_logic_vector(40, 8),
60973 => conv_std_logic_vector(41, 8),
60974 => conv_std_logic_vector(42, 8),
60975 => conv_std_logic_vector(43, 8),
60976 => conv_std_logic_vector(44, 8),
60977 => conv_std_logic_vector(45, 8),
60978 => conv_std_logic_vector(46, 8),
60979 => conv_std_logic_vector(47, 8),
60980 => conv_std_logic_vector(48, 8),
60981 => conv_std_logic_vector(49, 8),
60982 => conv_std_logic_vector(50, 8),
60983 => conv_std_logic_vector(51, 8),
60984 => conv_std_logic_vector(52, 8),
60985 => conv_std_logic_vector(52, 8),
60986 => conv_std_logic_vector(53, 8),
60987 => conv_std_logic_vector(54, 8),
60988 => conv_std_logic_vector(55, 8),
60989 => conv_std_logic_vector(56, 8),
60990 => conv_std_logic_vector(57, 8),
60991 => conv_std_logic_vector(58, 8),
60992 => conv_std_logic_vector(59, 8),
60993 => conv_std_logic_vector(60, 8),
60994 => conv_std_logic_vector(61, 8),
60995 => conv_std_logic_vector(62, 8),
60996 => conv_std_logic_vector(63, 8),
60997 => conv_std_logic_vector(64, 8),
60998 => conv_std_logic_vector(65, 8),
60999 => conv_std_logic_vector(66, 8),
61000 => conv_std_logic_vector(66, 8),
61001 => conv_std_logic_vector(67, 8),
61002 => conv_std_logic_vector(68, 8),
61003 => conv_std_logic_vector(69, 8),
61004 => conv_std_logic_vector(70, 8),
61005 => conv_std_logic_vector(71, 8),
61006 => conv_std_logic_vector(72, 8),
61007 => conv_std_logic_vector(73, 8),
61008 => conv_std_logic_vector(74, 8),
61009 => conv_std_logic_vector(75, 8),
61010 => conv_std_logic_vector(76, 8),
61011 => conv_std_logic_vector(77, 8),
61012 => conv_std_logic_vector(78, 8),
61013 => conv_std_logic_vector(79, 8),
61014 => conv_std_logic_vector(79, 8),
61015 => conv_std_logic_vector(80, 8),
61016 => conv_std_logic_vector(81, 8),
61017 => conv_std_logic_vector(82, 8),
61018 => conv_std_logic_vector(83, 8),
61019 => conv_std_logic_vector(84, 8),
61020 => conv_std_logic_vector(85, 8),
61021 => conv_std_logic_vector(86, 8),
61022 => conv_std_logic_vector(87, 8),
61023 => conv_std_logic_vector(88, 8),
61024 => conv_std_logic_vector(89, 8),
61025 => conv_std_logic_vector(90, 8),
61026 => conv_std_logic_vector(91, 8),
61027 => conv_std_logic_vector(92, 8),
61028 => conv_std_logic_vector(92, 8),
61029 => conv_std_logic_vector(93, 8),
61030 => conv_std_logic_vector(94, 8),
61031 => conv_std_logic_vector(95, 8),
61032 => conv_std_logic_vector(96, 8),
61033 => conv_std_logic_vector(97, 8),
61034 => conv_std_logic_vector(98, 8),
61035 => conv_std_logic_vector(99, 8),
61036 => conv_std_logic_vector(100, 8),
61037 => conv_std_logic_vector(101, 8),
61038 => conv_std_logic_vector(102, 8),
61039 => conv_std_logic_vector(103, 8),
61040 => conv_std_logic_vector(104, 8),
61041 => conv_std_logic_vector(105, 8),
61042 => conv_std_logic_vector(105, 8),
61043 => conv_std_logic_vector(106, 8),
61044 => conv_std_logic_vector(107, 8),
61045 => conv_std_logic_vector(108, 8),
61046 => conv_std_logic_vector(109, 8),
61047 => conv_std_logic_vector(110, 8),
61048 => conv_std_logic_vector(111, 8),
61049 => conv_std_logic_vector(112, 8),
61050 => conv_std_logic_vector(113, 8),
61051 => conv_std_logic_vector(114, 8),
61052 => conv_std_logic_vector(115, 8),
61053 => conv_std_logic_vector(116, 8),
61054 => conv_std_logic_vector(117, 8),
61055 => conv_std_logic_vector(118, 8),
61056 => conv_std_logic_vector(119, 8),
61057 => conv_std_logic_vector(119, 8),
61058 => conv_std_logic_vector(120, 8),
61059 => conv_std_logic_vector(121, 8),
61060 => conv_std_logic_vector(122, 8),
61061 => conv_std_logic_vector(123, 8),
61062 => conv_std_logic_vector(124, 8),
61063 => conv_std_logic_vector(125, 8),
61064 => conv_std_logic_vector(126, 8),
61065 => conv_std_logic_vector(127, 8),
61066 => conv_std_logic_vector(128, 8),
61067 => conv_std_logic_vector(129, 8),
61068 => conv_std_logic_vector(130, 8),
61069 => conv_std_logic_vector(131, 8),
61070 => conv_std_logic_vector(132, 8),
61071 => conv_std_logic_vector(132, 8),
61072 => conv_std_logic_vector(133, 8),
61073 => conv_std_logic_vector(134, 8),
61074 => conv_std_logic_vector(135, 8),
61075 => conv_std_logic_vector(136, 8),
61076 => conv_std_logic_vector(137, 8),
61077 => conv_std_logic_vector(138, 8),
61078 => conv_std_logic_vector(139, 8),
61079 => conv_std_logic_vector(140, 8),
61080 => conv_std_logic_vector(141, 8),
61081 => conv_std_logic_vector(142, 8),
61082 => conv_std_logic_vector(143, 8),
61083 => conv_std_logic_vector(144, 8),
61084 => conv_std_logic_vector(145, 8),
61085 => conv_std_logic_vector(145, 8),
61086 => conv_std_logic_vector(146, 8),
61087 => conv_std_logic_vector(147, 8),
61088 => conv_std_logic_vector(148, 8),
61089 => conv_std_logic_vector(149, 8),
61090 => conv_std_logic_vector(150, 8),
61091 => conv_std_logic_vector(151, 8),
61092 => conv_std_logic_vector(152, 8),
61093 => conv_std_logic_vector(153, 8),
61094 => conv_std_logic_vector(154, 8),
61095 => conv_std_logic_vector(155, 8),
61096 => conv_std_logic_vector(156, 8),
61097 => conv_std_logic_vector(157, 8),
61098 => conv_std_logic_vector(158, 8),
61099 => conv_std_logic_vector(158, 8),
61100 => conv_std_logic_vector(159, 8),
61101 => conv_std_logic_vector(160, 8),
61102 => conv_std_logic_vector(161, 8),
61103 => conv_std_logic_vector(162, 8),
61104 => conv_std_logic_vector(163, 8),
61105 => conv_std_logic_vector(164, 8),
61106 => conv_std_logic_vector(165, 8),
61107 => conv_std_logic_vector(166, 8),
61108 => conv_std_logic_vector(167, 8),
61109 => conv_std_logic_vector(168, 8),
61110 => conv_std_logic_vector(169, 8),
61111 => conv_std_logic_vector(170, 8),
61112 => conv_std_logic_vector(171, 8),
61113 => conv_std_logic_vector(171, 8),
61114 => conv_std_logic_vector(172, 8),
61115 => conv_std_logic_vector(173, 8),
61116 => conv_std_logic_vector(174, 8),
61117 => conv_std_logic_vector(175, 8),
61118 => conv_std_logic_vector(176, 8),
61119 => conv_std_logic_vector(177, 8),
61120 => conv_std_logic_vector(178, 8),
61121 => conv_std_logic_vector(179, 8),
61122 => conv_std_logic_vector(180, 8),
61123 => conv_std_logic_vector(181, 8),
61124 => conv_std_logic_vector(182, 8),
61125 => conv_std_logic_vector(183, 8),
61126 => conv_std_logic_vector(184, 8),
61127 => conv_std_logic_vector(185, 8),
61128 => conv_std_logic_vector(185, 8),
61129 => conv_std_logic_vector(186, 8),
61130 => conv_std_logic_vector(187, 8),
61131 => conv_std_logic_vector(188, 8),
61132 => conv_std_logic_vector(189, 8),
61133 => conv_std_logic_vector(190, 8),
61134 => conv_std_logic_vector(191, 8),
61135 => conv_std_logic_vector(192, 8),
61136 => conv_std_logic_vector(193, 8),
61137 => conv_std_logic_vector(194, 8),
61138 => conv_std_logic_vector(195, 8),
61139 => conv_std_logic_vector(196, 8),
61140 => conv_std_logic_vector(197, 8),
61141 => conv_std_logic_vector(198, 8),
61142 => conv_std_logic_vector(198, 8),
61143 => conv_std_logic_vector(199, 8),
61144 => conv_std_logic_vector(200, 8),
61145 => conv_std_logic_vector(201, 8),
61146 => conv_std_logic_vector(202, 8),
61147 => conv_std_logic_vector(203, 8),
61148 => conv_std_logic_vector(204, 8),
61149 => conv_std_logic_vector(205, 8),
61150 => conv_std_logic_vector(206, 8),
61151 => conv_std_logic_vector(207, 8),
61152 => conv_std_logic_vector(208, 8),
61153 => conv_std_logic_vector(209, 8),
61154 => conv_std_logic_vector(210, 8),
61155 => conv_std_logic_vector(211, 8),
61156 => conv_std_logic_vector(211, 8),
61157 => conv_std_logic_vector(212, 8),
61158 => conv_std_logic_vector(213, 8),
61159 => conv_std_logic_vector(214, 8),
61160 => conv_std_logic_vector(215, 8),
61161 => conv_std_logic_vector(216, 8),
61162 => conv_std_logic_vector(217, 8),
61163 => conv_std_logic_vector(218, 8),
61164 => conv_std_logic_vector(219, 8),
61165 => conv_std_logic_vector(220, 8),
61166 => conv_std_logic_vector(221, 8),
61167 => conv_std_logic_vector(222, 8),
61168 => conv_std_logic_vector(223, 8),
61169 => conv_std_logic_vector(224, 8),
61170 => conv_std_logic_vector(224, 8),
61171 => conv_std_logic_vector(225, 8),
61172 => conv_std_logic_vector(226, 8),
61173 => conv_std_logic_vector(227, 8),
61174 => conv_std_logic_vector(228, 8),
61175 => conv_std_logic_vector(229, 8),
61176 => conv_std_logic_vector(230, 8),
61177 => conv_std_logic_vector(231, 8),
61178 => conv_std_logic_vector(232, 8),
61179 => conv_std_logic_vector(233, 8),
61180 => conv_std_logic_vector(234, 8),
61181 => conv_std_logic_vector(235, 8),
61182 => conv_std_logic_vector(236, 8),
61183 => conv_std_logic_vector(237, 8),
61184 => conv_std_logic_vector(0, 8),
61185 => conv_std_logic_vector(0, 8),
61186 => conv_std_logic_vector(1, 8),
61187 => conv_std_logic_vector(2, 8),
61188 => conv_std_logic_vector(3, 8),
61189 => conv_std_logic_vector(4, 8),
61190 => conv_std_logic_vector(5, 8),
61191 => conv_std_logic_vector(6, 8),
61192 => conv_std_logic_vector(7, 8),
61193 => conv_std_logic_vector(8, 8),
61194 => conv_std_logic_vector(9, 8),
61195 => conv_std_logic_vector(10, 8),
61196 => conv_std_logic_vector(11, 8),
61197 => conv_std_logic_vector(12, 8),
61198 => conv_std_logic_vector(13, 8),
61199 => conv_std_logic_vector(14, 8),
61200 => conv_std_logic_vector(14, 8),
61201 => conv_std_logic_vector(15, 8),
61202 => conv_std_logic_vector(16, 8),
61203 => conv_std_logic_vector(17, 8),
61204 => conv_std_logic_vector(18, 8),
61205 => conv_std_logic_vector(19, 8),
61206 => conv_std_logic_vector(20, 8),
61207 => conv_std_logic_vector(21, 8),
61208 => conv_std_logic_vector(22, 8),
61209 => conv_std_logic_vector(23, 8),
61210 => conv_std_logic_vector(24, 8),
61211 => conv_std_logic_vector(25, 8),
61212 => conv_std_logic_vector(26, 8),
61213 => conv_std_logic_vector(27, 8),
61214 => conv_std_logic_vector(28, 8),
61215 => conv_std_logic_vector(28, 8),
61216 => conv_std_logic_vector(29, 8),
61217 => conv_std_logic_vector(30, 8),
61218 => conv_std_logic_vector(31, 8),
61219 => conv_std_logic_vector(32, 8),
61220 => conv_std_logic_vector(33, 8),
61221 => conv_std_logic_vector(34, 8),
61222 => conv_std_logic_vector(35, 8),
61223 => conv_std_logic_vector(36, 8),
61224 => conv_std_logic_vector(37, 8),
61225 => conv_std_logic_vector(38, 8),
61226 => conv_std_logic_vector(39, 8),
61227 => conv_std_logic_vector(40, 8),
61228 => conv_std_logic_vector(41, 8),
61229 => conv_std_logic_vector(42, 8),
61230 => conv_std_logic_vector(42, 8),
61231 => conv_std_logic_vector(43, 8),
61232 => conv_std_logic_vector(44, 8),
61233 => conv_std_logic_vector(45, 8),
61234 => conv_std_logic_vector(46, 8),
61235 => conv_std_logic_vector(47, 8),
61236 => conv_std_logic_vector(48, 8),
61237 => conv_std_logic_vector(49, 8),
61238 => conv_std_logic_vector(50, 8),
61239 => conv_std_logic_vector(51, 8),
61240 => conv_std_logic_vector(52, 8),
61241 => conv_std_logic_vector(53, 8),
61242 => conv_std_logic_vector(54, 8),
61243 => conv_std_logic_vector(55, 8),
61244 => conv_std_logic_vector(56, 8),
61245 => conv_std_logic_vector(56, 8),
61246 => conv_std_logic_vector(57, 8),
61247 => conv_std_logic_vector(58, 8),
61248 => conv_std_logic_vector(59, 8),
61249 => conv_std_logic_vector(60, 8),
61250 => conv_std_logic_vector(61, 8),
61251 => conv_std_logic_vector(62, 8),
61252 => conv_std_logic_vector(63, 8),
61253 => conv_std_logic_vector(64, 8),
61254 => conv_std_logic_vector(65, 8),
61255 => conv_std_logic_vector(66, 8),
61256 => conv_std_logic_vector(67, 8),
61257 => conv_std_logic_vector(68, 8),
61258 => conv_std_logic_vector(69, 8),
61259 => conv_std_logic_vector(70, 8),
61260 => conv_std_logic_vector(70, 8),
61261 => conv_std_logic_vector(71, 8),
61262 => conv_std_logic_vector(72, 8),
61263 => conv_std_logic_vector(73, 8),
61264 => conv_std_logic_vector(74, 8),
61265 => conv_std_logic_vector(75, 8),
61266 => conv_std_logic_vector(76, 8),
61267 => conv_std_logic_vector(77, 8),
61268 => conv_std_logic_vector(78, 8),
61269 => conv_std_logic_vector(79, 8),
61270 => conv_std_logic_vector(80, 8),
61271 => conv_std_logic_vector(81, 8),
61272 => conv_std_logic_vector(82, 8),
61273 => conv_std_logic_vector(83, 8),
61274 => conv_std_logic_vector(84, 8),
61275 => conv_std_logic_vector(84, 8),
61276 => conv_std_logic_vector(85, 8),
61277 => conv_std_logic_vector(86, 8),
61278 => conv_std_logic_vector(87, 8),
61279 => conv_std_logic_vector(88, 8),
61280 => conv_std_logic_vector(89, 8),
61281 => conv_std_logic_vector(90, 8),
61282 => conv_std_logic_vector(91, 8),
61283 => conv_std_logic_vector(92, 8),
61284 => conv_std_logic_vector(93, 8),
61285 => conv_std_logic_vector(94, 8),
61286 => conv_std_logic_vector(95, 8),
61287 => conv_std_logic_vector(96, 8),
61288 => conv_std_logic_vector(97, 8),
61289 => conv_std_logic_vector(98, 8),
61290 => conv_std_logic_vector(98, 8),
61291 => conv_std_logic_vector(99, 8),
61292 => conv_std_logic_vector(100, 8),
61293 => conv_std_logic_vector(101, 8),
61294 => conv_std_logic_vector(102, 8),
61295 => conv_std_logic_vector(103, 8),
61296 => conv_std_logic_vector(104, 8),
61297 => conv_std_logic_vector(105, 8),
61298 => conv_std_logic_vector(106, 8),
61299 => conv_std_logic_vector(107, 8),
61300 => conv_std_logic_vector(108, 8),
61301 => conv_std_logic_vector(109, 8),
61302 => conv_std_logic_vector(110, 8),
61303 => conv_std_logic_vector(111, 8),
61304 => conv_std_logic_vector(112, 8),
61305 => conv_std_logic_vector(112, 8),
61306 => conv_std_logic_vector(113, 8),
61307 => conv_std_logic_vector(114, 8),
61308 => conv_std_logic_vector(115, 8),
61309 => conv_std_logic_vector(116, 8),
61310 => conv_std_logic_vector(117, 8),
61311 => conv_std_logic_vector(118, 8),
61312 => conv_std_logic_vector(119, 8),
61313 => conv_std_logic_vector(120, 8),
61314 => conv_std_logic_vector(121, 8),
61315 => conv_std_logic_vector(122, 8),
61316 => conv_std_logic_vector(123, 8),
61317 => conv_std_logic_vector(124, 8),
61318 => conv_std_logic_vector(125, 8),
61319 => conv_std_logic_vector(126, 8),
61320 => conv_std_logic_vector(126, 8),
61321 => conv_std_logic_vector(127, 8),
61322 => conv_std_logic_vector(128, 8),
61323 => conv_std_logic_vector(129, 8),
61324 => conv_std_logic_vector(130, 8),
61325 => conv_std_logic_vector(131, 8),
61326 => conv_std_logic_vector(132, 8),
61327 => conv_std_logic_vector(133, 8),
61328 => conv_std_logic_vector(134, 8),
61329 => conv_std_logic_vector(135, 8),
61330 => conv_std_logic_vector(136, 8),
61331 => conv_std_logic_vector(137, 8),
61332 => conv_std_logic_vector(138, 8),
61333 => conv_std_logic_vector(139, 8),
61334 => conv_std_logic_vector(140, 8),
61335 => conv_std_logic_vector(140, 8),
61336 => conv_std_logic_vector(141, 8),
61337 => conv_std_logic_vector(142, 8),
61338 => conv_std_logic_vector(143, 8),
61339 => conv_std_logic_vector(144, 8),
61340 => conv_std_logic_vector(145, 8),
61341 => conv_std_logic_vector(146, 8),
61342 => conv_std_logic_vector(147, 8),
61343 => conv_std_logic_vector(148, 8),
61344 => conv_std_logic_vector(149, 8),
61345 => conv_std_logic_vector(150, 8),
61346 => conv_std_logic_vector(151, 8),
61347 => conv_std_logic_vector(152, 8),
61348 => conv_std_logic_vector(153, 8),
61349 => conv_std_logic_vector(154, 8),
61350 => conv_std_logic_vector(154, 8),
61351 => conv_std_logic_vector(155, 8),
61352 => conv_std_logic_vector(156, 8),
61353 => conv_std_logic_vector(157, 8),
61354 => conv_std_logic_vector(158, 8),
61355 => conv_std_logic_vector(159, 8),
61356 => conv_std_logic_vector(160, 8),
61357 => conv_std_logic_vector(161, 8),
61358 => conv_std_logic_vector(162, 8),
61359 => conv_std_logic_vector(163, 8),
61360 => conv_std_logic_vector(164, 8),
61361 => conv_std_logic_vector(165, 8),
61362 => conv_std_logic_vector(166, 8),
61363 => conv_std_logic_vector(167, 8),
61364 => conv_std_logic_vector(168, 8),
61365 => conv_std_logic_vector(168, 8),
61366 => conv_std_logic_vector(169, 8),
61367 => conv_std_logic_vector(170, 8),
61368 => conv_std_logic_vector(171, 8),
61369 => conv_std_logic_vector(172, 8),
61370 => conv_std_logic_vector(173, 8),
61371 => conv_std_logic_vector(174, 8),
61372 => conv_std_logic_vector(175, 8),
61373 => conv_std_logic_vector(176, 8),
61374 => conv_std_logic_vector(177, 8),
61375 => conv_std_logic_vector(178, 8),
61376 => conv_std_logic_vector(179, 8),
61377 => conv_std_logic_vector(180, 8),
61378 => conv_std_logic_vector(181, 8),
61379 => conv_std_logic_vector(182, 8),
61380 => conv_std_logic_vector(182, 8),
61381 => conv_std_logic_vector(183, 8),
61382 => conv_std_logic_vector(184, 8),
61383 => conv_std_logic_vector(185, 8),
61384 => conv_std_logic_vector(186, 8),
61385 => conv_std_logic_vector(187, 8),
61386 => conv_std_logic_vector(188, 8),
61387 => conv_std_logic_vector(189, 8),
61388 => conv_std_logic_vector(190, 8),
61389 => conv_std_logic_vector(191, 8),
61390 => conv_std_logic_vector(192, 8),
61391 => conv_std_logic_vector(193, 8),
61392 => conv_std_logic_vector(194, 8),
61393 => conv_std_logic_vector(195, 8),
61394 => conv_std_logic_vector(196, 8),
61395 => conv_std_logic_vector(196, 8),
61396 => conv_std_logic_vector(197, 8),
61397 => conv_std_logic_vector(198, 8),
61398 => conv_std_logic_vector(199, 8),
61399 => conv_std_logic_vector(200, 8),
61400 => conv_std_logic_vector(201, 8),
61401 => conv_std_logic_vector(202, 8),
61402 => conv_std_logic_vector(203, 8),
61403 => conv_std_logic_vector(204, 8),
61404 => conv_std_logic_vector(205, 8),
61405 => conv_std_logic_vector(206, 8),
61406 => conv_std_logic_vector(207, 8),
61407 => conv_std_logic_vector(208, 8),
61408 => conv_std_logic_vector(209, 8),
61409 => conv_std_logic_vector(210, 8),
61410 => conv_std_logic_vector(210, 8),
61411 => conv_std_logic_vector(211, 8),
61412 => conv_std_logic_vector(212, 8),
61413 => conv_std_logic_vector(213, 8),
61414 => conv_std_logic_vector(214, 8),
61415 => conv_std_logic_vector(215, 8),
61416 => conv_std_logic_vector(216, 8),
61417 => conv_std_logic_vector(217, 8),
61418 => conv_std_logic_vector(218, 8),
61419 => conv_std_logic_vector(219, 8),
61420 => conv_std_logic_vector(220, 8),
61421 => conv_std_logic_vector(221, 8),
61422 => conv_std_logic_vector(222, 8),
61423 => conv_std_logic_vector(223, 8),
61424 => conv_std_logic_vector(224, 8),
61425 => conv_std_logic_vector(224, 8),
61426 => conv_std_logic_vector(225, 8),
61427 => conv_std_logic_vector(226, 8),
61428 => conv_std_logic_vector(227, 8),
61429 => conv_std_logic_vector(228, 8),
61430 => conv_std_logic_vector(229, 8),
61431 => conv_std_logic_vector(230, 8),
61432 => conv_std_logic_vector(231, 8),
61433 => conv_std_logic_vector(232, 8),
61434 => conv_std_logic_vector(233, 8),
61435 => conv_std_logic_vector(234, 8),
61436 => conv_std_logic_vector(235, 8),
61437 => conv_std_logic_vector(236, 8),
61438 => conv_std_logic_vector(237, 8),
61439 => conv_std_logic_vector(238, 8),
61440 => conv_std_logic_vector(0, 8),
61441 => conv_std_logic_vector(0, 8),
61442 => conv_std_logic_vector(1, 8),
61443 => conv_std_logic_vector(2, 8),
61444 => conv_std_logic_vector(3, 8),
61445 => conv_std_logic_vector(4, 8),
61446 => conv_std_logic_vector(5, 8),
61447 => conv_std_logic_vector(6, 8),
61448 => conv_std_logic_vector(7, 8),
61449 => conv_std_logic_vector(8, 8),
61450 => conv_std_logic_vector(9, 8),
61451 => conv_std_logic_vector(10, 8),
61452 => conv_std_logic_vector(11, 8),
61453 => conv_std_logic_vector(12, 8),
61454 => conv_std_logic_vector(13, 8),
61455 => conv_std_logic_vector(14, 8),
61456 => conv_std_logic_vector(15, 8),
61457 => conv_std_logic_vector(15, 8),
61458 => conv_std_logic_vector(16, 8),
61459 => conv_std_logic_vector(17, 8),
61460 => conv_std_logic_vector(18, 8),
61461 => conv_std_logic_vector(19, 8),
61462 => conv_std_logic_vector(20, 8),
61463 => conv_std_logic_vector(21, 8),
61464 => conv_std_logic_vector(22, 8),
61465 => conv_std_logic_vector(23, 8),
61466 => conv_std_logic_vector(24, 8),
61467 => conv_std_logic_vector(25, 8),
61468 => conv_std_logic_vector(26, 8),
61469 => conv_std_logic_vector(27, 8),
61470 => conv_std_logic_vector(28, 8),
61471 => conv_std_logic_vector(29, 8),
61472 => conv_std_logic_vector(30, 8),
61473 => conv_std_logic_vector(30, 8),
61474 => conv_std_logic_vector(31, 8),
61475 => conv_std_logic_vector(32, 8),
61476 => conv_std_logic_vector(33, 8),
61477 => conv_std_logic_vector(34, 8),
61478 => conv_std_logic_vector(35, 8),
61479 => conv_std_logic_vector(36, 8),
61480 => conv_std_logic_vector(37, 8),
61481 => conv_std_logic_vector(38, 8),
61482 => conv_std_logic_vector(39, 8),
61483 => conv_std_logic_vector(40, 8),
61484 => conv_std_logic_vector(41, 8),
61485 => conv_std_logic_vector(42, 8),
61486 => conv_std_logic_vector(43, 8),
61487 => conv_std_logic_vector(44, 8),
61488 => conv_std_logic_vector(45, 8),
61489 => conv_std_logic_vector(45, 8),
61490 => conv_std_logic_vector(46, 8),
61491 => conv_std_logic_vector(47, 8),
61492 => conv_std_logic_vector(48, 8),
61493 => conv_std_logic_vector(49, 8),
61494 => conv_std_logic_vector(50, 8),
61495 => conv_std_logic_vector(51, 8),
61496 => conv_std_logic_vector(52, 8),
61497 => conv_std_logic_vector(53, 8),
61498 => conv_std_logic_vector(54, 8),
61499 => conv_std_logic_vector(55, 8),
61500 => conv_std_logic_vector(56, 8),
61501 => conv_std_logic_vector(57, 8),
61502 => conv_std_logic_vector(58, 8),
61503 => conv_std_logic_vector(59, 8),
61504 => conv_std_logic_vector(60, 8),
61505 => conv_std_logic_vector(60, 8),
61506 => conv_std_logic_vector(61, 8),
61507 => conv_std_logic_vector(62, 8),
61508 => conv_std_logic_vector(63, 8),
61509 => conv_std_logic_vector(64, 8),
61510 => conv_std_logic_vector(65, 8),
61511 => conv_std_logic_vector(66, 8),
61512 => conv_std_logic_vector(67, 8),
61513 => conv_std_logic_vector(68, 8),
61514 => conv_std_logic_vector(69, 8),
61515 => conv_std_logic_vector(70, 8),
61516 => conv_std_logic_vector(71, 8),
61517 => conv_std_logic_vector(72, 8),
61518 => conv_std_logic_vector(73, 8),
61519 => conv_std_logic_vector(74, 8),
61520 => conv_std_logic_vector(75, 8),
61521 => conv_std_logic_vector(75, 8),
61522 => conv_std_logic_vector(76, 8),
61523 => conv_std_logic_vector(77, 8),
61524 => conv_std_logic_vector(78, 8),
61525 => conv_std_logic_vector(79, 8),
61526 => conv_std_logic_vector(80, 8),
61527 => conv_std_logic_vector(81, 8),
61528 => conv_std_logic_vector(82, 8),
61529 => conv_std_logic_vector(83, 8),
61530 => conv_std_logic_vector(84, 8),
61531 => conv_std_logic_vector(85, 8),
61532 => conv_std_logic_vector(86, 8),
61533 => conv_std_logic_vector(87, 8),
61534 => conv_std_logic_vector(88, 8),
61535 => conv_std_logic_vector(89, 8),
61536 => conv_std_logic_vector(90, 8),
61537 => conv_std_logic_vector(90, 8),
61538 => conv_std_logic_vector(91, 8),
61539 => conv_std_logic_vector(92, 8),
61540 => conv_std_logic_vector(93, 8),
61541 => conv_std_logic_vector(94, 8),
61542 => conv_std_logic_vector(95, 8),
61543 => conv_std_logic_vector(96, 8),
61544 => conv_std_logic_vector(97, 8),
61545 => conv_std_logic_vector(98, 8),
61546 => conv_std_logic_vector(99, 8),
61547 => conv_std_logic_vector(100, 8),
61548 => conv_std_logic_vector(101, 8),
61549 => conv_std_logic_vector(102, 8),
61550 => conv_std_logic_vector(103, 8),
61551 => conv_std_logic_vector(104, 8),
61552 => conv_std_logic_vector(105, 8),
61553 => conv_std_logic_vector(105, 8),
61554 => conv_std_logic_vector(106, 8),
61555 => conv_std_logic_vector(107, 8),
61556 => conv_std_logic_vector(108, 8),
61557 => conv_std_logic_vector(109, 8),
61558 => conv_std_logic_vector(110, 8),
61559 => conv_std_logic_vector(111, 8),
61560 => conv_std_logic_vector(112, 8),
61561 => conv_std_logic_vector(113, 8),
61562 => conv_std_logic_vector(114, 8),
61563 => conv_std_logic_vector(115, 8),
61564 => conv_std_logic_vector(116, 8),
61565 => conv_std_logic_vector(117, 8),
61566 => conv_std_logic_vector(118, 8),
61567 => conv_std_logic_vector(119, 8),
61568 => conv_std_logic_vector(120, 8),
61569 => conv_std_logic_vector(120, 8),
61570 => conv_std_logic_vector(121, 8),
61571 => conv_std_logic_vector(122, 8),
61572 => conv_std_logic_vector(123, 8),
61573 => conv_std_logic_vector(124, 8),
61574 => conv_std_logic_vector(125, 8),
61575 => conv_std_logic_vector(126, 8),
61576 => conv_std_logic_vector(127, 8),
61577 => conv_std_logic_vector(128, 8),
61578 => conv_std_logic_vector(129, 8),
61579 => conv_std_logic_vector(130, 8),
61580 => conv_std_logic_vector(131, 8),
61581 => conv_std_logic_vector(132, 8),
61582 => conv_std_logic_vector(133, 8),
61583 => conv_std_logic_vector(134, 8),
61584 => conv_std_logic_vector(135, 8),
61585 => conv_std_logic_vector(135, 8),
61586 => conv_std_logic_vector(136, 8),
61587 => conv_std_logic_vector(137, 8),
61588 => conv_std_logic_vector(138, 8),
61589 => conv_std_logic_vector(139, 8),
61590 => conv_std_logic_vector(140, 8),
61591 => conv_std_logic_vector(141, 8),
61592 => conv_std_logic_vector(142, 8),
61593 => conv_std_logic_vector(143, 8),
61594 => conv_std_logic_vector(144, 8),
61595 => conv_std_logic_vector(145, 8),
61596 => conv_std_logic_vector(146, 8),
61597 => conv_std_logic_vector(147, 8),
61598 => conv_std_logic_vector(148, 8),
61599 => conv_std_logic_vector(149, 8),
61600 => conv_std_logic_vector(150, 8),
61601 => conv_std_logic_vector(150, 8),
61602 => conv_std_logic_vector(151, 8),
61603 => conv_std_logic_vector(152, 8),
61604 => conv_std_logic_vector(153, 8),
61605 => conv_std_logic_vector(154, 8),
61606 => conv_std_logic_vector(155, 8),
61607 => conv_std_logic_vector(156, 8),
61608 => conv_std_logic_vector(157, 8),
61609 => conv_std_logic_vector(158, 8),
61610 => conv_std_logic_vector(159, 8),
61611 => conv_std_logic_vector(160, 8),
61612 => conv_std_logic_vector(161, 8),
61613 => conv_std_logic_vector(162, 8),
61614 => conv_std_logic_vector(163, 8),
61615 => conv_std_logic_vector(164, 8),
61616 => conv_std_logic_vector(165, 8),
61617 => conv_std_logic_vector(165, 8),
61618 => conv_std_logic_vector(166, 8),
61619 => conv_std_logic_vector(167, 8),
61620 => conv_std_logic_vector(168, 8),
61621 => conv_std_logic_vector(169, 8),
61622 => conv_std_logic_vector(170, 8),
61623 => conv_std_logic_vector(171, 8),
61624 => conv_std_logic_vector(172, 8),
61625 => conv_std_logic_vector(173, 8),
61626 => conv_std_logic_vector(174, 8),
61627 => conv_std_logic_vector(175, 8),
61628 => conv_std_logic_vector(176, 8),
61629 => conv_std_logic_vector(177, 8),
61630 => conv_std_logic_vector(178, 8),
61631 => conv_std_logic_vector(179, 8),
61632 => conv_std_logic_vector(180, 8),
61633 => conv_std_logic_vector(180, 8),
61634 => conv_std_logic_vector(181, 8),
61635 => conv_std_logic_vector(182, 8),
61636 => conv_std_logic_vector(183, 8),
61637 => conv_std_logic_vector(184, 8),
61638 => conv_std_logic_vector(185, 8),
61639 => conv_std_logic_vector(186, 8),
61640 => conv_std_logic_vector(187, 8),
61641 => conv_std_logic_vector(188, 8),
61642 => conv_std_logic_vector(189, 8),
61643 => conv_std_logic_vector(190, 8),
61644 => conv_std_logic_vector(191, 8),
61645 => conv_std_logic_vector(192, 8),
61646 => conv_std_logic_vector(193, 8),
61647 => conv_std_logic_vector(194, 8),
61648 => conv_std_logic_vector(195, 8),
61649 => conv_std_logic_vector(195, 8),
61650 => conv_std_logic_vector(196, 8),
61651 => conv_std_logic_vector(197, 8),
61652 => conv_std_logic_vector(198, 8),
61653 => conv_std_logic_vector(199, 8),
61654 => conv_std_logic_vector(200, 8),
61655 => conv_std_logic_vector(201, 8),
61656 => conv_std_logic_vector(202, 8),
61657 => conv_std_logic_vector(203, 8),
61658 => conv_std_logic_vector(204, 8),
61659 => conv_std_logic_vector(205, 8),
61660 => conv_std_logic_vector(206, 8),
61661 => conv_std_logic_vector(207, 8),
61662 => conv_std_logic_vector(208, 8),
61663 => conv_std_logic_vector(209, 8),
61664 => conv_std_logic_vector(210, 8),
61665 => conv_std_logic_vector(210, 8),
61666 => conv_std_logic_vector(211, 8),
61667 => conv_std_logic_vector(212, 8),
61668 => conv_std_logic_vector(213, 8),
61669 => conv_std_logic_vector(214, 8),
61670 => conv_std_logic_vector(215, 8),
61671 => conv_std_logic_vector(216, 8),
61672 => conv_std_logic_vector(217, 8),
61673 => conv_std_logic_vector(218, 8),
61674 => conv_std_logic_vector(219, 8),
61675 => conv_std_logic_vector(220, 8),
61676 => conv_std_logic_vector(221, 8),
61677 => conv_std_logic_vector(222, 8),
61678 => conv_std_logic_vector(223, 8),
61679 => conv_std_logic_vector(224, 8),
61680 => conv_std_logic_vector(225, 8),
61681 => conv_std_logic_vector(225, 8),
61682 => conv_std_logic_vector(226, 8),
61683 => conv_std_logic_vector(227, 8),
61684 => conv_std_logic_vector(228, 8),
61685 => conv_std_logic_vector(229, 8),
61686 => conv_std_logic_vector(230, 8),
61687 => conv_std_logic_vector(231, 8),
61688 => conv_std_logic_vector(232, 8),
61689 => conv_std_logic_vector(233, 8),
61690 => conv_std_logic_vector(234, 8),
61691 => conv_std_logic_vector(235, 8),
61692 => conv_std_logic_vector(236, 8),
61693 => conv_std_logic_vector(237, 8),
61694 => conv_std_logic_vector(238, 8),
61695 => conv_std_logic_vector(239, 8),
61696 => conv_std_logic_vector(0, 8),
61697 => conv_std_logic_vector(0, 8),
61698 => conv_std_logic_vector(1, 8),
61699 => conv_std_logic_vector(2, 8),
61700 => conv_std_logic_vector(3, 8),
61701 => conv_std_logic_vector(4, 8),
61702 => conv_std_logic_vector(5, 8),
61703 => conv_std_logic_vector(6, 8),
61704 => conv_std_logic_vector(7, 8),
61705 => conv_std_logic_vector(8, 8),
61706 => conv_std_logic_vector(9, 8),
61707 => conv_std_logic_vector(10, 8),
61708 => conv_std_logic_vector(11, 8),
61709 => conv_std_logic_vector(12, 8),
61710 => conv_std_logic_vector(13, 8),
61711 => conv_std_logic_vector(14, 8),
61712 => conv_std_logic_vector(15, 8),
61713 => conv_std_logic_vector(16, 8),
61714 => conv_std_logic_vector(16, 8),
61715 => conv_std_logic_vector(17, 8),
61716 => conv_std_logic_vector(18, 8),
61717 => conv_std_logic_vector(19, 8),
61718 => conv_std_logic_vector(20, 8),
61719 => conv_std_logic_vector(21, 8),
61720 => conv_std_logic_vector(22, 8),
61721 => conv_std_logic_vector(23, 8),
61722 => conv_std_logic_vector(24, 8),
61723 => conv_std_logic_vector(25, 8),
61724 => conv_std_logic_vector(26, 8),
61725 => conv_std_logic_vector(27, 8),
61726 => conv_std_logic_vector(28, 8),
61727 => conv_std_logic_vector(29, 8),
61728 => conv_std_logic_vector(30, 8),
61729 => conv_std_logic_vector(31, 8),
61730 => conv_std_logic_vector(32, 8),
61731 => conv_std_logic_vector(32, 8),
61732 => conv_std_logic_vector(33, 8),
61733 => conv_std_logic_vector(34, 8),
61734 => conv_std_logic_vector(35, 8),
61735 => conv_std_logic_vector(36, 8),
61736 => conv_std_logic_vector(37, 8),
61737 => conv_std_logic_vector(38, 8),
61738 => conv_std_logic_vector(39, 8),
61739 => conv_std_logic_vector(40, 8),
61740 => conv_std_logic_vector(41, 8),
61741 => conv_std_logic_vector(42, 8),
61742 => conv_std_logic_vector(43, 8),
61743 => conv_std_logic_vector(44, 8),
61744 => conv_std_logic_vector(45, 8),
61745 => conv_std_logic_vector(46, 8),
61746 => conv_std_logic_vector(47, 8),
61747 => conv_std_logic_vector(48, 8),
61748 => conv_std_logic_vector(48, 8),
61749 => conv_std_logic_vector(49, 8),
61750 => conv_std_logic_vector(50, 8),
61751 => conv_std_logic_vector(51, 8),
61752 => conv_std_logic_vector(52, 8),
61753 => conv_std_logic_vector(53, 8),
61754 => conv_std_logic_vector(54, 8),
61755 => conv_std_logic_vector(55, 8),
61756 => conv_std_logic_vector(56, 8),
61757 => conv_std_logic_vector(57, 8),
61758 => conv_std_logic_vector(58, 8),
61759 => conv_std_logic_vector(59, 8),
61760 => conv_std_logic_vector(60, 8),
61761 => conv_std_logic_vector(61, 8),
61762 => conv_std_logic_vector(62, 8),
61763 => conv_std_logic_vector(63, 8),
61764 => conv_std_logic_vector(64, 8),
61765 => conv_std_logic_vector(64, 8),
61766 => conv_std_logic_vector(65, 8),
61767 => conv_std_logic_vector(66, 8),
61768 => conv_std_logic_vector(67, 8),
61769 => conv_std_logic_vector(68, 8),
61770 => conv_std_logic_vector(69, 8),
61771 => conv_std_logic_vector(70, 8),
61772 => conv_std_logic_vector(71, 8),
61773 => conv_std_logic_vector(72, 8),
61774 => conv_std_logic_vector(73, 8),
61775 => conv_std_logic_vector(74, 8),
61776 => conv_std_logic_vector(75, 8),
61777 => conv_std_logic_vector(76, 8),
61778 => conv_std_logic_vector(77, 8),
61779 => conv_std_logic_vector(78, 8),
61780 => conv_std_logic_vector(79, 8),
61781 => conv_std_logic_vector(80, 8),
61782 => conv_std_logic_vector(80, 8),
61783 => conv_std_logic_vector(81, 8),
61784 => conv_std_logic_vector(82, 8),
61785 => conv_std_logic_vector(83, 8),
61786 => conv_std_logic_vector(84, 8),
61787 => conv_std_logic_vector(85, 8),
61788 => conv_std_logic_vector(86, 8),
61789 => conv_std_logic_vector(87, 8),
61790 => conv_std_logic_vector(88, 8),
61791 => conv_std_logic_vector(89, 8),
61792 => conv_std_logic_vector(90, 8),
61793 => conv_std_logic_vector(91, 8),
61794 => conv_std_logic_vector(92, 8),
61795 => conv_std_logic_vector(93, 8),
61796 => conv_std_logic_vector(94, 8),
61797 => conv_std_logic_vector(95, 8),
61798 => conv_std_logic_vector(96, 8),
61799 => conv_std_logic_vector(96, 8),
61800 => conv_std_logic_vector(97, 8),
61801 => conv_std_logic_vector(98, 8),
61802 => conv_std_logic_vector(99, 8),
61803 => conv_std_logic_vector(100, 8),
61804 => conv_std_logic_vector(101, 8),
61805 => conv_std_logic_vector(102, 8),
61806 => conv_std_logic_vector(103, 8),
61807 => conv_std_logic_vector(104, 8),
61808 => conv_std_logic_vector(105, 8),
61809 => conv_std_logic_vector(106, 8),
61810 => conv_std_logic_vector(107, 8),
61811 => conv_std_logic_vector(108, 8),
61812 => conv_std_logic_vector(109, 8),
61813 => conv_std_logic_vector(110, 8),
61814 => conv_std_logic_vector(111, 8),
61815 => conv_std_logic_vector(112, 8),
61816 => conv_std_logic_vector(112, 8),
61817 => conv_std_logic_vector(113, 8),
61818 => conv_std_logic_vector(114, 8),
61819 => conv_std_logic_vector(115, 8),
61820 => conv_std_logic_vector(116, 8),
61821 => conv_std_logic_vector(117, 8),
61822 => conv_std_logic_vector(118, 8),
61823 => conv_std_logic_vector(119, 8),
61824 => conv_std_logic_vector(120, 8),
61825 => conv_std_logic_vector(121, 8),
61826 => conv_std_logic_vector(122, 8),
61827 => conv_std_logic_vector(123, 8),
61828 => conv_std_logic_vector(124, 8),
61829 => conv_std_logic_vector(125, 8),
61830 => conv_std_logic_vector(126, 8),
61831 => conv_std_logic_vector(127, 8),
61832 => conv_std_logic_vector(128, 8),
61833 => conv_std_logic_vector(128, 8),
61834 => conv_std_logic_vector(129, 8),
61835 => conv_std_logic_vector(130, 8),
61836 => conv_std_logic_vector(131, 8),
61837 => conv_std_logic_vector(132, 8),
61838 => conv_std_logic_vector(133, 8),
61839 => conv_std_logic_vector(134, 8),
61840 => conv_std_logic_vector(135, 8),
61841 => conv_std_logic_vector(136, 8),
61842 => conv_std_logic_vector(137, 8),
61843 => conv_std_logic_vector(138, 8),
61844 => conv_std_logic_vector(139, 8),
61845 => conv_std_logic_vector(140, 8),
61846 => conv_std_logic_vector(141, 8),
61847 => conv_std_logic_vector(142, 8),
61848 => conv_std_logic_vector(143, 8),
61849 => conv_std_logic_vector(144, 8),
61850 => conv_std_logic_vector(144, 8),
61851 => conv_std_logic_vector(145, 8),
61852 => conv_std_logic_vector(146, 8),
61853 => conv_std_logic_vector(147, 8),
61854 => conv_std_logic_vector(148, 8),
61855 => conv_std_logic_vector(149, 8),
61856 => conv_std_logic_vector(150, 8),
61857 => conv_std_logic_vector(151, 8),
61858 => conv_std_logic_vector(152, 8),
61859 => conv_std_logic_vector(153, 8),
61860 => conv_std_logic_vector(154, 8),
61861 => conv_std_logic_vector(155, 8),
61862 => conv_std_logic_vector(156, 8),
61863 => conv_std_logic_vector(157, 8),
61864 => conv_std_logic_vector(158, 8),
61865 => conv_std_logic_vector(159, 8),
61866 => conv_std_logic_vector(160, 8),
61867 => conv_std_logic_vector(160, 8),
61868 => conv_std_logic_vector(161, 8),
61869 => conv_std_logic_vector(162, 8),
61870 => conv_std_logic_vector(163, 8),
61871 => conv_std_logic_vector(164, 8),
61872 => conv_std_logic_vector(165, 8),
61873 => conv_std_logic_vector(166, 8),
61874 => conv_std_logic_vector(167, 8),
61875 => conv_std_logic_vector(168, 8),
61876 => conv_std_logic_vector(169, 8),
61877 => conv_std_logic_vector(170, 8),
61878 => conv_std_logic_vector(171, 8),
61879 => conv_std_logic_vector(172, 8),
61880 => conv_std_logic_vector(173, 8),
61881 => conv_std_logic_vector(174, 8),
61882 => conv_std_logic_vector(175, 8),
61883 => conv_std_logic_vector(176, 8),
61884 => conv_std_logic_vector(176, 8),
61885 => conv_std_logic_vector(177, 8),
61886 => conv_std_logic_vector(178, 8),
61887 => conv_std_logic_vector(179, 8),
61888 => conv_std_logic_vector(180, 8),
61889 => conv_std_logic_vector(181, 8),
61890 => conv_std_logic_vector(182, 8),
61891 => conv_std_logic_vector(183, 8),
61892 => conv_std_logic_vector(184, 8),
61893 => conv_std_logic_vector(185, 8),
61894 => conv_std_logic_vector(186, 8),
61895 => conv_std_logic_vector(187, 8),
61896 => conv_std_logic_vector(188, 8),
61897 => conv_std_logic_vector(189, 8),
61898 => conv_std_logic_vector(190, 8),
61899 => conv_std_logic_vector(191, 8),
61900 => conv_std_logic_vector(192, 8),
61901 => conv_std_logic_vector(192, 8),
61902 => conv_std_logic_vector(193, 8),
61903 => conv_std_logic_vector(194, 8),
61904 => conv_std_logic_vector(195, 8),
61905 => conv_std_logic_vector(196, 8),
61906 => conv_std_logic_vector(197, 8),
61907 => conv_std_logic_vector(198, 8),
61908 => conv_std_logic_vector(199, 8),
61909 => conv_std_logic_vector(200, 8),
61910 => conv_std_logic_vector(201, 8),
61911 => conv_std_logic_vector(202, 8),
61912 => conv_std_logic_vector(203, 8),
61913 => conv_std_logic_vector(204, 8),
61914 => conv_std_logic_vector(205, 8),
61915 => conv_std_logic_vector(206, 8),
61916 => conv_std_logic_vector(207, 8),
61917 => conv_std_logic_vector(208, 8),
61918 => conv_std_logic_vector(208, 8),
61919 => conv_std_logic_vector(209, 8),
61920 => conv_std_logic_vector(210, 8),
61921 => conv_std_logic_vector(211, 8),
61922 => conv_std_logic_vector(212, 8),
61923 => conv_std_logic_vector(213, 8),
61924 => conv_std_logic_vector(214, 8),
61925 => conv_std_logic_vector(215, 8),
61926 => conv_std_logic_vector(216, 8),
61927 => conv_std_logic_vector(217, 8),
61928 => conv_std_logic_vector(218, 8),
61929 => conv_std_logic_vector(219, 8),
61930 => conv_std_logic_vector(220, 8),
61931 => conv_std_logic_vector(221, 8),
61932 => conv_std_logic_vector(222, 8),
61933 => conv_std_logic_vector(223, 8),
61934 => conv_std_logic_vector(224, 8),
61935 => conv_std_logic_vector(224, 8),
61936 => conv_std_logic_vector(225, 8),
61937 => conv_std_logic_vector(226, 8),
61938 => conv_std_logic_vector(227, 8),
61939 => conv_std_logic_vector(228, 8),
61940 => conv_std_logic_vector(229, 8),
61941 => conv_std_logic_vector(230, 8),
61942 => conv_std_logic_vector(231, 8),
61943 => conv_std_logic_vector(232, 8),
61944 => conv_std_logic_vector(233, 8),
61945 => conv_std_logic_vector(234, 8),
61946 => conv_std_logic_vector(235, 8),
61947 => conv_std_logic_vector(236, 8),
61948 => conv_std_logic_vector(237, 8),
61949 => conv_std_logic_vector(238, 8),
61950 => conv_std_logic_vector(239, 8),
61951 => conv_std_logic_vector(240, 8),
61952 => conv_std_logic_vector(0, 8),
61953 => conv_std_logic_vector(0, 8),
61954 => conv_std_logic_vector(1, 8),
61955 => conv_std_logic_vector(2, 8),
61956 => conv_std_logic_vector(3, 8),
61957 => conv_std_logic_vector(4, 8),
61958 => conv_std_logic_vector(5, 8),
61959 => conv_std_logic_vector(6, 8),
61960 => conv_std_logic_vector(7, 8),
61961 => conv_std_logic_vector(8, 8),
61962 => conv_std_logic_vector(9, 8),
61963 => conv_std_logic_vector(10, 8),
61964 => conv_std_logic_vector(11, 8),
61965 => conv_std_logic_vector(12, 8),
61966 => conv_std_logic_vector(13, 8),
61967 => conv_std_logic_vector(14, 8),
61968 => conv_std_logic_vector(15, 8),
61969 => conv_std_logic_vector(16, 8),
61970 => conv_std_logic_vector(17, 8),
61971 => conv_std_logic_vector(17, 8),
61972 => conv_std_logic_vector(18, 8),
61973 => conv_std_logic_vector(19, 8),
61974 => conv_std_logic_vector(20, 8),
61975 => conv_std_logic_vector(21, 8),
61976 => conv_std_logic_vector(22, 8),
61977 => conv_std_logic_vector(23, 8),
61978 => conv_std_logic_vector(24, 8),
61979 => conv_std_logic_vector(25, 8),
61980 => conv_std_logic_vector(26, 8),
61981 => conv_std_logic_vector(27, 8),
61982 => conv_std_logic_vector(28, 8),
61983 => conv_std_logic_vector(29, 8),
61984 => conv_std_logic_vector(30, 8),
61985 => conv_std_logic_vector(31, 8),
61986 => conv_std_logic_vector(32, 8),
61987 => conv_std_logic_vector(33, 8),
61988 => conv_std_logic_vector(34, 8),
61989 => conv_std_logic_vector(34, 8),
61990 => conv_std_logic_vector(35, 8),
61991 => conv_std_logic_vector(36, 8),
61992 => conv_std_logic_vector(37, 8),
61993 => conv_std_logic_vector(38, 8),
61994 => conv_std_logic_vector(39, 8),
61995 => conv_std_logic_vector(40, 8),
61996 => conv_std_logic_vector(41, 8),
61997 => conv_std_logic_vector(42, 8),
61998 => conv_std_logic_vector(43, 8),
61999 => conv_std_logic_vector(44, 8),
62000 => conv_std_logic_vector(45, 8),
62001 => conv_std_logic_vector(46, 8),
62002 => conv_std_logic_vector(47, 8),
62003 => conv_std_logic_vector(48, 8),
62004 => conv_std_logic_vector(49, 8),
62005 => conv_std_logic_vector(50, 8),
62006 => conv_std_logic_vector(51, 8),
62007 => conv_std_logic_vector(51, 8),
62008 => conv_std_logic_vector(52, 8),
62009 => conv_std_logic_vector(53, 8),
62010 => conv_std_logic_vector(54, 8),
62011 => conv_std_logic_vector(55, 8),
62012 => conv_std_logic_vector(56, 8),
62013 => conv_std_logic_vector(57, 8),
62014 => conv_std_logic_vector(58, 8),
62015 => conv_std_logic_vector(59, 8),
62016 => conv_std_logic_vector(60, 8),
62017 => conv_std_logic_vector(61, 8),
62018 => conv_std_logic_vector(62, 8),
62019 => conv_std_logic_vector(63, 8),
62020 => conv_std_logic_vector(64, 8),
62021 => conv_std_logic_vector(65, 8),
62022 => conv_std_logic_vector(66, 8),
62023 => conv_std_logic_vector(67, 8),
62024 => conv_std_logic_vector(68, 8),
62025 => conv_std_logic_vector(69, 8),
62026 => conv_std_logic_vector(69, 8),
62027 => conv_std_logic_vector(70, 8),
62028 => conv_std_logic_vector(71, 8),
62029 => conv_std_logic_vector(72, 8),
62030 => conv_std_logic_vector(73, 8),
62031 => conv_std_logic_vector(74, 8),
62032 => conv_std_logic_vector(75, 8),
62033 => conv_std_logic_vector(76, 8),
62034 => conv_std_logic_vector(77, 8),
62035 => conv_std_logic_vector(78, 8),
62036 => conv_std_logic_vector(79, 8),
62037 => conv_std_logic_vector(80, 8),
62038 => conv_std_logic_vector(81, 8),
62039 => conv_std_logic_vector(82, 8),
62040 => conv_std_logic_vector(83, 8),
62041 => conv_std_logic_vector(84, 8),
62042 => conv_std_logic_vector(85, 8),
62043 => conv_std_logic_vector(86, 8),
62044 => conv_std_logic_vector(86, 8),
62045 => conv_std_logic_vector(87, 8),
62046 => conv_std_logic_vector(88, 8),
62047 => conv_std_logic_vector(89, 8),
62048 => conv_std_logic_vector(90, 8),
62049 => conv_std_logic_vector(91, 8),
62050 => conv_std_logic_vector(92, 8),
62051 => conv_std_logic_vector(93, 8),
62052 => conv_std_logic_vector(94, 8),
62053 => conv_std_logic_vector(95, 8),
62054 => conv_std_logic_vector(96, 8),
62055 => conv_std_logic_vector(97, 8),
62056 => conv_std_logic_vector(98, 8),
62057 => conv_std_logic_vector(99, 8),
62058 => conv_std_logic_vector(100, 8),
62059 => conv_std_logic_vector(101, 8),
62060 => conv_std_logic_vector(102, 8),
62061 => conv_std_logic_vector(103, 8),
62062 => conv_std_logic_vector(103, 8),
62063 => conv_std_logic_vector(104, 8),
62064 => conv_std_logic_vector(105, 8),
62065 => conv_std_logic_vector(106, 8),
62066 => conv_std_logic_vector(107, 8),
62067 => conv_std_logic_vector(108, 8),
62068 => conv_std_logic_vector(109, 8),
62069 => conv_std_logic_vector(110, 8),
62070 => conv_std_logic_vector(111, 8),
62071 => conv_std_logic_vector(112, 8),
62072 => conv_std_logic_vector(113, 8),
62073 => conv_std_logic_vector(114, 8),
62074 => conv_std_logic_vector(115, 8),
62075 => conv_std_logic_vector(116, 8),
62076 => conv_std_logic_vector(117, 8),
62077 => conv_std_logic_vector(118, 8),
62078 => conv_std_logic_vector(119, 8),
62079 => conv_std_logic_vector(120, 8),
62080 => conv_std_logic_vector(121, 8),
62081 => conv_std_logic_vector(121, 8),
62082 => conv_std_logic_vector(122, 8),
62083 => conv_std_logic_vector(123, 8),
62084 => conv_std_logic_vector(124, 8),
62085 => conv_std_logic_vector(125, 8),
62086 => conv_std_logic_vector(126, 8),
62087 => conv_std_logic_vector(127, 8),
62088 => conv_std_logic_vector(128, 8),
62089 => conv_std_logic_vector(129, 8),
62090 => conv_std_logic_vector(130, 8),
62091 => conv_std_logic_vector(131, 8),
62092 => conv_std_logic_vector(132, 8),
62093 => conv_std_logic_vector(133, 8),
62094 => conv_std_logic_vector(134, 8),
62095 => conv_std_logic_vector(135, 8),
62096 => conv_std_logic_vector(136, 8),
62097 => conv_std_logic_vector(137, 8),
62098 => conv_std_logic_vector(138, 8),
62099 => conv_std_logic_vector(138, 8),
62100 => conv_std_logic_vector(139, 8),
62101 => conv_std_logic_vector(140, 8),
62102 => conv_std_logic_vector(141, 8),
62103 => conv_std_logic_vector(142, 8),
62104 => conv_std_logic_vector(143, 8),
62105 => conv_std_logic_vector(144, 8),
62106 => conv_std_logic_vector(145, 8),
62107 => conv_std_logic_vector(146, 8),
62108 => conv_std_logic_vector(147, 8),
62109 => conv_std_logic_vector(148, 8),
62110 => conv_std_logic_vector(149, 8),
62111 => conv_std_logic_vector(150, 8),
62112 => conv_std_logic_vector(151, 8),
62113 => conv_std_logic_vector(152, 8),
62114 => conv_std_logic_vector(153, 8),
62115 => conv_std_logic_vector(154, 8),
62116 => conv_std_logic_vector(155, 8),
62117 => conv_std_logic_vector(155, 8),
62118 => conv_std_logic_vector(156, 8),
62119 => conv_std_logic_vector(157, 8),
62120 => conv_std_logic_vector(158, 8),
62121 => conv_std_logic_vector(159, 8),
62122 => conv_std_logic_vector(160, 8),
62123 => conv_std_logic_vector(161, 8),
62124 => conv_std_logic_vector(162, 8),
62125 => conv_std_logic_vector(163, 8),
62126 => conv_std_logic_vector(164, 8),
62127 => conv_std_logic_vector(165, 8),
62128 => conv_std_logic_vector(166, 8),
62129 => conv_std_logic_vector(167, 8),
62130 => conv_std_logic_vector(168, 8),
62131 => conv_std_logic_vector(169, 8),
62132 => conv_std_logic_vector(170, 8),
62133 => conv_std_logic_vector(171, 8),
62134 => conv_std_logic_vector(172, 8),
62135 => conv_std_logic_vector(172, 8),
62136 => conv_std_logic_vector(173, 8),
62137 => conv_std_logic_vector(174, 8),
62138 => conv_std_logic_vector(175, 8),
62139 => conv_std_logic_vector(176, 8),
62140 => conv_std_logic_vector(177, 8),
62141 => conv_std_logic_vector(178, 8),
62142 => conv_std_logic_vector(179, 8),
62143 => conv_std_logic_vector(180, 8),
62144 => conv_std_logic_vector(181, 8),
62145 => conv_std_logic_vector(182, 8),
62146 => conv_std_logic_vector(183, 8),
62147 => conv_std_logic_vector(184, 8),
62148 => conv_std_logic_vector(185, 8),
62149 => conv_std_logic_vector(186, 8),
62150 => conv_std_logic_vector(187, 8),
62151 => conv_std_logic_vector(188, 8),
62152 => conv_std_logic_vector(189, 8),
62153 => conv_std_logic_vector(190, 8),
62154 => conv_std_logic_vector(190, 8),
62155 => conv_std_logic_vector(191, 8),
62156 => conv_std_logic_vector(192, 8),
62157 => conv_std_logic_vector(193, 8),
62158 => conv_std_logic_vector(194, 8),
62159 => conv_std_logic_vector(195, 8),
62160 => conv_std_logic_vector(196, 8),
62161 => conv_std_logic_vector(197, 8),
62162 => conv_std_logic_vector(198, 8),
62163 => conv_std_logic_vector(199, 8),
62164 => conv_std_logic_vector(200, 8),
62165 => conv_std_logic_vector(201, 8),
62166 => conv_std_logic_vector(202, 8),
62167 => conv_std_logic_vector(203, 8),
62168 => conv_std_logic_vector(204, 8),
62169 => conv_std_logic_vector(205, 8),
62170 => conv_std_logic_vector(206, 8),
62171 => conv_std_logic_vector(207, 8),
62172 => conv_std_logic_vector(207, 8),
62173 => conv_std_logic_vector(208, 8),
62174 => conv_std_logic_vector(209, 8),
62175 => conv_std_logic_vector(210, 8),
62176 => conv_std_logic_vector(211, 8),
62177 => conv_std_logic_vector(212, 8),
62178 => conv_std_logic_vector(213, 8),
62179 => conv_std_logic_vector(214, 8),
62180 => conv_std_logic_vector(215, 8),
62181 => conv_std_logic_vector(216, 8),
62182 => conv_std_logic_vector(217, 8),
62183 => conv_std_logic_vector(218, 8),
62184 => conv_std_logic_vector(219, 8),
62185 => conv_std_logic_vector(220, 8),
62186 => conv_std_logic_vector(221, 8),
62187 => conv_std_logic_vector(222, 8),
62188 => conv_std_logic_vector(223, 8),
62189 => conv_std_logic_vector(224, 8),
62190 => conv_std_logic_vector(224, 8),
62191 => conv_std_logic_vector(225, 8),
62192 => conv_std_logic_vector(226, 8),
62193 => conv_std_logic_vector(227, 8),
62194 => conv_std_logic_vector(228, 8),
62195 => conv_std_logic_vector(229, 8),
62196 => conv_std_logic_vector(230, 8),
62197 => conv_std_logic_vector(231, 8),
62198 => conv_std_logic_vector(232, 8),
62199 => conv_std_logic_vector(233, 8),
62200 => conv_std_logic_vector(234, 8),
62201 => conv_std_logic_vector(235, 8),
62202 => conv_std_logic_vector(236, 8),
62203 => conv_std_logic_vector(237, 8),
62204 => conv_std_logic_vector(238, 8),
62205 => conv_std_logic_vector(239, 8),
62206 => conv_std_logic_vector(240, 8),
62207 => conv_std_logic_vector(241, 8),
62208 => conv_std_logic_vector(0, 8),
62209 => conv_std_logic_vector(0, 8),
62210 => conv_std_logic_vector(1, 8),
62211 => conv_std_logic_vector(2, 8),
62212 => conv_std_logic_vector(3, 8),
62213 => conv_std_logic_vector(4, 8),
62214 => conv_std_logic_vector(5, 8),
62215 => conv_std_logic_vector(6, 8),
62216 => conv_std_logic_vector(7, 8),
62217 => conv_std_logic_vector(8, 8),
62218 => conv_std_logic_vector(9, 8),
62219 => conv_std_logic_vector(10, 8),
62220 => conv_std_logic_vector(11, 8),
62221 => conv_std_logic_vector(12, 8),
62222 => conv_std_logic_vector(13, 8),
62223 => conv_std_logic_vector(14, 8),
62224 => conv_std_logic_vector(15, 8),
62225 => conv_std_logic_vector(16, 8),
62226 => conv_std_logic_vector(17, 8),
62227 => conv_std_logic_vector(18, 8),
62228 => conv_std_logic_vector(18, 8),
62229 => conv_std_logic_vector(19, 8),
62230 => conv_std_logic_vector(20, 8),
62231 => conv_std_logic_vector(21, 8),
62232 => conv_std_logic_vector(22, 8),
62233 => conv_std_logic_vector(23, 8),
62234 => conv_std_logic_vector(24, 8),
62235 => conv_std_logic_vector(25, 8),
62236 => conv_std_logic_vector(26, 8),
62237 => conv_std_logic_vector(27, 8),
62238 => conv_std_logic_vector(28, 8),
62239 => conv_std_logic_vector(29, 8),
62240 => conv_std_logic_vector(30, 8),
62241 => conv_std_logic_vector(31, 8),
62242 => conv_std_logic_vector(32, 8),
62243 => conv_std_logic_vector(33, 8),
62244 => conv_std_logic_vector(34, 8),
62245 => conv_std_logic_vector(35, 8),
62246 => conv_std_logic_vector(36, 8),
62247 => conv_std_logic_vector(37, 8),
62248 => conv_std_logic_vector(37, 8),
62249 => conv_std_logic_vector(38, 8),
62250 => conv_std_logic_vector(39, 8),
62251 => conv_std_logic_vector(40, 8),
62252 => conv_std_logic_vector(41, 8),
62253 => conv_std_logic_vector(42, 8),
62254 => conv_std_logic_vector(43, 8),
62255 => conv_std_logic_vector(44, 8),
62256 => conv_std_logic_vector(45, 8),
62257 => conv_std_logic_vector(46, 8),
62258 => conv_std_logic_vector(47, 8),
62259 => conv_std_logic_vector(48, 8),
62260 => conv_std_logic_vector(49, 8),
62261 => conv_std_logic_vector(50, 8),
62262 => conv_std_logic_vector(51, 8),
62263 => conv_std_logic_vector(52, 8),
62264 => conv_std_logic_vector(53, 8),
62265 => conv_std_logic_vector(54, 8),
62266 => conv_std_logic_vector(55, 8),
62267 => conv_std_logic_vector(56, 8),
62268 => conv_std_logic_vector(56, 8),
62269 => conv_std_logic_vector(57, 8),
62270 => conv_std_logic_vector(58, 8),
62271 => conv_std_logic_vector(59, 8),
62272 => conv_std_logic_vector(60, 8),
62273 => conv_std_logic_vector(61, 8),
62274 => conv_std_logic_vector(62, 8),
62275 => conv_std_logic_vector(63, 8),
62276 => conv_std_logic_vector(64, 8),
62277 => conv_std_logic_vector(65, 8),
62278 => conv_std_logic_vector(66, 8),
62279 => conv_std_logic_vector(67, 8),
62280 => conv_std_logic_vector(68, 8),
62281 => conv_std_logic_vector(69, 8),
62282 => conv_std_logic_vector(70, 8),
62283 => conv_std_logic_vector(71, 8),
62284 => conv_std_logic_vector(72, 8),
62285 => conv_std_logic_vector(73, 8),
62286 => conv_std_logic_vector(74, 8),
62287 => conv_std_logic_vector(74, 8),
62288 => conv_std_logic_vector(75, 8),
62289 => conv_std_logic_vector(76, 8),
62290 => conv_std_logic_vector(77, 8),
62291 => conv_std_logic_vector(78, 8),
62292 => conv_std_logic_vector(79, 8),
62293 => conv_std_logic_vector(80, 8),
62294 => conv_std_logic_vector(81, 8),
62295 => conv_std_logic_vector(82, 8),
62296 => conv_std_logic_vector(83, 8),
62297 => conv_std_logic_vector(84, 8),
62298 => conv_std_logic_vector(85, 8),
62299 => conv_std_logic_vector(86, 8),
62300 => conv_std_logic_vector(87, 8),
62301 => conv_std_logic_vector(88, 8),
62302 => conv_std_logic_vector(89, 8),
62303 => conv_std_logic_vector(90, 8),
62304 => conv_std_logic_vector(91, 8),
62305 => conv_std_logic_vector(92, 8),
62306 => conv_std_logic_vector(93, 8),
62307 => conv_std_logic_vector(93, 8),
62308 => conv_std_logic_vector(94, 8),
62309 => conv_std_logic_vector(95, 8),
62310 => conv_std_logic_vector(96, 8),
62311 => conv_std_logic_vector(97, 8),
62312 => conv_std_logic_vector(98, 8),
62313 => conv_std_logic_vector(99, 8),
62314 => conv_std_logic_vector(100, 8),
62315 => conv_std_logic_vector(101, 8),
62316 => conv_std_logic_vector(102, 8),
62317 => conv_std_logic_vector(103, 8),
62318 => conv_std_logic_vector(104, 8),
62319 => conv_std_logic_vector(105, 8),
62320 => conv_std_logic_vector(106, 8),
62321 => conv_std_logic_vector(107, 8),
62322 => conv_std_logic_vector(108, 8),
62323 => conv_std_logic_vector(109, 8),
62324 => conv_std_logic_vector(110, 8),
62325 => conv_std_logic_vector(111, 8),
62326 => conv_std_logic_vector(112, 8),
62327 => conv_std_logic_vector(112, 8),
62328 => conv_std_logic_vector(113, 8),
62329 => conv_std_logic_vector(114, 8),
62330 => conv_std_logic_vector(115, 8),
62331 => conv_std_logic_vector(116, 8),
62332 => conv_std_logic_vector(117, 8),
62333 => conv_std_logic_vector(118, 8),
62334 => conv_std_logic_vector(119, 8),
62335 => conv_std_logic_vector(120, 8),
62336 => conv_std_logic_vector(121, 8),
62337 => conv_std_logic_vector(122, 8),
62338 => conv_std_logic_vector(123, 8),
62339 => conv_std_logic_vector(124, 8),
62340 => conv_std_logic_vector(125, 8),
62341 => conv_std_logic_vector(126, 8),
62342 => conv_std_logic_vector(127, 8),
62343 => conv_std_logic_vector(128, 8),
62344 => conv_std_logic_vector(129, 8),
62345 => conv_std_logic_vector(130, 8),
62346 => conv_std_logic_vector(130, 8),
62347 => conv_std_logic_vector(131, 8),
62348 => conv_std_logic_vector(132, 8),
62349 => conv_std_logic_vector(133, 8),
62350 => conv_std_logic_vector(134, 8),
62351 => conv_std_logic_vector(135, 8),
62352 => conv_std_logic_vector(136, 8),
62353 => conv_std_logic_vector(137, 8),
62354 => conv_std_logic_vector(138, 8),
62355 => conv_std_logic_vector(139, 8),
62356 => conv_std_logic_vector(140, 8),
62357 => conv_std_logic_vector(141, 8),
62358 => conv_std_logic_vector(142, 8),
62359 => conv_std_logic_vector(143, 8),
62360 => conv_std_logic_vector(144, 8),
62361 => conv_std_logic_vector(145, 8),
62362 => conv_std_logic_vector(146, 8),
62363 => conv_std_logic_vector(147, 8),
62364 => conv_std_logic_vector(148, 8),
62365 => conv_std_logic_vector(149, 8),
62366 => conv_std_logic_vector(149, 8),
62367 => conv_std_logic_vector(150, 8),
62368 => conv_std_logic_vector(151, 8),
62369 => conv_std_logic_vector(152, 8),
62370 => conv_std_logic_vector(153, 8),
62371 => conv_std_logic_vector(154, 8),
62372 => conv_std_logic_vector(155, 8),
62373 => conv_std_logic_vector(156, 8),
62374 => conv_std_logic_vector(157, 8),
62375 => conv_std_logic_vector(158, 8),
62376 => conv_std_logic_vector(159, 8),
62377 => conv_std_logic_vector(160, 8),
62378 => conv_std_logic_vector(161, 8),
62379 => conv_std_logic_vector(162, 8),
62380 => conv_std_logic_vector(163, 8),
62381 => conv_std_logic_vector(164, 8),
62382 => conv_std_logic_vector(165, 8),
62383 => conv_std_logic_vector(166, 8),
62384 => conv_std_logic_vector(167, 8),
62385 => conv_std_logic_vector(168, 8),
62386 => conv_std_logic_vector(168, 8),
62387 => conv_std_logic_vector(169, 8),
62388 => conv_std_logic_vector(170, 8),
62389 => conv_std_logic_vector(171, 8),
62390 => conv_std_logic_vector(172, 8),
62391 => conv_std_logic_vector(173, 8),
62392 => conv_std_logic_vector(174, 8),
62393 => conv_std_logic_vector(175, 8),
62394 => conv_std_logic_vector(176, 8),
62395 => conv_std_logic_vector(177, 8),
62396 => conv_std_logic_vector(178, 8),
62397 => conv_std_logic_vector(179, 8),
62398 => conv_std_logic_vector(180, 8),
62399 => conv_std_logic_vector(181, 8),
62400 => conv_std_logic_vector(182, 8),
62401 => conv_std_logic_vector(183, 8),
62402 => conv_std_logic_vector(184, 8),
62403 => conv_std_logic_vector(185, 8),
62404 => conv_std_logic_vector(186, 8),
62405 => conv_std_logic_vector(186, 8),
62406 => conv_std_logic_vector(187, 8),
62407 => conv_std_logic_vector(188, 8),
62408 => conv_std_logic_vector(189, 8),
62409 => conv_std_logic_vector(190, 8),
62410 => conv_std_logic_vector(191, 8),
62411 => conv_std_logic_vector(192, 8),
62412 => conv_std_logic_vector(193, 8),
62413 => conv_std_logic_vector(194, 8),
62414 => conv_std_logic_vector(195, 8),
62415 => conv_std_logic_vector(196, 8),
62416 => conv_std_logic_vector(197, 8),
62417 => conv_std_logic_vector(198, 8),
62418 => conv_std_logic_vector(199, 8),
62419 => conv_std_logic_vector(200, 8),
62420 => conv_std_logic_vector(201, 8),
62421 => conv_std_logic_vector(202, 8),
62422 => conv_std_logic_vector(203, 8),
62423 => conv_std_logic_vector(204, 8),
62424 => conv_std_logic_vector(205, 8),
62425 => conv_std_logic_vector(205, 8),
62426 => conv_std_logic_vector(206, 8),
62427 => conv_std_logic_vector(207, 8),
62428 => conv_std_logic_vector(208, 8),
62429 => conv_std_logic_vector(209, 8),
62430 => conv_std_logic_vector(210, 8),
62431 => conv_std_logic_vector(211, 8),
62432 => conv_std_logic_vector(212, 8),
62433 => conv_std_logic_vector(213, 8),
62434 => conv_std_logic_vector(214, 8),
62435 => conv_std_logic_vector(215, 8),
62436 => conv_std_logic_vector(216, 8),
62437 => conv_std_logic_vector(217, 8),
62438 => conv_std_logic_vector(218, 8),
62439 => conv_std_logic_vector(219, 8),
62440 => conv_std_logic_vector(220, 8),
62441 => conv_std_logic_vector(221, 8),
62442 => conv_std_logic_vector(222, 8),
62443 => conv_std_logic_vector(223, 8),
62444 => conv_std_logic_vector(224, 8),
62445 => conv_std_logic_vector(224, 8),
62446 => conv_std_logic_vector(225, 8),
62447 => conv_std_logic_vector(226, 8),
62448 => conv_std_logic_vector(227, 8),
62449 => conv_std_logic_vector(228, 8),
62450 => conv_std_logic_vector(229, 8),
62451 => conv_std_logic_vector(230, 8),
62452 => conv_std_logic_vector(231, 8),
62453 => conv_std_logic_vector(232, 8),
62454 => conv_std_logic_vector(233, 8),
62455 => conv_std_logic_vector(234, 8),
62456 => conv_std_logic_vector(235, 8),
62457 => conv_std_logic_vector(236, 8),
62458 => conv_std_logic_vector(237, 8),
62459 => conv_std_logic_vector(238, 8),
62460 => conv_std_logic_vector(239, 8),
62461 => conv_std_logic_vector(240, 8),
62462 => conv_std_logic_vector(241, 8),
62463 => conv_std_logic_vector(242, 8),
62464 => conv_std_logic_vector(0, 8),
62465 => conv_std_logic_vector(0, 8),
62466 => conv_std_logic_vector(1, 8),
62467 => conv_std_logic_vector(2, 8),
62468 => conv_std_logic_vector(3, 8),
62469 => conv_std_logic_vector(4, 8),
62470 => conv_std_logic_vector(5, 8),
62471 => conv_std_logic_vector(6, 8),
62472 => conv_std_logic_vector(7, 8),
62473 => conv_std_logic_vector(8, 8),
62474 => conv_std_logic_vector(9, 8),
62475 => conv_std_logic_vector(10, 8),
62476 => conv_std_logic_vector(11, 8),
62477 => conv_std_logic_vector(12, 8),
62478 => conv_std_logic_vector(13, 8),
62479 => conv_std_logic_vector(14, 8),
62480 => conv_std_logic_vector(15, 8),
62481 => conv_std_logic_vector(16, 8),
62482 => conv_std_logic_vector(17, 8),
62483 => conv_std_logic_vector(18, 8),
62484 => conv_std_logic_vector(19, 8),
62485 => conv_std_logic_vector(20, 8),
62486 => conv_std_logic_vector(20, 8),
62487 => conv_std_logic_vector(21, 8),
62488 => conv_std_logic_vector(22, 8),
62489 => conv_std_logic_vector(23, 8),
62490 => conv_std_logic_vector(24, 8),
62491 => conv_std_logic_vector(25, 8),
62492 => conv_std_logic_vector(26, 8),
62493 => conv_std_logic_vector(27, 8),
62494 => conv_std_logic_vector(28, 8),
62495 => conv_std_logic_vector(29, 8),
62496 => conv_std_logic_vector(30, 8),
62497 => conv_std_logic_vector(31, 8),
62498 => conv_std_logic_vector(32, 8),
62499 => conv_std_logic_vector(33, 8),
62500 => conv_std_logic_vector(34, 8),
62501 => conv_std_logic_vector(35, 8),
62502 => conv_std_logic_vector(36, 8),
62503 => conv_std_logic_vector(37, 8),
62504 => conv_std_logic_vector(38, 8),
62505 => conv_std_logic_vector(39, 8),
62506 => conv_std_logic_vector(40, 8),
62507 => conv_std_logic_vector(40, 8),
62508 => conv_std_logic_vector(41, 8),
62509 => conv_std_logic_vector(42, 8),
62510 => conv_std_logic_vector(43, 8),
62511 => conv_std_logic_vector(44, 8),
62512 => conv_std_logic_vector(45, 8),
62513 => conv_std_logic_vector(46, 8),
62514 => conv_std_logic_vector(47, 8),
62515 => conv_std_logic_vector(48, 8),
62516 => conv_std_logic_vector(49, 8),
62517 => conv_std_logic_vector(50, 8),
62518 => conv_std_logic_vector(51, 8),
62519 => conv_std_logic_vector(52, 8),
62520 => conv_std_logic_vector(53, 8),
62521 => conv_std_logic_vector(54, 8),
62522 => conv_std_logic_vector(55, 8),
62523 => conv_std_logic_vector(56, 8),
62524 => conv_std_logic_vector(57, 8),
62525 => conv_std_logic_vector(58, 8),
62526 => conv_std_logic_vector(59, 8),
62527 => conv_std_logic_vector(60, 8),
62528 => conv_std_logic_vector(61, 8),
62529 => conv_std_logic_vector(61, 8),
62530 => conv_std_logic_vector(62, 8),
62531 => conv_std_logic_vector(63, 8),
62532 => conv_std_logic_vector(64, 8),
62533 => conv_std_logic_vector(65, 8),
62534 => conv_std_logic_vector(66, 8),
62535 => conv_std_logic_vector(67, 8),
62536 => conv_std_logic_vector(68, 8),
62537 => conv_std_logic_vector(69, 8),
62538 => conv_std_logic_vector(70, 8),
62539 => conv_std_logic_vector(71, 8),
62540 => conv_std_logic_vector(72, 8),
62541 => conv_std_logic_vector(73, 8),
62542 => conv_std_logic_vector(74, 8),
62543 => conv_std_logic_vector(75, 8),
62544 => conv_std_logic_vector(76, 8),
62545 => conv_std_logic_vector(77, 8),
62546 => conv_std_logic_vector(78, 8),
62547 => conv_std_logic_vector(79, 8),
62548 => conv_std_logic_vector(80, 8),
62549 => conv_std_logic_vector(81, 8),
62550 => conv_std_logic_vector(81, 8),
62551 => conv_std_logic_vector(82, 8),
62552 => conv_std_logic_vector(83, 8),
62553 => conv_std_logic_vector(84, 8),
62554 => conv_std_logic_vector(85, 8),
62555 => conv_std_logic_vector(86, 8),
62556 => conv_std_logic_vector(87, 8),
62557 => conv_std_logic_vector(88, 8),
62558 => conv_std_logic_vector(89, 8),
62559 => conv_std_logic_vector(90, 8),
62560 => conv_std_logic_vector(91, 8),
62561 => conv_std_logic_vector(92, 8),
62562 => conv_std_logic_vector(93, 8),
62563 => conv_std_logic_vector(94, 8),
62564 => conv_std_logic_vector(95, 8),
62565 => conv_std_logic_vector(96, 8),
62566 => conv_std_logic_vector(97, 8),
62567 => conv_std_logic_vector(98, 8),
62568 => conv_std_logic_vector(99, 8),
62569 => conv_std_logic_vector(100, 8),
62570 => conv_std_logic_vector(101, 8),
62571 => conv_std_logic_vector(101, 8),
62572 => conv_std_logic_vector(102, 8),
62573 => conv_std_logic_vector(103, 8),
62574 => conv_std_logic_vector(104, 8),
62575 => conv_std_logic_vector(105, 8),
62576 => conv_std_logic_vector(106, 8),
62577 => conv_std_logic_vector(107, 8),
62578 => conv_std_logic_vector(108, 8),
62579 => conv_std_logic_vector(109, 8),
62580 => conv_std_logic_vector(110, 8),
62581 => conv_std_logic_vector(111, 8),
62582 => conv_std_logic_vector(112, 8),
62583 => conv_std_logic_vector(113, 8),
62584 => conv_std_logic_vector(114, 8),
62585 => conv_std_logic_vector(115, 8),
62586 => conv_std_logic_vector(116, 8),
62587 => conv_std_logic_vector(117, 8),
62588 => conv_std_logic_vector(118, 8),
62589 => conv_std_logic_vector(119, 8),
62590 => conv_std_logic_vector(120, 8),
62591 => conv_std_logic_vector(121, 8),
62592 => conv_std_logic_vector(122, 8),
62593 => conv_std_logic_vector(122, 8),
62594 => conv_std_logic_vector(123, 8),
62595 => conv_std_logic_vector(124, 8),
62596 => conv_std_logic_vector(125, 8),
62597 => conv_std_logic_vector(126, 8),
62598 => conv_std_logic_vector(127, 8),
62599 => conv_std_logic_vector(128, 8),
62600 => conv_std_logic_vector(129, 8),
62601 => conv_std_logic_vector(130, 8),
62602 => conv_std_logic_vector(131, 8),
62603 => conv_std_logic_vector(132, 8),
62604 => conv_std_logic_vector(133, 8),
62605 => conv_std_logic_vector(134, 8),
62606 => conv_std_logic_vector(135, 8),
62607 => conv_std_logic_vector(136, 8),
62608 => conv_std_logic_vector(137, 8),
62609 => conv_std_logic_vector(138, 8),
62610 => conv_std_logic_vector(139, 8),
62611 => conv_std_logic_vector(140, 8),
62612 => conv_std_logic_vector(141, 8),
62613 => conv_std_logic_vector(142, 8),
62614 => conv_std_logic_vector(142, 8),
62615 => conv_std_logic_vector(143, 8),
62616 => conv_std_logic_vector(144, 8),
62617 => conv_std_logic_vector(145, 8),
62618 => conv_std_logic_vector(146, 8),
62619 => conv_std_logic_vector(147, 8),
62620 => conv_std_logic_vector(148, 8),
62621 => conv_std_logic_vector(149, 8),
62622 => conv_std_logic_vector(150, 8),
62623 => conv_std_logic_vector(151, 8),
62624 => conv_std_logic_vector(152, 8),
62625 => conv_std_logic_vector(153, 8),
62626 => conv_std_logic_vector(154, 8),
62627 => conv_std_logic_vector(155, 8),
62628 => conv_std_logic_vector(156, 8),
62629 => conv_std_logic_vector(157, 8),
62630 => conv_std_logic_vector(158, 8),
62631 => conv_std_logic_vector(159, 8),
62632 => conv_std_logic_vector(160, 8),
62633 => conv_std_logic_vector(161, 8),
62634 => conv_std_logic_vector(162, 8),
62635 => conv_std_logic_vector(162, 8),
62636 => conv_std_logic_vector(163, 8),
62637 => conv_std_logic_vector(164, 8),
62638 => conv_std_logic_vector(165, 8),
62639 => conv_std_logic_vector(166, 8),
62640 => conv_std_logic_vector(167, 8),
62641 => conv_std_logic_vector(168, 8),
62642 => conv_std_logic_vector(169, 8),
62643 => conv_std_logic_vector(170, 8),
62644 => conv_std_logic_vector(171, 8),
62645 => conv_std_logic_vector(172, 8),
62646 => conv_std_logic_vector(173, 8),
62647 => conv_std_logic_vector(174, 8),
62648 => conv_std_logic_vector(175, 8),
62649 => conv_std_logic_vector(176, 8),
62650 => conv_std_logic_vector(177, 8),
62651 => conv_std_logic_vector(178, 8),
62652 => conv_std_logic_vector(179, 8),
62653 => conv_std_logic_vector(180, 8),
62654 => conv_std_logic_vector(181, 8),
62655 => conv_std_logic_vector(182, 8),
62656 => conv_std_logic_vector(183, 8),
62657 => conv_std_logic_vector(183, 8),
62658 => conv_std_logic_vector(184, 8),
62659 => conv_std_logic_vector(185, 8),
62660 => conv_std_logic_vector(186, 8),
62661 => conv_std_logic_vector(187, 8),
62662 => conv_std_logic_vector(188, 8),
62663 => conv_std_logic_vector(189, 8),
62664 => conv_std_logic_vector(190, 8),
62665 => conv_std_logic_vector(191, 8),
62666 => conv_std_logic_vector(192, 8),
62667 => conv_std_logic_vector(193, 8),
62668 => conv_std_logic_vector(194, 8),
62669 => conv_std_logic_vector(195, 8),
62670 => conv_std_logic_vector(196, 8),
62671 => conv_std_logic_vector(197, 8),
62672 => conv_std_logic_vector(198, 8),
62673 => conv_std_logic_vector(199, 8),
62674 => conv_std_logic_vector(200, 8),
62675 => conv_std_logic_vector(201, 8),
62676 => conv_std_logic_vector(202, 8),
62677 => conv_std_logic_vector(203, 8),
62678 => conv_std_logic_vector(203, 8),
62679 => conv_std_logic_vector(204, 8),
62680 => conv_std_logic_vector(205, 8),
62681 => conv_std_logic_vector(206, 8),
62682 => conv_std_logic_vector(207, 8),
62683 => conv_std_logic_vector(208, 8),
62684 => conv_std_logic_vector(209, 8),
62685 => conv_std_logic_vector(210, 8),
62686 => conv_std_logic_vector(211, 8),
62687 => conv_std_logic_vector(212, 8),
62688 => conv_std_logic_vector(213, 8),
62689 => conv_std_logic_vector(214, 8),
62690 => conv_std_logic_vector(215, 8),
62691 => conv_std_logic_vector(216, 8),
62692 => conv_std_logic_vector(217, 8),
62693 => conv_std_logic_vector(218, 8),
62694 => conv_std_logic_vector(219, 8),
62695 => conv_std_logic_vector(220, 8),
62696 => conv_std_logic_vector(221, 8),
62697 => conv_std_logic_vector(222, 8),
62698 => conv_std_logic_vector(223, 8),
62699 => conv_std_logic_vector(223, 8),
62700 => conv_std_logic_vector(224, 8),
62701 => conv_std_logic_vector(225, 8),
62702 => conv_std_logic_vector(226, 8),
62703 => conv_std_logic_vector(227, 8),
62704 => conv_std_logic_vector(228, 8),
62705 => conv_std_logic_vector(229, 8),
62706 => conv_std_logic_vector(230, 8),
62707 => conv_std_logic_vector(231, 8),
62708 => conv_std_logic_vector(232, 8),
62709 => conv_std_logic_vector(233, 8),
62710 => conv_std_logic_vector(234, 8),
62711 => conv_std_logic_vector(235, 8),
62712 => conv_std_logic_vector(236, 8),
62713 => conv_std_logic_vector(237, 8),
62714 => conv_std_logic_vector(238, 8),
62715 => conv_std_logic_vector(239, 8),
62716 => conv_std_logic_vector(240, 8),
62717 => conv_std_logic_vector(241, 8),
62718 => conv_std_logic_vector(242, 8),
62719 => conv_std_logic_vector(243, 8),
62720 => conv_std_logic_vector(0, 8),
62721 => conv_std_logic_vector(0, 8),
62722 => conv_std_logic_vector(1, 8),
62723 => conv_std_logic_vector(2, 8),
62724 => conv_std_logic_vector(3, 8),
62725 => conv_std_logic_vector(4, 8),
62726 => conv_std_logic_vector(5, 8),
62727 => conv_std_logic_vector(6, 8),
62728 => conv_std_logic_vector(7, 8),
62729 => conv_std_logic_vector(8, 8),
62730 => conv_std_logic_vector(9, 8),
62731 => conv_std_logic_vector(10, 8),
62732 => conv_std_logic_vector(11, 8),
62733 => conv_std_logic_vector(12, 8),
62734 => conv_std_logic_vector(13, 8),
62735 => conv_std_logic_vector(14, 8),
62736 => conv_std_logic_vector(15, 8),
62737 => conv_std_logic_vector(16, 8),
62738 => conv_std_logic_vector(17, 8),
62739 => conv_std_logic_vector(18, 8),
62740 => conv_std_logic_vector(19, 8),
62741 => conv_std_logic_vector(20, 8),
62742 => conv_std_logic_vector(21, 8),
62743 => conv_std_logic_vector(22, 8),
62744 => conv_std_logic_vector(22, 8),
62745 => conv_std_logic_vector(23, 8),
62746 => conv_std_logic_vector(24, 8),
62747 => conv_std_logic_vector(25, 8),
62748 => conv_std_logic_vector(26, 8),
62749 => conv_std_logic_vector(27, 8),
62750 => conv_std_logic_vector(28, 8),
62751 => conv_std_logic_vector(29, 8),
62752 => conv_std_logic_vector(30, 8),
62753 => conv_std_logic_vector(31, 8),
62754 => conv_std_logic_vector(32, 8),
62755 => conv_std_logic_vector(33, 8),
62756 => conv_std_logic_vector(34, 8),
62757 => conv_std_logic_vector(35, 8),
62758 => conv_std_logic_vector(36, 8),
62759 => conv_std_logic_vector(37, 8),
62760 => conv_std_logic_vector(38, 8),
62761 => conv_std_logic_vector(39, 8),
62762 => conv_std_logic_vector(40, 8),
62763 => conv_std_logic_vector(41, 8),
62764 => conv_std_logic_vector(42, 8),
62765 => conv_std_logic_vector(43, 8),
62766 => conv_std_logic_vector(44, 8),
62767 => conv_std_logic_vector(44, 8),
62768 => conv_std_logic_vector(45, 8),
62769 => conv_std_logic_vector(46, 8),
62770 => conv_std_logic_vector(47, 8),
62771 => conv_std_logic_vector(48, 8),
62772 => conv_std_logic_vector(49, 8),
62773 => conv_std_logic_vector(50, 8),
62774 => conv_std_logic_vector(51, 8),
62775 => conv_std_logic_vector(52, 8),
62776 => conv_std_logic_vector(53, 8),
62777 => conv_std_logic_vector(54, 8),
62778 => conv_std_logic_vector(55, 8),
62779 => conv_std_logic_vector(56, 8),
62780 => conv_std_logic_vector(57, 8),
62781 => conv_std_logic_vector(58, 8),
62782 => conv_std_logic_vector(59, 8),
62783 => conv_std_logic_vector(60, 8),
62784 => conv_std_logic_vector(61, 8),
62785 => conv_std_logic_vector(62, 8),
62786 => conv_std_logic_vector(63, 8),
62787 => conv_std_logic_vector(64, 8),
62788 => conv_std_logic_vector(65, 8),
62789 => conv_std_logic_vector(66, 8),
62790 => conv_std_logic_vector(66, 8),
62791 => conv_std_logic_vector(67, 8),
62792 => conv_std_logic_vector(68, 8),
62793 => conv_std_logic_vector(69, 8),
62794 => conv_std_logic_vector(70, 8),
62795 => conv_std_logic_vector(71, 8),
62796 => conv_std_logic_vector(72, 8),
62797 => conv_std_logic_vector(73, 8),
62798 => conv_std_logic_vector(74, 8),
62799 => conv_std_logic_vector(75, 8),
62800 => conv_std_logic_vector(76, 8),
62801 => conv_std_logic_vector(77, 8),
62802 => conv_std_logic_vector(78, 8),
62803 => conv_std_logic_vector(79, 8),
62804 => conv_std_logic_vector(80, 8),
62805 => conv_std_logic_vector(81, 8),
62806 => conv_std_logic_vector(82, 8),
62807 => conv_std_logic_vector(83, 8),
62808 => conv_std_logic_vector(84, 8),
62809 => conv_std_logic_vector(85, 8),
62810 => conv_std_logic_vector(86, 8),
62811 => conv_std_logic_vector(87, 8),
62812 => conv_std_logic_vector(88, 8),
62813 => conv_std_logic_vector(89, 8),
62814 => conv_std_logic_vector(89, 8),
62815 => conv_std_logic_vector(90, 8),
62816 => conv_std_logic_vector(91, 8),
62817 => conv_std_logic_vector(92, 8),
62818 => conv_std_logic_vector(93, 8),
62819 => conv_std_logic_vector(94, 8),
62820 => conv_std_logic_vector(95, 8),
62821 => conv_std_logic_vector(96, 8),
62822 => conv_std_logic_vector(97, 8),
62823 => conv_std_logic_vector(98, 8),
62824 => conv_std_logic_vector(99, 8),
62825 => conv_std_logic_vector(100, 8),
62826 => conv_std_logic_vector(101, 8),
62827 => conv_std_logic_vector(102, 8),
62828 => conv_std_logic_vector(103, 8),
62829 => conv_std_logic_vector(104, 8),
62830 => conv_std_logic_vector(105, 8),
62831 => conv_std_logic_vector(106, 8),
62832 => conv_std_logic_vector(107, 8),
62833 => conv_std_logic_vector(108, 8),
62834 => conv_std_logic_vector(109, 8),
62835 => conv_std_logic_vector(110, 8),
62836 => conv_std_logic_vector(111, 8),
62837 => conv_std_logic_vector(111, 8),
62838 => conv_std_logic_vector(112, 8),
62839 => conv_std_logic_vector(113, 8),
62840 => conv_std_logic_vector(114, 8),
62841 => conv_std_logic_vector(115, 8),
62842 => conv_std_logic_vector(116, 8),
62843 => conv_std_logic_vector(117, 8),
62844 => conv_std_logic_vector(118, 8),
62845 => conv_std_logic_vector(119, 8),
62846 => conv_std_logic_vector(120, 8),
62847 => conv_std_logic_vector(121, 8),
62848 => conv_std_logic_vector(122, 8),
62849 => conv_std_logic_vector(123, 8),
62850 => conv_std_logic_vector(124, 8),
62851 => conv_std_logic_vector(125, 8),
62852 => conv_std_logic_vector(126, 8),
62853 => conv_std_logic_vector(127, 8),
62854 => conv_std_logic_vector(128, 8),
62855 => conv_std_logic_vector(129, 8),
62856 => conv_std_logic_vector(130, 8),
62857 => conv_std_logic_vector(131, 8),
62858 => conv_std_logic_vector(132, 8),
62859 => conv_std_logic_vector(133, 8),
62860 => conv_std_logic_vector(133, 8),
62861 => conv_std_logic_vector(134, 8),
62862 => conv_std_logic_vector(135, 8),
62863 => conv_std_logic_vector(136, 8),
62864 => conv_std_logic_vector(137, 8),
62865 => conv_std_logic_vector(138, 8),
62866 => conv_std_logic_vector(139, 8),
62867 => conv_std_logic_vector(140, 8),
62868 => conv_std_logic_vector(141, 8),
62869 => conv_std_logic_vector(142, 8),
62870 => conv_std_logic_vector(143, 8),
62871 => conv_std_logic_vector(144, 8),
62872 => conv_std_logic_vector(145, 8),
62873 => conv_std_logic_vector(146, 8),
62874 => conv_std_logic_vector(147, 8),
62875 => conv_std_logic_vector(148, 8),
62876 => conv_std_logic_vector(149, 8),
62877 => conv_std_logic_vector(150, 8),
62878 => conv_std_logic_vector(151, 8),
62879 => conv_std_logic_vector(152, 8),
62880 => conv_std_logic_vector(153, 8),
62881 => conv_std_logic_vector(154, 8),
62882 => conv_std_logic_vector(155, 8),
62883 => conv_std_logic_vector(155, 8),
62884 => conv_std_logic_vector(156, 8),
62885 => conv_std_logic_vector(157, 8),
62886 => conv_std_logic_vector(158, 8),
62887 => conv_std_logic_vector(159, 8),
62888 => conv_std_logic_vector(160, 8),
62889 => conv_std_logic_vector(161, 8),
62890 => conv_std_logic_vector(162, 8),
62891 => conv_std_logic_vector(163, 8),
62892 => conv_std_logic_vector(164, 8),
62893 => conv_std_logic_vector(165, 8),
62894 => conv_std_logic_vector(166, 8),
62895 => conv_std_logic_vector(167, 8),
62896 => conv_std_logic_vector(168, 8),
62897 => conv_std_logic_vector(169, 8),
62898 => conv_std_logic_vector(170, 8),
62899 => conv_std_logic_vector(171, 8),
62900 => conv_std_logic_vector(172, 8),
62901 => conv_std_logic_vector(173, 8),
62902 => conv_std_logic_vector(174, 8),
62903 => conv_std_logic_vector(175, 8),
62904 => conv_std_logic_vector(176, 8),
62905 => conv_std_logic_vector(177, 8),
62906 => conv_std_logic_vector(178, 8),
62907 => conv_std_logic_vector(178, 8),
62908 => conv_std_logic_vector(179, 8),
62909 => conv_std_logic_vector(180, 8),
62910 => conv_std_logic_vector(181, 8),
62911 => conv_std_logic_vector(182, 8),
62912 => conv_std_logic_vector(183, 8),
62913 => conv_std_logic_vector(184, 8),
62914 => conv_std_logic_vector(185, 8),
62915 => conv_std_logic_vector(186, 8),
62916 => conv_std_logic_vector(187, 8),
62917 => conv_std_logic_vector(188, 8),
62918 => conv_std_logic_vector(189, 8),
62919 => conv_std_logic_vector(190, 8),
62920 => conv_std_logic_vector(191, 8),
62921 => conv_std_logic_vector(192, 8),
62922 => conv_std_logic_vector(193, 8),
62923 => conv_std_logic_vector(194, 8),
62924 => conv_std_logic_vector(195, 8),
62925 => conv_std_logic_vector(196, 8),
62926 => conv_std_logic_vector(197, 8),
62927 => conv_std_logic_vector(198, 8),
62928 => conv_std_logic_vector(199, 8),
62929 => conv_std_logic_vector(200, 8),
62930 => conv_std_logic_vector(200, 8),
62931 => conv_std_logic_vector(201, 8),
62932 => conv_std_logic_vector(202, 8),
62933 => conv_std_logic_vector(203, 8),
62934 => conv_std_logic_vector(204, 8),
62935 => conv_std_logic_vector(205, 8),
62936 => conv_std_logic_vector(206, 8),
62937 => conv_std_logic_vector(207, 8),
62938 => conv_std_logic_vector(208, 8),
62939 => conv_std_logic_vector(209, 8),
62940 => conv_std_logic_vector(210, 8),
62941 => conv_std_logic_vector(211, 8),
62942 => conv_std_logic_vector(212, 8),
62943 => conv_std_logic_vector(213, 8),
62944 => conv_std_logic_vector(214, 8),
62945 => conv_std_logic_vector(215, 8),
62946 => conv_std_logic_vector(216, 8),
62947 => conv_std_logic_vector(217, 8),
62948 => conv_std_logic_vector(218, 8),
62949 => conv_std_logic_vector(219, 8),
62950 => conv_std_logic_vector(220, 8),
62951 => conv_std_logic_vector(221, 8),
62952 => conv_std_logic_vector(222, 8),
62953 => conv_std_logic_vector(222, 8),
62954 => conv_std_logic_vector(223, 8),
62955 => conv_std_logic_vector(224, 8),
62956 => conv_std_logic_vector(225, 8),
62957 => conv_std_logic_vector(226, 8),
62958 => conv_std_logic_vector(227, 8),
62959 => conv_std_logic_vector(228, 8),
62960 => conv_std_logic_vector(229, 8),
62961 => conv_std_logic_vector(230, 8),
62962 => conv_std_logic_vector(231, 8),
62963 => conv_std_logic_vector(232, 8),
62964 => conv_std_logic_vector(233, 8),
62965 => conv_std_logic_vector(234, 8),
62966 => conv_std_logic_vector(235, 8),
62967 => conv_std_logic_vector(236, 8),
62968 => conv_std_logic_vector(237, 8),
62969 => conv_std_logic_vector(238, 8),
62970 => conv_std_logic_vector(239, 8),
62971 => conv_std_logic_vector(240, 8),
62972 => conv_std_logic_vector(241, 8),
62973 => conv_std_logic_vector(242, 8),
62974 => conv_std_logic_vector(243, 8),
62975 => conv_std_logic_vector(244, 8),
62976 => conv_std_logic_vector(0, 8),
62977 => conv_std_logic_vector(0, 8),
62978 => conv_std_logic_vector(1, 8),
62979 => conv_std_logic_vector(2, 8),
62980 => conv_std_logic_vector(3, 8),
62981 => conv_std_logic_vector(4, 8),
62982 => conv_std_logic_vector(5, 8),
62983 => conv_std_logic_vector(6, 8),
62984 => conv_std_logic_vector(7, 8),
62985 => conv_std_logic_vector(8, 8),
62986 => conv_std_logic_vector(9, 8),
62987 => conv_std_logic_vector(10, 8),
62988 => conv_std_logic_vector(11, 8),
62989 => conv_std_logic_vector(12, 8),
62990 => conv_std_logic_vector(13, 8),
62991 => conv_std_logic_vector(14, 8),
62992 => conv_std_logic_vector(15, 8),
62993 => conv_std_logic_vector(16, 8),
62994 => conv_std_logic_vector(17, 8),
62995 => conv_std_logic_vector(18, 8),
62996 => conv_std_logic_vector(19, 8),
62997 => conv_std_logic_vector(20, 8),
62998 => conv_std_logic_vector(21, 8),
62999 => conv_std_logic_vector(22, 8),
63000 => conv_std_logic_vector(23, 8),
63001 => conv_std_logic_vector(24, 8),
63002 => conv_std_logic_vector(24, 8),
63003 => conv_std_logic_vector(25, 8),
63004 => conv_std_logic_vector(26, 8),
63005 => conv_std_logic_vector(27, 8),
63006 => conv_std_logic_vector(28, 8),
63007 => conv_std_logic_vector(29, 8),
63008 => conv_std_logic_vector(30, 8),
63009 => conv_std_logic_vector(31, 8),
63010 => conv_std_logic_vector(32, 8),
63011 => conv_std_logic_vector(33, 8),
63012 => conv_std_logic_vector(34, 8),
63013 => conv_std_logic_vector(35, 8),
63014 => conv_std_logic_vector(36, 8),
63015 => conv_std_logic_vector(37, 8),
63016 => conv_std_logic_vector(38, 8),
63017 => conv_std_logic_vector(39, 8),
63018 => conv_std_logic_vector(40, 8),
63019 => conv_std_logic_vector(41, 8),
63020 => conv_std_logic_vector(42, 8),
63021 => conv_std_logic_vector(43, 8),
63022 => conv_std_logic_vector(44, 8),
63023 => conv_std_logic_vector(45, 8),
63024 => conv_std_logic_vector(46, 8),
63025 => conv_std_logic_vector(47, 8),
63026 => conv_std_logic_vector(48, 8),
63027 => conv_std_logic_vector(49, 8),
63028 => conv_std_logic_vector(49, 8),
63029 => conv_std_logic_vector(50, 8),
63030 => conv_std_logic_vector(51, 8),
63031 => conv_std_logic_vector(52, 8),
63032 => conv_std_logic_vector(53, 8),
63033 => conv_std_logic_vector(54, 8),
63034 => conv_std_logic_vector(55, 8),
63035 => conv_std_logic_vector(56, 8),
63036 => conv_std_logic_vector(57, 8),
63037 => conv_std_logic_vector(58, 8),
63038 => conv_std_logic_vector(59, 8),
63039 => conv_std_logic_vector(60, 8),
63040 => conv_std_logic_vector(61, 8),
63041 => conv_std_logic_vector(62, 8),
63042 => conv_std_logic_vector(63, 8),
63043 => conv_std_logic_vector(64, 8),
63044 => conv_std_logic_vector(65, 8),
63045 => conv_std_logic_vector(66, 8),
63046 => conv_std_logic_vector(67, 8),
63047 => conv_std_logic_vector(68, 8),
63048 => conv_std_logic_vector(69, 8),
63049 => conv_std_logic_vector(70, 8),
63050 => conv_std_logic_vector(71, 8),
63051 => conv_std_logic_vector(72, 8),
63052 => conv_std_logic_vector(73, 8),
63053 => conv_std_logic_vector(73, 8),
63054 => conv_std_logic_vector(74, 8),
63055 => conv_std_logic_vector(75, 8),
63056 => conv_std_logic_vector(76, 8),
63057 => conv_std_logic_vector(77, 8),
63058 => conv_std_logic_vector(78, 8),
63059 => conv_std_logic_vector(79, 8),
63060 => conv_std_logic_vector(80, 8),
63061 => conv_std_logic_vector(81, 8),
63062 => conv_std_logic_vector(82, 8),
63063 => conv_std_logic_vector(83, 8),
63064 => conv_std_logic_vector(84, 8),
63065 => conv_std_logic_vector(85, 8),
63066 => conv_std_logic_vector(86, 8),
63067 => conv_std_logic_vector(87, 8),
63068 => conv_std_logic_vector(88, 8),
63069 => conv_std_logic_vector(89, 8),
63070 => conv_std_logic_vector(90, 8),
63071 => conv_std_logic_vector(91, 8),
63072 => conv_std_logic_vector(92, 8),
63073 => conv_std_logic_vector(93, 8),
63074 => conv_std_logic_vector(94, 8),
63075 => conv_std_logic_vector(95, 8),
63076 => conv_std_logic_vector(96, 8),
63077 => conv_std_logic_vector(97, 8),
63078 => conv_std_logic_vector(98, 8),
63079 => conv_std_logic_vector(98, 8),
63080 => conv_std_logic_vector(99, 8),
63081 => conv_std_logic_vector(100, 8),
63082 => conv_std_logic_vector(101, 8),
63083 => conv_std_logic_vector(102, 8),
63084 => conv_std_logic_vector(103, 8),
63085 => conv_std_logic_vector(104, 8),
63086 => conv_std_logic_vector(105, 8),
63087 => conv_std_logic_vector(106, 8),
63088 => conv_std_logic_vector(107, 8),
63089 => conv_std_logic_vector(108, 8),
63090 => conv_std_logic_vector(109, 8),
63091 => conv_std_logic_vector(110, 8),
63092 => conv_std_logic_vector(111, 8),
63093 => conv_std_logic_vector(112, 8),
63094 => conv_std_logic_vector(113, 8),
63095 => conv_std_logic_vector(114, 8),
63096 => conv_std_logic_vector(115, 8),
63097 => conv_std_logic_vector(116, 8),
63098 => conv_std_logic_vector(117, 8),
63099 => conv_std_logic_vector(118, 8),
63100 => conv_std_logic_vector(119, 8),
63101 => conv_std_logic_vector(120, 8),
63102 => conv_std_logic_vector(121, 8),
63103 => conv_std_logic_vector(122, 8),
63104 => conv_std_logic_vector(123, 8),
63105 => conv_std_logic_vector(123, 8),
63106 => conv_std_logic_vector(124, 8),
63107 => conv_std_logic_vector(125, 8),
63108 => conv_std_logic_vector(126, 8),
63109 => conv_std_logic_vector(127, 8),
63110 => conv_std_logic_vector(128, 8),
63111 => conv_std_logic_vector(129, 8),
63112 => conv_std_logic_vector(130, 8),
63113 => conv_std_logic_vector(131, 8),
63114 => conv_std_logic_vector(132, 8),
63115 => conv_std_logic_vector(133, 8),
63116 => conv_std_logic_vector(134, 8),
63117 => conv_std_logic_vector(135, 8),
63118 => conv_std_logic_vector(136, 8),
63119 => conv_std_logic_vector(137, 8),
63120 => conv_std_logic_vector(138, 8),
63121 => conv_std_logic_vector(139, 8),
63122 => conv_std_logic_vector(140, 8),
63123 => conv_std_logic_vector(141, 8),
63124 => conv_std_logic_vector(142, 8),
63125 => conv_std_logic_vector(143, 8),
63126 => conv_std_logic_vector(144, 8),
63127 => conv_std_logic_vector(145, 8),
63128 => conv_std_logic_vector(146, 8),
63129 => conv_std_logic_vector(147, 8),
63130 => conv_std_logic_vector(147, 8),
63131 => conv_std_logic_vector(148, 8),
63132 => conv_std_logic_vector(149, 8),
63133 => conv_std_logic_vector(150, 8),
63134 => conv_std_logic_vector(151, 8),
63135 => conv_std_logic_vector(152, 8),
63136 => conv_std_logic_vector(153, 8),
63137 => conv_std_logic_vector(154, 8),
63138 => conv_std_logic_vector(155, 8),
63139 => conv_std_logic_vector(156, 8),
63140 => conv_std_logic_vector(157, 8),
63141 => conv_std_logic_vector(158, 8),
63142 => conv_std_logic_vector(159, 8),
63143 => conv_std_logic_vector(160, 8),
63144 => conv_std_logic_vector(161, 8),
63145 => conv_std_logic_vector(162, 8),
63146 => conv_std_logic_vector(163, 8),
63147 => conv_std_logic_vector(164, 8),
63148 => conv_std_logic_vector(165, 8),
63149 => conv_std_logic_vector(166, 8),
63150 => conv_std_logic_vector(167, 8),
63151 => conv_std_logic_vector(168, 8),
63152 => conv_std_logic_vector(169, 8),
63153 => conv_std_logic_vector(170, 8),
63154 => conv_std_logic_vector(171, 8),
63155 => conv_std_logic_vector(172, 8),
63156 => conv_std_logic_vector(172, 8),
63157 => conv_std_logic_vector(173, 8),
63158 => conv_std_logic_vector(174, 8),
63159 => conv_std_logic_vector(175, 8),
63160 => conv_std_logic_vector(176, 8),
63161 => conv_std_logic_vector(177, 8),
63162 => conv_std_logic_vector(178, 8),
63163 => conv_std_logic_vector(179, 8),
63164 => conv_std_logic_vector(180, 8),
63165 => conv_std_logic_vector(181, 8),
63166 => conv_std_logic_vector(182, 8),
63167 => conv_std_logic_vector(183, 8),
63168 => conv_std_logic_vector(184, 8),
63169 => conv_std_logic_vector(185, 8),
63170 => conv_std_logic_vector(186, 8),
63171 => conv_std_logic_vector(187, 8),
63172 => conv_std_logic_vector(188, 8),
63173 => conv_std_logic_vector(189, 8),
63174 => conv_std_logic_vector(190, 8),
63175 => conv_std_logic_vector(191, 8),
63176 => conv_std_logic_vector(192, 8),
63177 => conv_std_logic_vector(193, 8),
63178 => conv_std_logic_vector(194, 8),
63179 => conv_std_logic_vector(195, 8),
63180 => conv_std_logic_vector(196, 8),
63181 => conv_std_logic_vector(196, 8),
63182 => conv_std_logic_vector(197, 8),
63183 => conv_std_logic_vector(198, 8),
63184 => conv_std_logic_vector(199, 8),
63185 => conv_std_logic_vector(200, 8),
63186 => conv_std_logic_vector(201, 8),
63187 => conv_std_logic_vector(202, 8),
63188 => conv_std_logic_vector(203, 8),
63189 => conv_std_logic_vector(204, 8),
63190 => conv_std_logic_vector(205, 8),
63191 => conv_std_logic_vector(206, 8),
63192 => conv_std_logic_vector(207, 8),
63193 => conv_std_logic_vector(208, 8),
63194 => conv_std_logic_vector(209, 8),
63195 => conv_std_logic_vector(210, 8),
63196 => conv_std_logic_vector(211, 8),
63197 => conv_std_logic_vector(212, 8),
63198 => conv_std_logic_vector(213, 8),
63199 => conv_std_logic_vector(214, 8),
63200 => conv_std_logic_vector(215, 8),
63201 => conv_std_logic_vector(216, 8),
63202 => conv_std_logic_vector(217, 8),
63203 => conv_std_logic_vector(218, 8),
63204 => conv_std_logic_vector(219, 8),
63205 => conv_std_logic_vector(220, 8),
63206 => conv_std_logic_vector(221, 8),
63207 => conv_std_logic_vector(221, 8),
63208 => conv_std_logic_vector(222, 8),
63209 => conv_std_logic_vector(223, 8),
63210 => conv_std_logic_vector(224, 8),
63211 => conv_std_logic_vector(225, 8),
63212 => conv_std_logic_vector(226, 8),
63213 => conv_std_logic_vector(227, 8),
63214 => conv_std_logic_vector(228, 8),
63215 => conv_std_logic_vector(229, 8),
63216 => conv_std_logic_vector(230, 8),
63217 => conv_std_logic_vector(231, 8),
63218 => conv_std_logic_vector(232, 8),
63219 => conv_std_logic_vector(233, 8),
63220 => conv_std_logic_vector(234, 8),
63221 => conv_std_logic_vector(235, 8),
63222 => conv_std_logic_vector(236, 8),
63223 => conv_std_logic_vector(237, 8),
63224 => conv_std_logic_vector(238, 8),
63225 => conv_std_logic_vector(239, 8),
63226 => conv_std_logic_vector(240, 8),
63227 => conv_std_logic_vector(241, 8),
63228 => conv_std_logic_vector(242, 8),
63229 => conv_std_logic_vector(243, 8),
63230 => conv_std_logic_vector(244, 8),
63231 => conv_std_logic_vector(245, 8),
63232 => conv_std_logic_vector(0, 8),
63233 => conv_std_logic_vector(0, 8),
63234 => conv_std_logic_vector(1, 8),
63235 => conv_std_logic_vector(2, 8),
63236 => conv_std_logic_vector(3, 8),
63237 => conv_std_logic_vector(4, 8),
63238 => conv_std_logic_vector(5, 8),
63239 => conv_std_logic_vector(6, 8),
63240 => conv_std_logic_vector(7, 8),
63241 => conv_std_logic_vector(8, 8),
63242 => conv_std_logic_vector(9, 8),
63243 => conv_std_logic_vector(10, 8),
63244 => conv_std_logic_vector(11, 8),
63245 => conv_std_logic_vector(12, 8),
63246 => conv_std_logic_vector(13, 8),
63247 => conv_std_logic_vector(14, 8),
63248 => conv_std_logic_vector(15, 8),
63249 => conv_std_logic_vector(16, 8),
63250 => conv_std_logic_vector(17, 8),
63251 => conv_std_logic_vector(18, 8),
63252 => conv_std_logic_vector(19, 8),
63253 => conv_std_logic_vector(20, 8),
63254 => conv_std_logic_vector(21, 8),
63255 => conv_std_logic_vector(22, 8),
63256 => conv_std_logic_vector(23, 8),
63257 => conv_std_logic_vector(24, 8),
63258 => conv_std_logic_vector(25, 8),
63259 => conv_std_logic_vector(26, 8),
63260 => conv_std_logic_vector(27, 8),
63261 => conv_std_logic_vector(27, 8),
63262 => conv_std_logic_vector(28, 8),
63263 => conv_std_logic_vector(29, 8),
63264 => conv_std_logic_vector(30, 8),
63265 => conv_std_logic_vector(31, 8),
63266 => conv_std_logic_vector(32, 8),
63267 => conv_std_logic_vector(33, 8),
63268 => conv_std_logic_vector(34, 8),
63269 => conv_std_logic_vector(35, 8),
63270 => conv_std_logic_vector(36, 8),
63271 => conv_std_logic_vector(37, 8),
63272 => conv_std_logic_vector(38, 8),
63273 => conv_std_logic_vector(39, 8),
63274 => conv_std_logic_vector(40, 8),
63275 => conv_std_logic_vector(41, 8),
63276 => conv_std_logic_vector(42, 8),
63277 => conv_std_logic_vector(43, 8),
63278 => conv_std_logic_vector(44, 8),
63279 => conv_std_logic_vector(45, 8),
63280 => conv_std_logic_vector(46, 8),
63281 => conv_std_logic_vector(47, 8),
63282 => conv_std_logic_vector(48, 8),
63283 => conv_std_logic_vector(49, 8),
63284 => conv_std_logic_vector(50, 8),
63285 => conv_std_logic_vector(51, 8),
63286 => conv_std_logic_vector(52, 8),
63287 => conv_std_logic_vector(53, 8),
63288 => conv_std_logic_vector(54, 8),
63289 => conv_std_logic_vector(54, 8),
63290 => conv_std_logic_vector(55, 8),
63291 => conv_std_logic_vector(56, 8),
63292 => conv_std_logic_vector(57, 8),
63293 => conv_std_logic_vector(58, 8),
63294 => conv_std_logic_vector(59, 8),
63295 => conv_std_logic_vector(60, 8),
63296 => conv_std_logic_vector(61, 8),
63297 => conv_std_logic_vector(62, 8),
63298 => conv_std_logic_vector(63, 8),
63299 => conv_std_logic_vector(64, 8),
63300 => conv_std_logic_vector(65, 8),
63301 => conv_std_logic_vector(66, 8),
63302 => conv_std_logic_vector(67, 8),
63303 => conv_std_logic_vector(68, 8),
63304 => conv_std_logic_vector(69, 8),
63305 => conv_std_logic_vector(70, 8),
63306 => conv_std_logic_vector(71, 8),
63307 => conv_std_logic_vector(72, 8),
63308 => conv_std_logic_vector(73, 8),
63309 => conv_std_logic_vector(74, 8),
63310 => conv_std_logic_vector(75, 8),
63311 => conv_std_logic_vector(76, 8),
63312 => conv_std_logic_vector(77, 8),
63313 => conv_std_logic_vector(78, 8),
63314 => conv_std_logic_vector(79, 8),
63315 => conv_std_logic_vector(80, 8),
63316 => conv_std_logic_vector(81, 8),
63317 => conv_std_logic_vector(82, 8),
63318 => conv_std_logic_vector(82, 8),
63319 => conv_std_logic_vector(83, 8),
63320 => conv_std_logic_vector(84, 8),
63321 => conv_std_logic_vector(85, 8),
63322 => conv_std_logic_vector(86, 8),
63323 => conv_std_logic_vector(87, 8),
63324 => conv_std_logic_vector(88, 8),
63325 => conv_std_logic_vector(89, 8),
63326 => conv_std_logic_vector(90, 8),
63327 => conv_std_logic_vector(91, 8),
63328 => conv_std_logic_vector(92, 8),
63329 => conv_std_logic_vector(93, 8),
63330 => conv_std_logic_vector(94, 8),
63331 => conv_std_logic_vector(95, 8),
63332 => conv_std_logic_vector(96, 8),
63333 => conv_std_logic_vector(97, 8),
63334 => conv_std_logic_vector(98, 8),
63335 => conv_std_logic_vector(99, 8),
63336 => conv_std_logic_vector(100, 8),
63337 => conv_std_logic_vector(101, 8),
63338 => conv_std_logic_vector(102, 8),
63339 => conv_std_logic_vector(103, 8),
63340 => conv_std_logic_vector(104, 8),
63341 => conv_std_logic_vector(105, 8),
63342 => conv_std_logic_vector(106, 8),
63343 => conv_std_logic_vector(107, 8),
63344 => conv_std_logic_vector(108, 8),
63345 => conv_std_logic_vector(109, 8),
63346 => conv_std_logic_vector(109, 8),
63347 => conv_std_logic_vector(110, 8),
63348 => conv_std_logic_vector(111, 8),
63349 => conv_std_logic_vector(112, 8),
63350 => conv_std_logic_vector(113, 8),
63351 => conv_std_logic_vector(114, 8),
63352 => conv_std_logic_vector(115, 8),
63353 => conv_std_logic_vector(116, 8),
63354 => conv_std_logic_vector(117, 8),
63355 => conv_std_logic_vector(118, 8),
63356 => conv_std_logic_vector(119, 8),
63357 => conv_std_logic_vector(120, 8),
63358 => conv_std_logic_vector(121, 8),
63359 => conv_std_logic_vector(122, 8),
63360 => conv_std_logic_vector(123, 8),
63361 => conv_std_logic_vector(124, 8),
63362 => conv_std_logic_vector(125, 8),
63363 => conv_std_logic_vector(126, 8),
63364 => conv_std_logic_vector(127, 8),
63365 => conv_std_logic_vector(128, 8),
63366 => conv_std_logic_vector(129, 8),
63367 => conv_std_logic_vector(130, 8),
63368 => conv_std_logic_vector(131, 8),
63369 => conv_std_logic_vector(132, 8),
63370 => conv_std_logic_vector(133, 8),
63371 => conv_std_logic_vector(134, 8),
63372 => conv_std_logic_vector(135, 8),
63373 => conv_std_logic_vector(136, 8),
63374 => conv_std_logic_vector(137, 8),
63375 => conv_std_logic_vector(137, 8),
63376 => conv_std_logic_vector(138, 8),
63377 => conv_std_logic_vector(139, 8),
63378 => conv_std_logic_vector(140, 8),
63379 => conv_std_logic_vector(141, 8),
63380 => conv_std_logic_vector(142, 8),
63381 => conv_std_logic_vector(143, 8),
63382 => conv_std_logic_vector(144, 8),
63383 => conv_std_logic_vector(145, 8),
63384 => conv_std_logic_vector(146, 8),
63385 => conv_std_logic_vector(147, 8),
63386 => conv_std_logic_vector(148, 8),
63387 => conv_std_logic_vector(149, 8),
63388 => conv_std_logic_vector(150, 8),
63389 => conv_std_logic_vector(151, 8),
63390 => conv_std_logic_vector(152, 8),
63391 => conv_std_logic_vector(153, 8),
63392 => conv_std_logic_vector(154, 8),
63393 => conv_std_logic_vector(155, 8),
63394 => conv_std_logic_vector(156, 8),
63395 => conv_std_logic_vector(157, 8),
63396 => conv_std_logic_vector(158, 8),
63397 => conv_std_logic_vector(159, 8),
63398 => conv_std_logic_vector(160, 8),
63399 => conv_std_logic_vector(161, 8),
63400 => conv_std_logic_vector(162, 8),
63401 => conv_std_logic_vector(163, 8),
63402 => conv_std_logic_vector(164, 8),
63403 => conv_std_logic_vector(164, 8),
63404 => conv_std_logic_vector(165, 8),
63405 => conv_std_logic_vector(166, 8),
63406 => conv_std_logic_vector(167, 8),
63407 => conv_std_logic_vector(168, 8),
63408 => conv_std_logic_vector(169, 8),
63409 => conv_std_logic_vector(170, 8),
63410 => conv_std_logic_vector(171, 8),
63411 => conv_std_logic_vector(172, 8),
63412 => conv_std_logic_vector(173, 8),
63413 => conv_std_logic_vector(174, 8),
63414 => conv_std_logic_vector(175, 8),
63415 => conv_std_logic_vector(176, 8),
63416 => conv_std_logic_vector(177, 8),
63417 => conv_std_logic_vector(178, 8),
63418 => conv_std_logic_vector(179, 8),
63419 => conv_std_logic_vector(180, 8),
63420 => conv_std_logic_vector(181, 8),
63421 => conv_std_logic_vector(182, 8),
63422 => conv_std_logic_vector(183, 8),
63423 => conv_std_logic_vector(184, 8),
63424 => conv_std_logic_vector(185, 8),
63425 => conv_std_logic_vector(186, 8),
63426 => conv_std_logic_vector(187, 8),
63427 => conv_std_logic_vector(188, 8),
63428 => conv_std_logic_vector(189, 8),
63429 => conv_std_logic_vector(190, 8),
63430 => conv_std_logic_vector(191, 8),
63431 => conv_std_logic_vector(192, 8),
63432 => conv_std_logic_vector(192, 8),
63433 => conv_std_logic_vector(193, 8),
63434 => conv_std_logic_vector(194, 8),
63435 => conv_std_logic_vector(195, 8),
63436 => conv_std_logic_vector(196, 8),
63437 => conv_std_logic_vector(197, 8),
63438 => conv_std_logic_vector(198, 8),
63439 => conv_std_logic_vector(199, 8),
63440 => conv_std_logic_vector(200, 8),
63441 => conv_std_logic_vector(201, 8),
63442 => conv_std_logic_vector(202, 8),
63443 => conv_std_logic_vector(203, 8),
63444 => conv_std_logic_vector(204, 8),
63445 => conv_std_logic_vector(205, 8),
63446 => conv_std_logic_vector(206, 8),
63447 => conv_std_logic_vector(207, 8),
63448 => conv_std_logic_vector(208, 8),
63449 => conv_std_logic_vector(209, 8),
63450 => conv_std_logic_vector(210, 8),
63451 => conv_std_logic_vector(211, 8),
63452 => conv_std_logic_vector(212, 8),
63453 => conv_std_logic_vector(213, 8),
63454 => conv_std_logic_vector(214, 8),
63455 => conv_std_logic_vector(215, 8),
63456 => conv_std_logic_vector(216, 8),
63457 => conv_std_logic_vector(217, 8),
63458 => conv_std_logic_vector(218, 8),
63459 => conv_std_logic_vector(219, 8),
63460 => conv_std_logic_vector(219, 8),
63461 => conv_std_logic_vector(220, 8),
63462 => conv_std_logic_vector(221, 8),
63463 => conv_std_logic_vector(222, 8),
63464 => conv_std_logic_vector(223, 8),
63465 => conv_std_logic_vector(224, 8),
63466 => conv_std_logic_vector(225, 8),
63467 => conv_std_logic_vector(226, 8),
63468 => conv_std_logic_vector(227, 8),
63469 => conv_std_logic_vector(228, 8),
63470 => conv_std_logic_vector(229, 8),
63471 => conv_std_logic_vector(230, 8),
63472 => conv_std_logic_vector(231, 8),
63473 => conv_std_logic_vector(232, 8),
63474 => conv_std_logic_vector(233, 8),
63475 => conv_std_logic_vector(234, 8),
63476 => conv_std_logic_vector(235, 8),
63477 => conv_std_logic_vector(236, 8),
63478 => conv_std_logic_vector(237, 8),
63479 => conv_std_logic_vector(238, 8),
63480 => conv_std_logic_vector(239, 8),
63481 => conv_std_logic_vector(240, 8),
63482 => conv_std_logic_vector(241, 8),
63483 => conv_std_logic_vector(242, 8),
63484 => conv_std_logic_vector(243, 8),
63485 => conv_std_logic_vector(244, 8),
63486 => conv_std_logic_vector(245, 8),
63487 => conv_std_logic_vector(246, 8),
63488 => conv_std_logic_vector(0, 8),
63489 => conv_std_logic_vector(0, 8),
63490 => conv_std_logic_vector(1, 8),
63491 => conv_std_logic_vector(2, 8),
63492 => conv_std_logic_vector(3, 8),
63493 => conv_std_logic_vector(4, 8),
63494 => conv_std_logic_vector(5, 8),
63495 => conv_std_logic_vector(6, 8),
63496 => conv_std_logic_vector(7, 8),
63497 => conv_std_logic_vector(8, 8),
63498 => conv_std_logic_vector(9, 8),
63499 => conv_std_logic_vector(10, 8),
63500 => conv_std_logic_vector(11, 8),
63501 => conv_std_logic_vector(12, 8),
63502 => conv_std_logic_vector(13, 8),
63503 => conv_std_logic_vector(14, 8),
63504 => conv_std_logic_vector(15, 8),
63505 => conv_std_logic_vector(16, 8),
63506 => conv_std_logic_vector(17, 8),
63507 => conv_std_logic_vector(18, 8),
63508 => conv_std_logic_vector(19, 8),
63509 => conv_std_logic_vector(20, 8),
63510 => conv_std_logic_vector(21, 8),
63511 => conv_std_logic_vector(22, 8),
63512 => conv_std_logic_vector(23, 8),
63513 => conv_std_logic_vector(24, 8),
63514 => conv_std_logic_vector(25, 8),
63515 => conv_std_logic_vector(26, 8),
63516 => conv_std_logic_vector(27, 8),
63517 => conv_std_logic_vector(28, 8),
63518 => conv_std_logic_vector(29, 8),
63519 => conv_std_logic_vector(30, 8),
63520 => conv_std_logic_vector(31, 8),
63521 => conv_std_logic_vector(31, 8),
63522 => conv_std_logic_vector(32, 8),
63523 => conv_std_logic_vector(33, 8),
63524 => conv_std_logic_vector(34, 8),
63525 => conv_std_logic_vector(35, 8),
63526 => conv_std_logic_vector(36, 8),
63527 => conv_std_logic_vector(37, 8),
63528 => conv_std_logic_vector(38, 8),
63529 => conv_std_logic_vector(39, 8),
63530 => conv_std_logic_vector(40, 8),
63531 => conv_std_logic_vector(41, 8),
63532 => conv_std_logic_vector(42, 8),
63533 => conv_std_logic_vector(43, 8),
63534 => conv_std_logic_vector(44, 8),
63535 => conv_std_logic_vector(45, 8),
63536 => conv_std_logic_vector(46, 8),
63537 => conv_std_logic_vector(47, 8),
63538 => conv_std_logic_vector(48, 8),
63539 => conv_std_logic_vector(49, 8),
63540 => conv_std_logic_vector(50, 8),
63541 => conv_std_logic_vector(51, 8),
63542 => conv_std_logic_vector(52, 8),
63543 => conv_std_logic_vector(53, 8),
63544 => conv_std_logic_vector(54, 8),
63545 => conv_std_logic_vector(55, 8),
63546 => conv_std_logic_vector(56, 8),
63547 => conv_std_logic_vector(57, 8),
63548 => conv_std_logic_vector(58, 8),
63549 => conv_std_logic_vector(59, 8),
63550 => conv_std_logic_vector(60, 8),
63551 => conv_std_logic_vector(61, 8),
63552 => conv_std_logic_vector(62, 8),
63553 => conv_std_logic_vector(62, 8),
63554 => conv_std_logic_vector(63, 8),
63555 => conv_std_logic_vector(64, 8),
63556 => conv_std_logic_vector(65, 8),
63557 => conv_std_logic_vector(66, 8),
63558 => conv_std_logic_vector(67, 8),
63559 => conv_std_logic_vector(68, 8),
63560 => conv_std_logic_vector(69, 8),
63561 => conv_std_logic_vector(70, 8),
63562 => conv_std_logic_vector(71, 8),
63563 => conv_std_logic_vector(72, 8),
63564 => conv_std_logic_vector(73, 8),
63565 => conv_std_logic_vector(74, 8),
63566 => conv_std_logic_vector(75, 8),
63567 => conv_std_logic_vector(76, 8),
63568 => conv_std_logic_vector(77, 8),
63569 => conv_std_logic_vector(78, 8),
63570 => conv_std_logic_vector(79, 8),
63571 => conv_std_logic_vector(80, 8),
63572 => conv_std_logic_vector(81, 8),
63573 => conv_std_logic_vector(82, 8),
63574 => conv_std_logic_vector(83, 8),
63575 => conv_std_logic_vector(84, 8),
63576 => conv_std_logic_vector(85, 8),
63577 => conv_std_logic_vector(86, 8),
63578 => conv_std_logic_vector(87, 8),
63579 => conv_std_logic_vector(88, 8),
63580 => conv_std_logic_vector(89, 8),
63581 => conv_std_logic_vector(90, 8),
63582 => conv_std_logic_vector(91, 8),
63583 => conv_std_logic_vector(92, 8),
63584 => conv_std_logic_vector(93, 8),
63585 => conv_std_logic_vector(93, 8),
63586 => conv_std_logic_vector(94, 8),
63587 => conv_std_logic_vector(95, 8),
63588 => conv_std_logic_vector(96, 8),
63589 => conv_std_logic_vector(97, 8),
63590 => conv_std_logic_vector(98, 8),
63591 => conv_std_logic_vector(99, 8),
63592 => conv_std_logic_vector(100, 8),
63593 => conv_std_logic_vector(101, 8),
63594 => conv_std_logic_vector(102, 8),
63595 => conv_std_logic_vector(103, 8),
63596 => conv_std_logic_vector(104, 8),
63597 => conv_std_logic_vector(105, 8),
63598 => conv_std_logic_vector(106, 8),
63599 => conv_std_logic_vector(107, 8),
63600 => conv_std_logic_vector(108, 8),
63601 => conv_std_logic_vector(109, 8),
63602 => conv_std_logic_vector(110, 8),
63603 => conv_std_logic_vector(111, 8),
63604 => conv_std_logic_vector(112, 8),
63605 => conv_std_logic_vector(113, 8),
63606 => conv_std_logic_vector(114, 8),
63607 => conv_std_logic_vector(115, 8),
63608 => conv_std_logic_vector(116, 8),
63609 => conv_std_logic_vector(117, 8),
63610 => conv_std_logic_vector(118, 8),
63611 => conv_std_logic_vector(119, 8),
63612 => conv_std_logic_vector(120, 8),
63613 => conv_std_logic_vector(121, 8),
63614 => conv_std_logic_vector(122, 8),
63615 => conv_std_logic_vector(123, 8),
63616 => conv_std_logic_vector(124, 8),
63617 => conv_std_logic_vector(124, 8),
63618 => conv_std_logic_vector(125, 8),
63619 => conv_std_logic_vector(126, 8),
63620 => conv_std_logic_vector(127, 8),
63621 => conv_std_logic_vector(128, 8),
63622 => conv_std_logic_vector(129, 8),
63623 => conv_std_logic_vector(130, 8),
63624 => conv_std_logic_vector(131, 8),
63625 => conv_std_logic_vector(132, 8),
63626 => conv_std_logic_vector(133, 8),
63627 => conv_std_logic_vector(134, 8),
63628 => conv_std_logic_vector(135, 8),
63629 => conv_std_logic_vector(136, 8),
63630 => conv_std_logic_vector(137, 8),
63631 => conv_std_logic_vector(138, 8),
63632 => conv_std_logic_vector(139, 8),
63633 => conv_std_logic_vector(140, 8),
63634 => conv_std_logic_vector(141, 8),
63635 => conv_std_logic_vector(142, 8),
63636 => conv_std_logic_vector(143, 8),
63637 => conv_std_logic_vector(144, 8),
63638 => conv_std_logic_vector(145, 8),
63639 => conv_std_logic_vector(146, 8),
63640 => conv_std_logic_vector(147, 8),
63641 => conv_std_logic_vector(148, 8),
63642 => conv_std_logic_vector(149, 8),
63643 => conv_std_logic_vector(150, 8),
63644 => conv_std_logic_vector(151, 8),
63645 => conv_std_logic_vector(152, 8),
63646 => conv_std_logic_vector(153, 8),
63647 => conv_std_logic_vector(154, 8),
63648 => conv_std_logic_vector(155, 8),
63649 => conv_std_logic_vector(155, 8),
63650 => conv_std_logic_vector(156, 8),
63651 => conv_std_logic_vector(157, 8),
63652 => conv_std_logic_vector(158, 8),
63653 => conv_std_logic_vector(159, 8),
63654 => conv_std_logic_vector(160, 8),
63655 => conv_std_logic_vector(161, 8),
63656 => conv_std_logic_vector(162, 8),
63657 => conv_std_logic_vector(163, 8),
63658 => conv_std_logic_vector(164, 8),
63659 => conv_std_logic_vector(165, 8),
63660 => conv_std_logic_vector(166, 8),
63661 => conv_std_logic_vector(167, 8),
63662 => conv_std_logic_vector(168, 8),
63663 => conv_std_logic_vector(169, 8),
63664 => conv_std_logic_vector(170, 8),
63665 => conv_std_logic_vector(171, 8),
63666 => conv_std_logic_vector(172, 8),
63667 => conv_std_logic_vector(173, 8),
63668 => conv_std_logic_vector(174, 8),
63669 => conv_std_logic_vector(175, 8),
63670 => conv_std_logic_vector(176, 8),
63671 => conv_std_logic_vector(177, 8),
63672 => conv_std_logic_vector(178, 8),
63673 => conv_std_logic_vector(179, 8),
63674 => conv_std_logic_vector(180, 8),
63675 => conv_std_logic_vector(181, 8),
63676 => conv_std_logic_vector(182, 8),
63677 => conv_std_logic_vector(183, 8),
63678 => conv_std_logic_vector(184, 8),
63679 => conv_std_logic_vector(185, 8),
63680 => conv_std_logic_vector(186, 8),
63681 => conv_std_logic_vector(186, 8),
63682 => conv_std_logic_vector(187, 8),
63683 => conv_std_logic_vector(188, 8),
63684 => conv_std_logic_vector(189, 8),
63685 => conv_std_logic_vector(190, 8),
63686 => conv_std_logic_vector(191, 8),
63687 => conv_std_logic_vector(192, 8),
63688 => conv_std_logic_vector(193, 8),
63689 => conv_std_logic_vector(194, 8),
63690 => conv_std_logic_vector(195, 8),
63691 => conv_std_logic_vector(196, 8),
63692 => conv_std_logic_vector(197, 8),
63693 => conv_std_logic_vector(198, 8),
63694 => conv_std_logic_vector(199, 8),
63695 => conv_std_logic_vector(200, 8),
63696 => conv_std_logic_vector(201, 8),
63697 => conv_std_logic_vector(202, 8),
63698 => conv_std_logic_vector(203, 8),
63699 => conv_std_logic_vector(204, 8),
63700 => conv_std_logic_vector(205, 8),
63701 => conv_std_logic_vector(206, 8),
63702 => conv_std_logic_vector(207, 8),
63703 => conv_std_logic_vector(208, 8),
63704 => conv_std_logic_vector(209, 8),
63705 => conv_std_logic_vector(210, 8),
63706 => conv_std_logic_vector(211, 8),
63707 => conv_std_logic_vector(212, 8),
63708 => conv_std_logic_vector(213, 8),
63709 => conv_std_logic_vector(214, 8),
63710 => conv_std_logic_vector(215, 8),
63711 => conv_std_logic_vector(216, 8),
63712 => conv_std_logic_vector(217, 8),
63713 => conv_std_logic_vector(217, 8),
63714 => conv_std_logic_vector(218, 8),
63715 => conv_std_logic_vector(219, 8),
63716 => conv_std_logic_vector(220, 8),
63717 => conv_std_logic_vector(221, 8),
63718 => conv_std_logic_vector(222, 8),
63719 => conv_std_logic_vector(223, 8),
63720 => conv_std_logic_vector(224, 8),
63721 => conv_std_logic_vector(225, 8),
63722 => conv_std_logic_vector(226, 8),
63723 => conv_std_logic_vector(227, 8),
63724 => conv_std_logic_vector(228, 8),
63725 => conv_std_logic_vector(229, 8),
63726 => conv_std_logic_vector(230, 8),
63727 => conv_std_logic_vector(231, 8),
63728 => conv_std_logic_vector(232, 8),
63729 => conv_std_logic_vector(233, 8),
63730 => conv_std_logic_vector(234, 8),
63731 => conv_std_logic_vector(235, 8),
63732 => conv_std_logic_vector(236, 8),
63733 => conv_std_logic_vector(237, 8),
63734 => conv_std_logic_vector(238, 8),
63735 => conv_std_logic_vector(239, 8),
63736 => conv_std_logic_vector(240, 8),
63737 => conv_std_logic_vector(241, 8),
63738 => conv_std_logic_vector(242, 8),
63739 => conv_std_logic_vector(243, 8),
63740 => conv_std_logic_vector(244, 8),
63741 => conv_std_logic_vector(245, 8),
63742 => conv_std_logic_vector(246, 8),
63743 => conv_std_logic_vector(247, 8),
63744 => conv_std_logic_vector(0, 8),
63745 => conv_std_logic_vector(0, 8),
63746 => conv_std_logic_vector(1, 8),
63747 => conv_std_logic_vector(2, 8),
63748 => conv_std_logic_vector(3, 8),
63749 => conv_std_logic_vector(4, 8),
63750 => conv_std_logic_vector(5, 8),
63751 => conv_std_logic_vector(6, 8),
63752 => conv_std_logic_vector(7, 8),
63753 => conv_std_logic_vector(8, 8),
63754 => conv_std_logic_vector(9, 8),
63755 => conv_std_logic_vector(10, 8),
63756 => conv_std_logic_vector(11, 8),
63757 => conv_std_logic_vector(12, 8),
63758 => conv_std_logic_vector(13, 8),
63759 => conv_std_logic_vector(14, 8),
63760 => conv_std_logic_vector(15, 8),
63761 => conv_std_logic_vector(16, 8),
63762 => conv_std_logic_vector(17, 8),
63763 => conv_std_logic_vector(18, 8),
63764 => conv_std_logic_vector(19, 8),
63765 => conv_std_logic_vector(20, 8),
63766 => conv_std_logic_vector(21, 8),
63767 => conv_std_logic_vector(22, 8),
63768 => conv_std_logic_vector(23, 8),
63769 => conv_std_logic_vector(24, 8),
63770 => conv_std_logic_vector(25, 8),
63771 => conv_std_logic_vector(26, 8),
63772 => conv_std_logic_vector(27, 8),
63773 => conv_std_logic_vector(28, 8),
63774 => conv_std_logic_vector(29, 8),
63775 => conv_std_logic_vector(30, 8),
63776 => conv_std_logic_vector(31, 8),
63777 => conv_std_logic_vector(32, 8),
63778 => conv_std_logic_vector(33, 8),
63779 => conv_std_logic_vector(34, 8),
63780 => conv_std_logic_vector(35, 8),
63781 => conv_std_logic_vector(35, 8),
63782 => conv_std_logic_vector(36, 8),
63783 => conv_std_logic_vector(37, 8),
63784 => conv_std_logic_vector(38, 8),
63785 => conv_std_logic_vector(39, 8),
63786 => conv_std_logic_vector(40, 8),
63787 => conv_std_logic_vector(41, 8),
63788 => conv_std_logic_vector(42, 8),
63789 => conv_std_logic_vector(43, 8),
63790 => conv_std_logic_vector(44, 8),
63791 => conv_std_logic_vector(45, 8),
63792 => conv_std_logic_vector(46, 8),
63793 => conv_std_logic_vector(47, 8),
63794 => conv_std_logic_vector(48, 8),
63795 => conv_std_logic_vector(49, 8),
63796 => conv_std_logic_vector(50, 8),
63797 => conv_std_logic_vector(51, 8),
63798 => conv_std_logic_vector(52, 8),
63799 => conv_std_logic_vector(53, 8),
63800 => conv_std_logic_vector(54, 8),
63801 => conv_std_logic_vector(55, 8),
63802 => conv_std_logic_vector(56, 8),
63803 => conv_std_logic_vector(57, 8),
63804 => conv_std_logic_vector(58, 8),
63805 => conv_std_logic_vector(59, 8),
63806 => conv_std_logic_vector(60, 8),
63807 => conv_std_logic_vector(61, 8),
63808 => conv_std_logic_vector(62, 8),
63809 => conv_std_logic_vector(63, 8),
63810 => conv_std_logic_vector(64, 8),
63811 => conv_std_logic_vector(65, 8),
63812 => conv_std_logic_vector(66, 8),
63813 => conv_std_logic_vector(67, 8),
63814 => conv_std_logic_vector(68, 8),
63815 => conv_std_logic_vector(69, 8),
63816 => conv_std_logic_vector(70, 8),
63817 => conv_std_logic_vector(71, 8),
63818 => conv_std_logic_vector(71, 8),
63819 => conv_std_logic_vector(72, 8),
63820 => conv_std_logic_vector(73, 8),
63821 => conv_std_logic_vector(74, 8),
63822 => conv_std_logic_vector(75, 8),
63823 => conv_std_logic_vector(76, 8),
63824 => conv_std_logic_vector(77, 8),
63825 => conv_std_logic_vector(78, 8),
63826 => conv_std_logic_vector(79, 8),
63827 => conv_std_logic_vector(80, 8),
63828 => conv_std_logic_vector(81, 8),
63829 => conv_std_logic_vector(82, 8),
63830 => conv_std_logic_vector(83, 8),
63831 => conv_std_logic_vector(84, 8),
63832 => conv_std_logic_vector(85, 8),
63833 => conv_std_logic_vector(86, 8),
63834 => conv_std_logic_vector(87, 8),
63835 => conv_std_logic_vector(88, 8),
63836 => conv_std_logic_vector(89, 8),
63837 => conv_std_logic_vector(90, 8),
63838 => conv_std_logic_vector(91, 8),
63839 => conv_std_logic_vector(92, 8),
63840 => conv_std_logic_vector(93, 8),
63841 => conv_std_logic_vector(94, 8),
63842 => conv_std_logic_vector(95, 8),
63843 => conv_std_logic_vector(96, 8),
63844 => conv_std_logic_vector(97, 8),
63845 => conv_std_logic_vector(98, 8),
63846 => conv_std_logic_vector(99, 8),
63847 => conv_std_logic_vector(100, 8),
63848 => conv_std_logic_vector(101, 8),
63849 => conv_std_logic_vector(102, 8),
63850 => conv_std_logic_vector(103, 8),
63851 => conv_std_logic_vector(104, 8),
63852 => conv_std_logic_vector(105, 8),
63853 => conv_std_logic_vector(106, 8),
63854 => conv_std_logic_vector(106, 8),
63855 => conv_std_logic_vector(107, 8),
63856 => conv_std_logic_vector(108, 8),
63857 => conv_std_logic_vector(109, 8),
63858 => conv_std_logic_vector(110, 8),
63859 => conv_std_logic_vector(111, 8),
63860 => conv_std_logic_vector(112, 8),
63861 => conv_std_logic_vector(113, 8),
63862 => conv_std_logic_vector(114, 8),
63863 => conv_std_logic_vector(115, 8),
63864 => conv_std_logic_vector(116, 8),
63865 => conv_std_logic_vector(117, 8),
63866 => conv_std_logic_vector(118, 8),
63867 => conv_std_logic_vector(119, 8),
63868 => conv_std_logic_vector(120, 8),
63869 => conv_std_logic_vector(121, 8),
63870 => conv_std_logic_vector(122, 8),
63871 => conv_std_logic_vector(123, 8),
63872 => conv_std_logic_vector(124, 8),
63873 => conv_std_logic_vector(125, 8),
63874 => conv_std_logic_vector(126, 8),
63875 => conv_std_logic_vector(127, 8),
63876 => conv_std_logic_vector(128, 8),
63877 => conv_std_logic_vector(129, 8),
63878 => conv_std_logic_vector(130, 8),
63879 => conv_std_logic_vector(131, 8),
63880 => conv_std_logic_vector(132, 8),
63881 => conv_std_logic_vector(133, 8),
63882 => conv_std_logic_vector(134, 8),
63883 => conv_std_logic_vector(135, 8),
63884 => conv_std_logic_vector(136, 8),
63885 => conv_std_logic_vector(137, 8),
63886 => conv_std_logic_vector(138, 8),
63887 => conv_std_logic_vector(139, 8),
63888 => conv_std_logic_vector(140, 8),
63889 => conv_std_logic_vector(141, 8),
63890 => conv_std_logic_vector(142, 8),
63891 => conv_std_logic_vector(142, 8),
63892 => conv_std_logic_vector(143, 8),
63893 => conv_std_logic_vector(144, 8),
63894 => conv_std_logic_vector(145, 8),
63895 => conv_std_logic_vector(146, 8),
63896 => conv_std_logic_vector(147, 8),
63897 => conv_std_logic_vector(148, 8),
63898 => conv_std_logic_vector(149, 8),
63899 => conv_std_logic_vector(150, 8),
63900 => conv_std_logic_vector(151, 8),
63901 => conv_std_logic_vector(152, 8),
63902 => conv_std_logic_vector(153, 8),
63903 => conv_std_logic_vector(154, 8),
63904 => conv_std_logic_vector(155, 8),
63905 => conv_std_logic_vector(156, 8),
63906 => conv_std_logic_vector(157, 8),
63907 => conv_std_logic_vector(158, 8),
63908 => conv_std_logic_vector(159, 8),
63909 => conv_std_logic_vector(160, 8),
63910 => conv_std_logic_vector(161, 8),
63911 => conv_std_logic_vector(162, 8),
63912 => conv_std_logic_vector(163, 8),
63913 => conv_std_logic_vector(164, 8),
63914 => conv_std_logic_vector(165, 8),
63915 => conv_std_logic_vector(166, 8),
63916 => conv_std_logic_vector(167, 8),
63917 => conv_std_logic_vector(168, 8),
63918 => conv_std_logic_vector(169, 8),
63919 => conv_std_logic_vector(170, 8),
63920 => conv_std_logic_vector(171, 8),
63921 => conv_std_logic_vector(172, 8),
63922 => conv_std_logic_vector(173, 8),
63923 => conv_std_logic_vector(174, 8),
63924 => conv_std_logic_vector(175, 8),
63925 => conv_std_logic_vector(176, 8),
63926 => conv_std_logic_vector(177, 8),
63927 => conv_std_logic_vector(177, 8),
63928 => conv_std_logic_vector(178, 8),
63929 => conv_std_logic_vector(179, 8),
63930 => conv_std_logic_vector(180, 8),
63931 => conv_std_logic_vector(181, 8),
63932 => conv_std_logic_vector(182, 8),
63933 => conv_std_logic_vector(183, 8),
63934 => conv_std_logic_vector(184, 8),
63935 => conv_std_logic_vector(185, 8),
63936 => conv_std_logic_vector(186, 8),
63937 => conv_std_logic_vector(187, 8),
63938 => conv_std_logic_vector(188, 8),
63939 => conv_std_logic_vector(189, 8),
63940 => conv_std_logic_vector(190, 8),
63941 => conv_std_logic_vector(191, 8),
63942 => conv_std_logic_vector(192, 8),
63943 => conv_std_logic_vector(193, 8),
63944 => conv_std_logic_vector(194, 8),
63945 => conv_std_logic_vector(195, 8),
63946 => conv_std_logic_vector(196, 8),
63947 => conv_std_logic_vector(197, 8),
63948 => conv_std_logic_vector(198, 8),
63949 => conv_std_logic_vector(199, 8),
63950 => conv_std_logic_vector(200, 8),
63951 => conv_std_logic_vector(201, 8),
63952 => conv_std_logic_vector(202, 8),
63953 => conv_std_logic_vector(203, 8),
63954 => conv_std_logic_vector(204, 8),
63955 => conv_std_logic_vector(205, 8),
63956 => conv_std_logic_vector(206, 8),
63957 => conv_std_logic_vector(207, 8),
63958 => conv_std_logic_vector(208, 8),
63959 => conv_std_logic_vector(209, 8),
63960 => conv_std_logic_vector(210, 8),
63961 => conv_std_logic_vector(211, 8),
63962 => conv_std_logic_vector(212, 8),
63963 => conv_std_logic_vector(213, 8),
63964 => conv_std_logic_vector(213, 8),
63965 => conv_std_logic_vector(214, 8),
63966 => conv_std_logic_vector(215, 8),
63967 => conv_std_logic_vector(216, 8),
63968 => conv_std_logic_vector(217, 8),
63969 => conv_std_logic_vector(218, 8),
63970 => conv_std_logic_vector(219, 8),
63971 => conv_std_logic_vector(220, 8),
63972 => conv_std_logic_vector(221, 8),
63973 => conv_std_logic_vector(222, 8),
63974 => conv_std_logic_vector(223, 8),
63975 => conv_std_logic_vector(224, 8),
63976 => conv_std_logic_vector(225, 8),
63977 => conv_std_logic_vector(226, 8),
63978 => conv_std_logic_vector(227, 8),
63979 => conv_std_logic_vector(228, 8),
63980 => conv_std_logic_vector(229, 8),
63981 => conv_std_logic_vector(230, 8),
63982 => conv_std_logic_vector(231, 8),
63983 => conv_std_logic_vector(232, 8),
63984 => conv_std_logic_vector(233, 8),
63985 => conv_std_logic_vector(234, 8),
63986 => conv_std_logic_vector(235, 8),
63987 => conv_std_logic_vector(236, 8),
63988 => conv_std_logic_vector(237, 8),
63989 => conv_std_logic_vector(238, 8),
63990 => conv_std_logic_vector(239, 8),
63991 => conv_std_logic_vector(240, 8),
63992 => conv_std_logic_vector(241, 8),
63993 => conv_std_logic_vector(242, 8),
63994 => conv_std_logic_vector(243, 8),
63995 => conv_std_logic_vector(244, 8),
63996 => conv_std_logic_vector(245, 8),
63997 => conv_std_logic_vector(246, 8),
63998 => conv_std_logic_vector(247, 8),
63999 => conv_std_logic_vector(248, 8),
64000 => conv_std_logic_vector(0, 8),
64001 => conv_std_logic_vector(0, 8),
64002 => conv_std_logic_vector(1, 8),
64003 => conv_std_logic_vector(2, 8),
64004 => conv_std_logic_vector(3, 8),
64005 => conv_std_logic_vector(4, 8),
64006 => conv_std_logic_vector(5, 8),
64007 => conv_std_logic_vector(6, 8),
64008 => conv_std_logic_vector(7, 8),
64009 => conv_std_logic_vector(8, 8),
64010 => conv_std_logic_vector(9, 8),
64011 => conv_std_logic_vector(10, 8),
64012 => conv_std_logic_vector(11, 8),
64013 => conv_std_logic_vector(12, 8),
64014 => conv_std_logic_vector(13, 8),
64015 => conv_std_logic_vector(14, 8),
64016 => conv_std_logic_vector(15, 8),
64017 => conv_std_logic_vector(16, 8),
64018 => conv_std_logic_vector(17, 8),
64019 => conv_std_logic_vector(18, 8),
64020 => conv_std_logic_vector(19, 8),
64021 => conv_std_logic_vector(20, 8),
64022 => conv_std_logic_vector(21, 8),
64023 => conv_std_logic_vector(22, 8),
64024 => conv_std_logic_vector(23, 8),
64025 => conv_std_logic_vector(24, 8),
64026 => conv_std_logic_vector(25, 8),
64027 => conv_std_logic_vector(26, 8),
64028 => conv_std_logic_vector(27, 8),
64029 => conv_std_logic_vector(28, 8),
64030 => conv_std_logic_vector(29, 8),
64031 => conv_std_logic_vector(30, 8),
64032 => conv_std_logic_vector(31, 8),
64033 => conv_std_logic_vector(32, 8),
64034 => conv_std_logic_vector(33, 8),
64035 => conv_std_logic_vector(34, 8),
64036 => conv_std_logic_vector(35, 8),
64037 => conv_std_logic_vector(36, 8),
64038 => conv_std_logic_vector(37, 8),
64039 => conv_std_logic_vector(38, 8),
64040 => conv_std_logic_vector(39, 8),
64041 => conv_std_logic_vector(40, 8),
64042 => conv_std_logic_vector(41, 8),
64043 => conv_std_logic_vector(41, 8),
64044 => conv_std_logic_vector(42, 8),
64045 => conv_std_logic_vector(43, 8),
64046 => conv_std_logic_vector(44, 8),
64047 => conv_std_logic_vector(45, 8),
64048 => conv_std_logic_vector(46, 8),
64049 => conv_std_logic_vector(47, 8),
64050 => conv_std_logic_vector(48, 8),
64051 => conv_std_logic_vector(49, 8),
64052 => conv_std_logic_vector(50, 8),
64053 => conv_std_logic_vector(51, 8),
64054 => conv_std_logic_vector(52, 8),
64055 => conv_std_logic_vector(53, 8),
64056 => conv_std_logic_vector(54, 8),
64057 => conv_std_logic_vector(55, 8),
64058 => conv_std_logic_vector(56, 8),
64059 => conv_std_logic_vector(57, 8),
64060 => conv_std_logic_vector(58, 8),
64061 => conv_std_logic_vector(59, 8),
64062 => conv_std_logic_vector(60, 8),
64063 => conv_std_logic_vector(61, 8),
64064 => conv_std_logic_vector(62, 8),
64065 => conv_std_logic_vector(63, 8),
64066 => conv_std_logic_vector(64, 8),
64067 => conv_std_logic_vector(65, 8),
64068 => conv_std_logic_vector(66, 8),
64069 => conv_std_logic_vector(67, 8),
64070 => conv_std_logic_vector(68, 8),
64071 => conv_std_logic_vector(69, 8),
64072 => conv_std_logic_vector(70, 8),
64073 => conv_std_logic_vector(71, 8),
64074 => conv_std_logic_vector(72, 8),
64075 => conv_std_logic_vector(73, 8),
64076 => conv_std_logic_vector(74, 8),
64077 => conv_std_logic_vector(75, 8),
64078 => conv_std_logic_vector(76, 8),
64079 => conv_std_logic_vector(77, 8),
64080 => conv_std_logic_vector(78, 8),
64081 => conv_std_logic_vector(79, 8),
64082 => conv_std_logic_vector(80, 8),
64083 => conv_std_logic_vector(81, 8),
64084 => conv_std_logic_vector(82, 8),
64085 => conv_std_logic_vector(83, 8),
64086 => conv_std_logic_vector(83, 8),
64087 => conv_std_logic_vector(84, 8),
64088 => conv_std_logic_vector(85, 8),
64089 => conv_std_logic_vector(86, 8),
64090 => conv_std_logic_vector(87, 8),
64091 => conv_std_logic_vector(88, 8),
64092 => conv_std_logic_vector(89, 8),
64093 => conv_std_logic_vector(90, 8),
64094 => conv_std_logic_vector(91, 8),
64095 => conv_std_logic_vector(92, 8),
64096 => conv_std_logic_vector(93, 8),
64097 => conv_std_logic_vector(94, 8),
64098 => conv_std_logic_vector(95, 8),
64099 => conv_std_logic_vector(96, 8),
64100 => conv_std_logic_vector(97, 8),
64101 => conv_std_logic_vector(98, 8),
64102 => conv_std_logic_vector(99, 8),
64103 => conv_std_logic_vector(100, 8),
64104 => conv_std_logic_vector(101, 8),
64105 => conv_std_logic_vector(102, 8),
64106 => conv_std_logic_vector(103, 8),
64107 => conv_std_logic_vector(104, 8),
64108 => conv_std_logic_vector(105, 8),
64109 => conv_std_logic_vector(106, 8),
64110 => conv_std_logic_vector(107, 8),
64111 => conv_std_logic_vector(108, 8),
64112 => conv_std_logic_vector(109, 8),
64113 => conv_std_logic_vector(110, 8),
64114 => conv_std_logic_vector(111, 8),
64115 => conv_std_logic_vector(112, 8),
64116 => conv_std_logic_vector(113, 8),
64117 => conv_std_logic_vector(114, 8),
64118 => conv_std_logic_vector(115, 8),
64119 => conv_std_logic_vector(116, 8),
64120 => conv_std_logic_vector(117, 8),
64121 => conv_std_logic_vector(118, 8),
64122 => conv_std_logic_vector(119, 8),
64123 => conv_std_logic_vector(120, 8),
64124 => conv_std_logic_vector(121, 8),
64125 => conv_std_logic_vector(122, 8),
64126 => conv_std_logic_vector(123, 8),
64127 => conv_std_logic_vector(124, 8),
64128 => conv_std_logic_vector(125, 8),
64129 => conv_std_logic_vector(125, 8),
64130 => conv_std_logic_vector(126, 8),
64131 => conv_std_logic_vector(127, 8),
64132 => conv_std_logic_vector(128, 8),
64133 => conv_std_logic_vector(129, 8),
64134 => conv_std_logic_vector(130, 8),
64135 => conv_std_logic_vector(131, 8),
64136 => conv_std_logic_vector(132, 8),
64137 => conv_std_logic_vector(133, 8),
64138 => conv_std_logic_vector(134, 8),
64139 => conv_std_logic_vector(135, 8),
64140 => conv_std_logic_vector(136, 8),
64141 => conv_std_logic_vector(137, 8),
64142 => conv_std_logic_vector(138, 8),
64143 => conv_std_logic_vector(139, 8),
64144 => conv_std_logic_vector(140, 8),
64145 => conv_std_logic_vector(141, 8),
64146 => conv_std_logic_vector(142, 8),
64147 => conv_std_logic_vector(143, 8),
64148 => conv_std_logic_vector(144, 8),
64149 => conv_std_logic_vector(145, 8),
64150 => conv_std_logic_vector(146, 8),
64151 => conv_std_logic_vector(147, 8),
64152 => conv_std_logic_vector(148, 8),
64153 => conv_std_logic_vector(149, 8),
64154 => conv_std_logic_vector(150, 8),
64155 => conv_std_logic_vector(151, 8),
64156 => conv_std_logic_vector(152, 8),
64157 => conv_std_logic_vector(153, 8),
64158 => conv_std_logic_vector(154, 8),
64159 => conv_std_logic_vector(155, 8),
64160 => conv_std_logic_vector(156, 8),
64161 => conv_std_logic_vector(157, 8),
64162 => conv_std_logic_vector(158, 8),
64163 => conv_std_logic_vector(159, 8),
64164 => conv_std_logic_vector(160, 8),
64165 => conv_std_logic_vector(161, 8),
64166 => conv_std_logic_vector(162, 8),
64167 => conv_std_logic_vector(163, 8),
64168 => conv_std_logic_vector(164, 8),
64169 => conv_std_logic_vector(165, 8),
64170 => conv_std_logic_vector(166, 8),
64171 => conv_std_logic_vector(166, 8),
64172 => conv_std_logic_vector(167, 8),
64173 => conv_std_logic_vector(168, 8),
64174 => conv_std_logic_vector(169, 8),
64175 => conv_std_logic_vector(170, 8),
64176 => conv_std_logic_vector(171, 8),
64177 => conv_std_logic_vector(172, 8),
64178 => conv_std_logic_vector(173, 8),
64179 => conv_std_logic_vector(174, 8),
64180 => conv_std_logic_vector(175, 8),
64181 => conv_std_logic_vector(176, 8),
64182 => conv_std_logic_vector(177, 8),
64183 => conv_std_logic_vector(178, 8),
64184 => conv_std_logic_vector(179, 8),
64185 => conv_std_logic_vector(180, 8),
64186 => conv_std_logic_vector(181, 8),
64187 => conv_std_logic_vector(182, 8),
64188 => conv_std_logic_vector(183, 8),
64189 => conv_std_logic_vector(184, 8),
64190 => conv_std_logic_vector(185, 8),
64191 => conv_std_logic_vector(186, 8),
64192 => conv_std_logic_vector(187, 8),
64193 => conv_std_logic_vector(188, 8),
64194 => conv_std_logic_vector(189, 8),
64195 => conv_std_logic_vector(190, 8),
64196 => conv_std_logic_vector(191, 8),
64197 => conv_std_logic_vector(192, 8),
64198 => conv_std_logic_vector(193, 8),
64199 => conv_std_logic_vector(194, 8),
64200 => conv_std_logic_vector(195, 8),
64201 => conv_std_logic_vector(196, 8),
64202 => conv_std_logic_vector(197, 8),
64203 => conv_std_logic_vector(198, 8),
64204 => conv_std_logic_vector(199, 8),
64205 => conv_std_logic_vector(200, 8),
64206 => conv_std_logic_vector(201, 8),
64207 => conv_std_logic_vector(202, 8),
64208 => conv_std_logic_vector(203, 8),
64209 => conv_std_logic_vector(204, 8),
64210 => conv_std_logic_vector(205, 8),
64211 => conv_std_logic_vector(206, 8),
64212 => conv_std_logic_vector(207, 8),
64213 => conv_std_logic_vector(208, 8),
64214 => conv_std_logic_vector(208, 8),
64215 => conv_std_logic_vector(209, 8),
64216 => conv_std_logic_vector(210, 8),
64217 => conv_std_logic_vector(211, 8),
64218 => conv_std_logic_vector(212, 8),
64219 => conv_std_logic_vector(213, 8),
64220 => conv_std_logic_vector(214, 8),
64221 => conv_std_logic_vector(215, 8),
64222 => conv_std_logic_vector(216, 8),
64223 => conv_std_logic_vector(217, 8),
64224 => conv_std_logic_vector(218, 8),
64225 => conv_std_logic_vector(219, 8),
64226 => conv_std_logic_vector(220, 8),
64227 => conv_std_logic_vector(221, 8),
64228 => conv_std_logic_vector(222, 8),
64229 => conv_std_logic_vector(223, 8),
64230 => conv_std_logic_vector(224, 8),
64231 => conv_std_logic_vector(225, 8),
64232 => conv_std_logic_vector(226, 8),
64233 => conv_std_logic_vector(227, 8),
64234 => conv_std_logic_vector(228, 8),
64235 => conv_std_logic_vector(229, 8),
64236 => conv_std_logic_vector(230, 8),
64237 => conv_std_logic_vector(231, 8),
64238 => conv_std_logic_vector(232, 8),
64239 => conv_std_logic_vector(233, 8),
64240 => conv_std_logic_vector(234, 8),
64241 => conv_std_logic_vector(235, 8),
64242 => conv_std_logic_vector(236, 8),
64243 => conv_std_logic_vector(237, 8),
64244 => conv_std_logic_vector(238, 8),
64245 => conv_std_logic_vector(239, 8),
64246 => conv_std_logic_vector(240, 8),
64247 => conv_std_logic_vector(241, 8),
64248 => conv_std_logic_vector(242, 8),
64249 => conv_std_logic_vector(243, 8),
64250 => conv_std_logic_vector(244, 8),
64251 => conv_std_logic_vector(245, 8),
64252 => conv_std_logic_vector(246, 8),
64253 => conv_std_logic_vector(247, 8),
64254 => conv_std_logic_vector(248, 8),
64255 => conv_std_logic_vector(249, 8),
64256 => conv_std_logic_vector(0, 8),
64257 => conv_std_logic_vector(0, 8),
64258 => conv_std_logic_vector(1, 8),
64259 => conv_std_logic_vector(2, 8),
64260 => conv_std_logic_vector(3, 8),
64261 => conv_std_logic_vector(4, 8),
64262 => conv_std_logic_vector(5, 8),
64263 => conv_std_logic_vector(6, 8),
64264 => conv_std_logic_vector(7, 8),
64265 => conv_std_logic_vector(8, 8),
64266 => conv_std_logic_vector(9, 8),
64267 => conv_std_logic_vector(10, 8),
64268 => conv_std_logic_vector(11, 8),
64269 => conv_std_logic_vector(12, 8),
64270 => conv_std_logic_vector(13, 8),
64271 => conv_std_logic_vector(14, 8),
64272 => conv_std_logic_vector(15, 8),
64273 => conv_std_logic_vector(16, 8),
64274 => conv_std_logic_vector(17, 8),
64275 => conv_std_logic_vector(18, 8),
64276 => conv_std_logic_vector(19, 8),
64277 => conv_std_logic_vector(20, 8),
64278 => conv_std_logic_vector(21, 8),
64279 => conv_std_logic_vector(22, 8),
64280 => conv_std_logic_vector(23, 8),
64281 => conv_std_logic_vector(24, 8),
64282 => conv_std_logic_vector(25, 8),
64283 => conv_std_logic_vector(26, 8),
64284 => conv_std_logic_vector(27, 8),
64285 => conv_std_logic_vector(28, 8),
64286 => conv_std_logic_vector(29, 8),
64287 => conv_std_logic_vector(30, 8),
64288 => conv_std_logic_vector(31, 8),
64289 => conv_std_logic_vector(32, 8),
64290 => conv_std_logic_vector(33, 8),
64291 => conv_std_logic_vector(34, 8),
64292 => conv_std_logic_vector(35, 8),
64293 => conv_std_logic_vector(36, 8),
64294 => conv_std_logic_vector(37, 8),
64295 => conv_std_logic_vector(38, 8),
64296 => conv_std_logic_vector(39, 8),
64297 => conv_std_logic_vector(40, 8),
64298 => conv_std_logic_vector(41, 8),
64299 => conv_std_logic_vector(42, 8),
64300 => conv_std_logic_vector(43, 8),
64301 => conv_std_logic_vector(44, 8),
64302 => conv_std_logic_vector(45, 8),
64303 => conv_std_logic_vector(46, 8),
64304 => conv_std_logic_vector(47, 8),
64305 => conv_std_logic_vector(48, 8),
64306 => conv_std_logic_vector(49, 8),
64307 => conv_std_logic_vector(50, 8),
64308 => conv_std_logic_vector(50, 8),
64309 => conv_std_logic_vector(51, 8),
64310 => conv_std_logic_vector(52, 8),
64311 => conv_std_logic_vector(53, 8),
64312 => conv_std_logic_vector(54, 8),
64313 => conv_std_logic_vector(55, 8),
64314 => conv_std_logic_vector(56, 8),
64315 => conv_std_logic_vector(57, 8),
64316 => conv_std_logic_vector(58, 8),
64317 => conv_std_logic_vector(59, 8),
64318 => conv_std_logic_vector(60, 8),
64319 => conv_std_logic_vector(61, 8),
64320 => conv_std_logic_vector(62, 8),
64321 => conv_std_logic_vector(63, 8),
64322 => conv_std_logic_vector(64, 8),
64323 => conv_std_logic_vector(65, 8),
64324 => conv_std_logic_vector(66, 8),
64325 => conv_std_logic_vector(67, 8),
64326 => conv_std_logic_vector(68, 8),
64327 => conv_std_logic_vector(69, 8),
64328 => conv_std_logic_vector(70, 8),
64329 => conv_std_logic_vector(71, 8),
64330 => conv_std_logic_vector(72, 8),
64331 => conv_std_logic_vector(73, 8),
64332 => conv_std_logic_vector(74, 8),
64333 => conv_std_logic_vector(75, 8),
64334 => conv_std_logic_vector(76, 8),
64335 => conv_std_logic_vector(77, 8),
64336 => conv_std_logic_vector(78, 8),
64337 => conv_std_logic_vector(79, 8),
64338 => conv_std_logic_vector(80, 8),
64339 => conv_std_logic_vector(81, 8),
64340 => conv_std_logic_vector(82, 8),
64341 => conv_std_logic_vector(83, 8),
64342 => conv_std_logic_vector(84, 8),
64343 => conv_std_logic_vector(85, 8),
64344 => conv_std_logic_vector(86, 8),
64345 => conv_std_logic_vector(87, 8),
64346 => conv_std_logic_vector(88, 8),
64347 => conv_std_logic_vector(89, 8),
64348 => conv_std_logic_vector(90, 8),
64349 => conv_std_logic_vector(91, 8),
64350 => conv_std_logic_vector(92, 8),
64351 => conv_std_logic_vector(93, 8),
64352 => conv_std_logic_vector(94, 8),
64353 => conv_std_logic_vector(95, 8),
64354 => conv_std_logic_vector(96, 8),
64355 => conv_std_logic_vector(97, 8),
64356 => conv_std_logic_vector(98, 8),
64357 => conv_std_logic_vector(99, 8),
64358 => conv_std_logic_vector(100, 8),
64359 => conv_std_logic_vector(100, 8),
64360 => conv_std_logic_vector(101, 8),
64361 => conv_std_logic_vector(102, 8),
64362 => conv_std_logic_vector(103, 8),
64363 => conv_std_logic_vector(104, 8),
64364 => conv_std_logic_vector(105, 8),
64365 => conv_std_logic_vector(106, 8),
64366 => conv_std_logic_vector(107, 8),
64367 => conv_std_logic_vector(108, 8),
64368 => conv_std_logic_vector(109, 8),
64369 => conv_std_logic_vector(110, 8),
64370 => conv_std_logic_vector(111, 8),
64371 => conv_std_logic_vector(112, 8),
64372 => conv_std_logic_vector(113, 8),
64373 => conv_std_logic_vector(114, 8),
64374 => conv_std_logic_vector(115, 8),
64375 => conv_std_logic_vector(116, 8),
64376 => conv_std_logic_vector(117, 8),
64377 => conv_std_logic_vector(118, 8),
64378 => conv_std_logic_vector(119, 8),
64379 => conv_std_logic_vector(120, 8),
64380 => conv_std_logic_vector(121, 8),
64381 => conv_std_logic_vector(122, 8),
64382 => conv_std_logic_vector(123, 8),
64383 => conv_std_logic_vector(124, 8),
64384 => conv_std_logic_vector(125, 8),
64385 => conv_std_logic_vector(126, 8),
64386 => conv_std_logic_vector(127, 8),
64387 => conv_std_logic_vector(128, 8),
64388 => conv_std_logic_vector(129, 8),
64389 => conv_std_logic_vector(130, 8),
64390 => conv_std_logic_vector(131, 8),
64391 => conv_std_logic_vector(132, 8),
64392 => conv_std_logic_vector(133, 8),
64393 => conv_std_logic_vector(134, 8),
64394 => conv_std_logic_vector(135, 8),
64395 => conv_std_logic_vector(136, 8),
64396 => conv_std_logic_vector(137, 8),
64397 => conv_std_logic_vector(138, 8),
64398 => conv_std_logic_vector(139, 8),
64399 => conv_std_logic_vector(140, 8),
64400 => conv_std_logic_vector(141, 8),
64401 => conv_std_logic_vector(142, 8),
64402 => conv_std_logic_vector(143, 8),
64403 => conv_std_logic_vector(144, 8),
64404 => conv_std_logic_vector(145, 8),
64405 => conv_std_logic_vector(146, 8),
64406 => conv_std_logic_vector(147, 8),
64407 => conv_std_logic_vector(148, 8),
64408 => conv_std_logic_vector(149, 8),
64409 => conv_std_logic_vector(150, 8),
64410 => conv_std_logic_vector(150, 8),
64411 => conv_std_logic_vector(151, 8),
64412 => conv_std_logic_vector(152, 8),
64413 => conv_std_logic_vector(153, 8),
64414 => conv_std_logic_vector(154, 8),
64415 => conv_std_logic_vector(155, 8),
64416 => conv_std_logic_vector(156, 8),
64417 => conv_std_logic_vector(157, 8),
64418 => conv_std_logic_vector(158, 8),
64419 => conv_std_logic_vector(159, 8),
64420 => conv_std_logic_vector(160, 8),
64421 => conv_std_logic_vector(161, 8),
64422 => conv_std_logic_vector(162, 8),
64423 => conv_std_logic_vector(163, 8),
64424 => conv_std_logic_vector(164, 8),
64425 => conv_std_logic_vector(165, 8),
64426 => conv_std_logic_vector(166, 8),
64427 => conv_std_logic_vector(167, 8),
64428 => conv_std_logic_vector(168, 8),
64429 => conv_std_logic_vector(169, 8),
64430 => conv_std_logic_vector(170, 8),
64431 => conv_std_logic_vector(171, 8),
64432 => conv_std_logic_vector(172, 8),
64433 => conv_std_logic_vector(173, 8),
64434 => conv_std_logic_vector(174, 8),
64435 => conv_std_logic_vector(175, 8),
64436 => conv_std_logic_vector(176, 8),
64437 => conv_std_logic_vector(177, 8),
64438 => conv_std_logic_vector(178, 8),
64439 => conv_std_logic_vector(179, 8),
64440 => conv_std_logic_vector(180, 8),
64441 => conv_std_logic_vector(181, 8),
64442 => conv_std_logic_vector(182, 8),
64443 => conv_std_logic_vector(183, 8),
64444 => conv_std_logic_vector(184, 8),
64445 => conv_std_logic_vector(185, 8),
64446 => conv_std_logic_vector(186, 8),
64447 => conv_std_logic_vector(187, 8),
64448 => conv_std_logic_vector(188, 8),
64449 => conv_std_logic_vector(189, 8),
64450 => conv_std_logic_vector(190, 8),
64451 => conv_std_logic_vector(191, 8),
64452 => conv_std_logic_vector(192, 8),
64453 => conv_std_logic_vector(193, 8),
64454 => conv_std_logic_vector(194, 8),
64455 => conv_std_logic_vector(195, 8),
64456 => conv_std_logic_vector(196, 8),
64457 => conv_std_logic_vector(197, 8),
64458 => conv_std_logic_vector(198, 8),
64459 => conv_std_logic_vector(199, 8),
64460 => conv_std_logic_vector(200, 8),
64461 => conv_std_logic_vector(200, 8),
64462 => conv_std_logic_vector(201, 8),
64463 => conv_std_logic_vector(202, 8),
64464 => conv_std_logic_vector(203, 8),
64465 => conv_std_logic_vector(204, 8),
64466 => conv_std_logic_vector(205, 8),
64467 => conv_std_logic_vector(206, 8),
64468 => conv_std_logic_vector(207, 8),
64469 => conv_std_logic_vector(208, 8),
64470 => conv_std_logic_vector(209, 8),
64471 => conv_std_logic_vector(210, 8),
64472 => conv_std_logic_vector(211, 8),
64473 => conv_std_logic_vector(212, 8),
64474 => conv_std_logic_vector(213, 8),
64475 => conv_std_logic_vector(214, 8),
64476 => conv_std_logic_vector(215, 8),
64477 => conv_std_logic_vector(216, 8),
64478 => conv_std_logic_vector(217, 8),
64479 => conv_std_logic_vector(218, 8),
64480 => conv_std_logic_vector(219, 8),
64481 => conv_std_logic_vector(220, 8),
64482 => conv_std_logic_vector(221, 8),
64483 => conv_std_logic_vector(222, 8),
64484 => conv_std_logic_vector(223, 8),
64485 => conv_std_logic_vector(224, 8),
64486 => conv_std_logic_vector(225, 8),
64487 => conv_std_logic_vector(226, 8),
64488 => conv_std_logic_vector(227, 8),
64489 => conv_std_logic_vector(228, 8),
64490 => conv_std_logic_vector(229, 8),
64491 => conv_std_logic_vector(230, 8),
64492 => conv_std_logic_vector(231, 8),
64493 => conv_std_logic_vector(232, 8),
64494 => conv_std_logic_vector(233, 8),
64495 => conv_std_logic_vector(234, 8),
64496 => conv_std_logic_vector(235, 8),
64497 => conv_std_logic_vector(236, 8),
64498 => conv_std_logic_vector(237, 8),
64499 => conv_std_logic_vector(238, 8),
64500 => conv_std_logic_vector(239, 8),
64501 => conv_std_logic_vector(240, 8),
64502 => conv_std_logic_vector(241, 8),
64503 => conv_std_logic_vector(242, 8),
64504 => conv_std_logic_vector(243, 8),
64505 => conv_std_logic_vector(244, 8),
64506 => conv_std_logic_vector(245, 8),
64507 => conv_std_logic_vector(246, 8),
64508 => conv_std_logic_vector(247, 8),
64509 => conv_std_logic_vector(248, 8),
64510 => conv_std_logic_vector(249, 8),
64511 => conv_std_logic_vector(250, 8),
64512 => conv_std_logic_vector(0, 8),
64513 => conv_std_logic_vector(0, 8),
64514 => conv_std_logic_vector(1, 8),
64515 => conv_std_logic_vector(2, 8),
64516 => conv_std_logic_vector(3, 8),
64517 => conv_std_logic_vector(4, 8),
64518 => conv_std_logic_vector(5, 8),
64519 => conv_std_logic_vector(6, 8),
64520 => conv_std_logic_vector(7, 8),
64521 => conv_std_logic_vector(8, 8),
64522 => conv_std_logic_vector(9, 8),
64523 => conv_std_logic_vector(10, 8),
64524 => conv_std_logic_vector(11, 8),
64525 => conv_std_logic_vector(12, 8),
64526 => conv_std_logic_vector(13, 8),
64527 => conv_std_logic_vector(14, 8),
64528 => conv_std_logic_vector(15, 8),
64529 => conv_std_logic_vector(16, 8),
64530 => conv_std_logic_vector(17, 8),
64531 => conv_std_logic_vector(18, 8),
64532 => conv_std_logic_vector(19, 8),
64533 => conv_std_logic_vector(20, 8),
64534 => conv_std_logic_vector(21, 8),
64535 => conv_std_logic_vector(22, 8),
64536 => conv_std_logic_vector(23, 8),
64537 => conv_std_logic_vector(24, 8),
64538 => conv_std_logic_vector(25, 8),
64539 => conv_std_logic_vector(26, 8),
64540 => conv_std_logic_vector(27, 8),
64541 => conv_std_logic_vector(28, 8),
64542 => conv_std_logic_vector(29, 8),
64543 => conv_std_logic_vector(30, 8),
64544 => conv_std_logic_vector(31, 8),
64545 => conv_std_logic_vector(32, 8),
64546 => conv_std_logic_vector(33, 8),
64547 => conv_std_logic_vector(34, 8),
64548 => conv_std_logic_vector(35, 8),
64549 => conv_std_logic_vector(36, 8),
64550 => conv_std_logic_vector(37, 8),
64551 => conv_std_logic_vector(38, 8),
64552 => conv_std_logic_vector(39, 8),
64553 => conv_std_logic_vector(40, 8),
64554 => conv_std_logic_vector(41, 8),
64555 => conv_std_logic_vector(42, 8),
64556 => conv_std_logic_vector(43, 8),
64557 => conv_std_logic_vector(44, 8),
64558 => conv_std_logic_vector(45, 8),
64559 => conv_std_logic_vector(46, 8),
64560 => conv_std_logic_vector(47, 8),
64561 => conv_std_logic_vector(48, 8),
64562 => conv_std_logic_vector(49, 8),
64563 => conv_std_logic_vector(50, 8),
64564 => conv_std_logic_vector(51, 8),
64565 => conv_std_logic_vector(52, 8),
64566 => conv_std_logic_vector(53, 8),
64567 => conv_std_logic_vector(54, 8),
64568 => conv_std_logic_vector(55, 8),
64569 => conv_std_logic_vector(56, 8),
64570 => conv_std_logic_vector(57, 8),
64571 => conv_std_logic_vector(58, 8),
64572 => conv_std_logic_vector(59, 8),
64573 => conv_std_logic_vector(60, 8),
64574 => conv_std_logic_vector(61, 8),
64575 => conv_std_logic_vector(62, 8),
64576 => conv_std_logic_vector(63, 8),
64577 => conv_std_logic_vector(63, 8),
64578 => conv_std_logic_vector(64, 8),
64579 => conv_std_logic_vector(65, 8),
64580 => conv_std_logic_vector(66, 8),
64581 => conv_std_logic_vector(67, 8),
64582 => conv_std_logic_vector(68, 8),
64583 => conv_std_logic_vector(69, 8),
64584 => conv_std_logic_vector(70, 8),
64585 => conv_std_logic_vector(71, 8),
64586 => conv_std_logic_vector(72, 8),
64587 => conv_std_logic_vector(73, 8),
64588 => conv_std_logic_vector(74, 8),
64589 => conv_std_logic_vector(75, 8),
64590 => conv_std_logic_vector(76, 8),
64591 => conv_std_logic_vector(77, 8),
64592 => conv_std_logic_vector(78, 8),
64593 => conv_std_logic_vector(79, 8),
64594 => conv_std_logic_vector(80, 8),
64595 => conv_std_logic_vector(81, 8),
64596 => conv_std_logic_vector(82, 8),
64597 => conv_std_logic_vector(83, 8),
64598 => conv_std_logic_vector(84, 8),
64599 => conv_std_logic_vector(85, 8),
64600 => conv_std_logic_vector(86, 8),
64601 => conv_std_logic_vector(87, 8),
64602 => conv_std_logic_vector(88, 8),
64603 => conv_std_logic_vector(89, 8),
64604 => conv_std_logic_vector(90, 8),
64605 => conv_std_logic_vector(91, 8),
64606 => conv_std_logic_vector(92, 8),
64607 => conv_std_logic_vector(93, 8),
64608 => conv_std_logic_vector(94, 8),
64609 => conv_std_logic_vector(95, 8),
64610 => conv_std_logic_vector(96, 8),
64611 => conv_std_logic_vector(97, 8),
64612 => conv_std_logic_vector(98, 8),
64613 => conv_std_logic_vector(99, 8),
64614 => conv_std_logic_vector(100, 8),
64615 => conv_std_logic_vector(101, 8),
64616 => conv_std_logic_vector(102, 8),
64617 => conv_std_logic_vector(103, 8),
64618 => conv_std_logic_vector(104, 8),
64619 => conv_std_logic_vector(105, 8),
64620 => conv_std_logic_vector(106, 8),
64621 => conv_std_logic_vector(107, 8),
64622 => conv_std_logic_vector(108, 8),
64623 => conv_std_logic_vector(109, 8),
64624 => conv_std_logic_vector(110, 8),
64625 => conv_std_logic_vector(111, 8),
64626 => conv_std_logic_vector(112, 8),
64627 => conv_std_logic_vector(113, 8),
64628 => conv_std_logic_vector(114, 8),
64629 => conv_std_logic_vector(115, 8),
64630 => conv_std_logic_vector(116, 8),
64631 => conv_std_logic_vector(117, 8),
64632 => conv_std_logic_vector(118, 8),
64633 => conv_std_logic_vector(119, 8),
64634 => conv_std_logic_vector(120, 8),
64635 => conv_std_logic_vector(121, 8),
64636 => conv_std_logic_vector(122, 8),
64637 => conv_std_logic_vector(123, 8),
64638 => conv_std_logic_vector(124, 8),
64639 => conv_std_logic_vector(125, 8),
64640 => conv_std_logic_vector(126, 8),
64641 => conv_std_logic_vector(126, 8),
64642 => conv_std_logic_vector(127, 8),
64643 => conv_std_logic_vector(128, 8),
64644 => conv_std_logic_vector(129, 8),
64645 => conv_std_logic_vector(130, 8),
64646 => conv_std_logic_vector(131, 8),
64647 => conv_std_logic_vector(132, 8),
64648 => conv_std_logic_vector(133, 8),
64649 => conv_std_logic_vector(134, 8),
64650 => conv_std_logic_vector(135, 8),
64651 => conv_std_logic_vector(136, 8),
64652 => conv_std_logic_vector(137, 8),
64653 => conv_std_logic_vector(138, 8),
64654 => conv_std_logic_vector(139, 8),
64655 => conv_std_logic_vector(140, 8),
64656 => conv_std_logic_vector(141, 8),
64657 => conv_std_logic_vector(142, 8),
64658 => conv_std_logic_vector(143, 8),
64659 => conv_std_logic_vector(144, 8),
64660 => conv_std_logic_vector(145, 8),
64661 => conv_std_logic_vector(146, 8),
64662 => conv_std_logic_vector(147, 8),
64663 => conv_std_logic_vector(148, 8),
64664 => conv_std_logic_vector(149, 8),
64665 => conv_std_logic_vector(150, 8),
64666 => conv_std_logic_vector(151, 8),
64667 => conv_std_logic_vector(152, 8),
64668 => conv_std_logic_vector(153, 8),
64669 => conv_std_logic_vector(154, 8),
64670 => conv_std_logic_vector(155, 8),
64671 => conv_std_logic_vector(156, 8),
64672 => conv_std_logic_vector(157, 8),
64673 => conv_std_logic_vector(158, 8),
64674 => conv_std_logic_vector(159, 8),
64675 => conv_std_logic_vector(160, 8),
64676 => conv_std_logic_vector(161, 8),
64677 => conv_std_logic_vector(162, 8),
64678 => conv_std_logic_vector(163, 8),
64679 => conv_std_logic_vector(164, 8),
64680 => conv_std_logic_vector(165, 8),
64681 => conv_std_logic_vector(166, 8),
64682 => conv_std_logic_vector(167, 8),
64683 => conv_std_logic_vector(168, 8),
64684 => conv_std_logic_vector(169, 8),
64685 => conv_std_logic_vector(170, 8),
64686 => conv_std_logic_vector(171, 8),
64687 => conv_std_logic_vector(172, 8),
64688 => conv_std_logic_vector(173, 8),
64689 => conv_std_logic_vector(174, 8),
64690 => conv_std_logic_vector(175, 8),
64691 => conv_std_logic_vector(176, 8),
64692 => conv_std_logic_vector(177, 8),
64693 => conv_std_logic_vector(178, 8),
64694 => conv_std_logic_vector(179, 8),
64695 => conv_std_logic_vector(180, 8),
64696 => conv_std_logic_vector(181, 8),
64697 => conv_std_logic_vector(182, 8),
64698 => conv_std_logic_vector(183, 8),
64699 => conv_std_logic_vector(184, 8),
64700 => conv_std_logic_vector(185, 8),
64701 => conv_std_logic_vector(186, 8),
64702 => conv_std_logic_vector(187, 8),
64703 => conv_std_logic_vector(188, 8),
64704 => conv_std_logic_vector(189, 8),
64705 => conv_std_logic_vector(189, 8),
64706 => conv_std_logic_vector(190, 8),
64707 => conv_std_logic_vector(191, 8),
64708 => conv_std_logic_vector(192, 8),
64709 => conv_std_logic_vector(193, 8),
64710 => conv_std_logic_vector(194, 8),
64711 => conv_std_logic_vector(195, 8),
64712 => conv_std_logic_vector(196, 8),
64713 => conv_std_logic_vector(197, 8),
64714 => conv_std_logic_vector(198, 8),
64715 => conv_std_logic_vector(199, 8),
64716 => conv_std_logic_vector(200, 8),
64717 => conv_std_logic_vector(201, 8),
64718 => conv_std_logic_vector(202, 8),
64719 => conv_std_logic_vector(203, 8),
64720 => conv_std_logic_vector(204, 8),
64721 => conv_std_logic_vector(205, 8),
64722 => conv_std_logic_vector(206, 8),
64723 => conv_std_logic_vector(207, 8),
64724 => conv_std_logic_vector(208, 8),
64725 => conv_std_logic_vector(209, 8),
64726 => conv_std_logic_vector(210, 8),
64727 => conv_std_logic_vector(211, 8),
64728 => conv_std_logic_vector(212, 8),
64729 => conv_std_logic_vector(213, 8),
64730 => conv_std_logic_vector(214, 8),
64731 => conv_std_logic_vector(215, 8),
64732 => conv_std_logic_vector(216, 8),
64733 => conv_std_logic_vector(217, 8),
64734 => conv_std_logic_vector(218, 8),
64735 => conv_std_logic_vector(219, 8),
64736 => conv_std_logic_vector(220, 8),
64737 => conv_std_logic_vector(221, 8),
64738 => conv_std_logic_vector(222, 8),
64739 => conv_std_logic_vector(223, 8),
64740 => conv_std_logic_vector(224, 8),
64741 => conv_std_logic_vector(225, 8),
64742 => conv_std_logic_vector(226, 8),
64743 => conv_std_logic_vector(227, 8),
64744 => conv_std_logic_vector(228, 8),
64745 => conv_std_logic_vector(229, 8),
64746 => conv_std_logic_vector(230, 8),
64747 => conv_std_logic_vector(231, 8),
64748 => conv_std_logic_vector(232, 8),
64749 => conv_std_logic_vector(233, 8),
64750 => conv_std_logic_vector(234, 8),
64751 => conv_std_logic_vector(235, 8),
64752 => conv_std_logic_vector(236, 8),
64753 => conv_std_logic_vector(237, 8),
64754 => conv_std_logic_vector(238, 8),
64755 => conv_std_logic_vector(239, 8),
64756 => conv_std_logic_vector(240, 8),
64757 => conv_std_logic_vector(241, 8),
64758 => conv_std_logic_vector(242, 8),
64759 => conv_std_logic_vector(243, 8),
64760 => conv_std_logic_vector(244, 8),
64761 => conv_std_logic_vector(245, 8),
64762 => conv_std_logic_vector(246, 8),
64763 => conv_std_logic_vector(247, 8),
64764 => conv_std_logic_vector(248, 8),
64765 => conv_std_logic_vector(249, 8),
64766 => conv_std_logic_vector(250, 8),
64767 => conv_std_logic_vector(251, 8),
64768 => conv_std_logic_vector(0, 8),
64769 => conv_std_logic_vector(0, 8),
64770 => conv_std_logic_vector(1, 8),
64771 => conv_std_logic_vector(2, 8),
64772 => conv_std_logic_vector(3, 8),
64773 => conv_std_logic_vector(4, 8),
64774 => conv_std_logic_vector(5, 8),
64775 => conv_std_logic_vector(6, 8),
64776 => conv_std_logic_vector(7, 8),
64777 => conv_std_logic_vector(8, 8),
64778 => conv_std_logic_vector(9, 8),
64779 => conv_std_logic_vector(10, 8),
64780 => conv_std_logic_vector(11, 8),
64781 => conv_std_logic_vector(12, 8),
64782 => conv_std_logic_vector(13, 8),
64783 => conv_std_logic_vector(14, 8),
64784 => conv_std_logic_vector(15, 8),
64785 => conv_std_logic_vector(16, 8),
64786 => conv_std_logic_vector(17, 8),
64787 => conv_std_logic_vector(18, 8),
64788 => conv_std_logic_vector(19, 8),
64789 => conv_std_logic_vector(20, 8),
64790 => conv_std_logic_vector(21, 8),
64791 => conv_std_logic_vector(22, 8),
64792 => conv_std_logic_vector(23, 8),
64793 => conv_std_logic_vector(24, 8),
64794 => conv_std_logic_vector(25, 8),
64795 => conv_std_logic_vector(26, 8),
64796 => conv_std_logic_vector(27, 8),
64797 => conv_std_logic_vector(28, 8),
64798 => conv_std_logic_vector(29, 8),
64799 => conv_std_logic_vector(30, 8),
64800 => conv_std_logic_vector(31, 8),
64801 => conv_std_logic_vector(32, 8),
64802 => conv_std_logic_vector(33, 8),
64803 => conv_std_logic_vector(34, 8),
64804 => conv_std_logic_vector(35, 8),
64805 => conv_std_logic_vector(36, 8),
64806 => conv_std_logic_vector(37, 8),
64807 => conv_std_logic_vector(38, 8),
64808 => conv_std_logic_vector(39, 8),
64809 => conv_std_logic_vector(40, 8),
64810 => conv_std_logic_vector(41, 8),
64811 => conv_std_logic_vector(42, 8),
64812 => conv_std_logic_vector(43, 8),
64813 => conv_std_logic_vector(44, 8),
64814 => conv_std_logic_vector(45, 8),
64815 => conv_std_logic_vector(46, 8),
64816 => conv_std_logic_vector(47, 8),
64817 => conv_std_logic_vector(48, 8),
64818 => conv_std_logic_vector(49, 8),
64819 => conv_std_logic_vector(50, 8),
64820 => conv_std_logic_vector(51, 8),
64821 => conv_std_logic_vector(52, 8),
64822 => conv_std_logic_vector(53, 8),
64823 => conv_std_logic_vector(54, 8),
64824 => conv_std_logic_vector(55, 8),
64825 => conv_std_logic_vector(56, 8),
64826 => conv_std_logic_vector(57, 8),
64827 => conv_std_logic_vector(58, 8),
64828 => conv_std_logic_vector(59, 8),
64829 => conv_std_logic_vector(60, 8),
64830 => conv_std_logic_vector(61, 8),
64831 => conv_std_logic_vector(62, 8),
64832 => conv_std_logic_vector(63, 8),
64833 => conv_std_logic_vector(64, 8),
64834 => conv_std_logic_vector(65, 8),
64835 => conv_std_logic_vector(66, 8),
64836 => conv_std_logic_vector(67, 8),
64837 => conv_std_logic_vector(68, 8),
64838 => conv_std_logic_vector(69, 8),
64839 => conv_std_logic_vector(70, 8),
64840 => conv_std_logic_vector(71, 8),
64841 => conv_std_logic_vector(72, 8),
64842 => conv_std_logic_vector(73, 8),
64843 => conv_std_logic_vector(74, 8),
64844 => conv_std_logic_vector(75, 8),
64845 => conv_std_logic_vector(76, 8),
64846 => conv_std_logic_vector(77, 8),
64847 => conv_std_logic_vector(78, 8),
64848 => conv_std_logic_vector(79, 8),
64849 => conv_std_logic_vector(80, 8),
64850 => conv_std_logic_vector(81, 8),
64851 => conv_std_logic_vector(82, 8),
64852 => conv_std_logic_vector(83, 8),
64853 => conv_std_logic_vector(84, 8),
64854 => conv_std_logic_vector(84, 8),
64855 => conv_std_logic_vector(85, 8),
64856 => conv_std_logic_vector(86, 8),
64857 => conv_std_logic_vector(87, 8),
64858 => conv_std_logic_vector(88, 8),
64859 => conv_std_logic_vector(89, 8),
64860 => conv_std_logic_vector(90, 8),
64861 => conv_std_logic_vector(91, 8),
64862 => conv_std_logic_vector(92, 8),
64863 => conv_std_logic_vector(93, 8),
64864 => conv_std_logic_vector(94, 8),
64865 => conv_std_logic_vector(95, 8),
64866 => conv_std_logic_vector(96, 8),
64867 => conv_std_logic_vector(97, 8),
64868 => conv_std_logic_vector(98, 8),
64869 => conv_std_logic_vector(99, 8),
64870 => conv_std_logic_vector(100, 8),
64871 => conv_std_logic_vector(101, 8),
64872 => conv_std_logic_vector(102, 8),
64873 => conv_std_logic_vector(103, 8),
64874 => conv_std_logic_vector(104, 8),
64875 => conv_std_logic_vector(105, 8),
64876 => conv_std_logic_vector(106, 8),
64877 => conv_std_logic_vector(107, 8),
64878 => conv_std_logic_vector(108, 8),
64879 => conv_std_logic_vector(109, 8),
64880 => conv_std_logic_vector(110, 8),
64881 => conv_std_logic_vector(111, 8),
64882 => conv_std_logic_vector(112, 8),
64883 => conv_std_logic_vector(113, 8),
64884 => conv_std_logic_vector(114, 8),
64885 => conv_std_logic_vector(115, 8),
64886 => conv_std_logic_vector(116, 8),
64887 => conv_std_logic_vector(117, 8),
64888 => conv_std_logic_vector(118, 8),
64889 => conv_std_logic_vector(119, 8),
64890 => conv_std_logic_vector(120, 8),
64891 => conv_std_logic_vector(121, 8),
64892 => conv_std_logic_vector(122, 8),
64893 => conv_std_logic_vector(123, 8),
64894 => conv_std_logic_vector(124, 8),
64895 => conv_std_logic_vector(125, 8),
64896 => conv_std_logic_vector(126, 8),
64897 => conv_std_logic_vector(127, 8),
64898 => conv_std_logic_vector(128, 8),
64899 => conv_std_logic_vector(129, 8),
64900 => conv_std_logic_vector(130, 8),
64901 => conv_std_logic_vector(131, 8),
64902 => conv_std_logic_vector(132, 8),
64903 => conv_std_logic_vector(133, 8),
64904 => conv_std_logic_vector(134, 8),
64905 => conv_std_logic_vector(135, 8),
64906 => conv_std_logic_vector(136, 8),
64907 => conv_std_logic_vector(137, 8),
64908 => conv_std_logic_vector(138, 8),
64909 => conv_std_logic_vector(139, 8),
64910 => conv_std_logic_vector(140, 8),
64911 => conv_std_logic_vector(141, 8),
64912 => conv_std_logic_vector(142, 8),
64913 => conv_std_logic_vector(143, 8),
64914 => conv_std_logic_vector(144, 8),
64915 => conv_std_logic_vector(145, 8),
64916 => conv_std_logic_vector(146, 8),
64917 => conv_std_logic_vector(147, 8),
64918 => conv_std_logic_vector(148, 8),
64919 => conv_std_logic_vector(149, 8),
64920 => conv_std_logic_vector(150, 8),
64921 => conv_std_logic_vector(151, 8),
64922 => conv_std_logic_vector(152, 8),
64923 => conv_std_logic_vector(153, 8),
64924 => conv_std_logic_vector(154, 8),
64925 => conv_std_logic_vector(155, 8),
64926 => conv_std_logic_vector(156, 8),
64927 => conv_std_logic_vector(157, 8),
64928 => conv_std_logic_vector(158, 8),
64929 => conv_std_logic_vector(159, 8),
64930 => conv_std_logic_vector(160, 8),
64931 => conv_std_logic_vector(161, 8),
64932 => conv_std_logic_vector(162, 8),
64933 => conv_std_logic_vector(163, 8),
64934 => conv_std_logic_vector(164, 8),
64935 => conv_std_logic_vector(165, 8),
64936 => conv_std_logic_vector(166, 8),
64937 => conv_std_logic_vector(167, 8),
64938 => conv_std_logic_vector(168, 8),
64939 => conv_std_logic_vector(168, 8),
64940 => conv_std_logic_vector(169, 8),
64941 => conv_std_logic_vector(170, 8),
64942 => conv_std_logic_vector(171, 8),
64943 => conv_std_logic_vector(172, 8),
64944 => conv_std_logic_vector(173, 8),
64945 => conv_std_logic_vector(174, 8),
64946 => conv_std_logic_vector(175, 8),
64947 => conv_std_logic_vector(176, 8),
64948 => conv_std_logic_vector(177, 8),
64949 => conv_std_logic_vector(178, 8),
64950 => conv_std_logic_vector(179, 8),
64951 => conv_std_logic_vector(180, 8),
64952 => conv_std_logic_vector(181, 8),
64953 => conv_std_logic_vector(182, 8),
64954 => conv_std_logic_vector(183, 8),
64955 => conv_std_logic_vector(184, 8),
64956 => conv_std_logic_vector(185, 8),
64957 => conv_std_logic_vector(186, 8),
64958 => conv_std_logic_vector(187, 8),
64959 => conv_std_logic_vector(188, 8),
64960 => conv_std_logic_vector(189, 8),
64961 => conv_std_logic_vector(190, 8),
64962 => conv_std_logic_vector(191, 8),
64963 => conv_std_logic_vector(192, 8),
64964 => conv_std_logic_vector(193, 8),
64965 => conv_std_logic_vector(194, 8),
64966 => conv_std_logic_vector(195, 8),
64967 => conv_std_logic_vector(196, 8),
64968 => conv_std_logic_vector(197, 8),
64969 => conv_std_logic_vector(198, 8),
64970 => conv_std_logic_vector(199, 8),
64971 => conv_std_logic_vector(200, 8),
64972 => conv_std_logic_vector(201, 8),
64973 => conv_std_logic_vector(202, 8),
64974 => conv_std_logic_vector(203, 8),
64975 => conv_std_logic_vector(204, 8),
64976 => conv_std_logic_vector(205, 8),
64977 => conv_std_logic_vector(206, 8),
64978 => conv_std_logic_vector(207, 8),
64979 => conv_std_logic_vector(208, 8),
64980 => conv_std_logic_vector(209, 8),
64981 => conv_std_logic_vector(210, 8),
64982 => conv_std_logic_vector(211, 8),
64983 => conv_std_logic_vector(212, 8),
64984 => conv_std_logic_vector(213, 8),
64985 => conv_std_logic_vector(214, 8),
64986 => conv_std_logic_vector(215, 8),
64987 => conv_std_logic_vector(216, 8),
64988 => conv_std_logic_vector(217, 8),
64989 => conv_std_logic_vector(218, 8),
64990 => conv_std_logic_vector(219, 8),
64991 => conv_std_logic_vector(220, 8),
64992 => conv_std_logic_vector(221, 8),
64993 => conv_std_logic_vector(222, 8),
64994 => conv_std_logic_vector(223, 8),
64995 => conv_std_logic_vector(224, 8),
64996 => conv_std_logic_vector(225, 8),
64997 => conv_std_logic_vector(226, 8),
64998 => conv_std_logic_vector(227, 8),
64999 => conv_std_logic_vector(228, 8),
65000 => conv_std_logic_vector(229, 8),
65001 => conv_std_logic_vector(230, 8),
65002 => conv_std_logic_vector(231, 8),
65003 => conv_std_logic_vector(232, 8),
65004 => conv_std_logic_vector(233, 8),
65005 => conv_std_logic_vector(234, 8),
65006 => conv_std_logic_vector(235, 8),
65007 => conv_std_logic_vector(236, 8),
65008 => conv_std_logic_vector(237, 8),
65009 => conv_std_logic_vector(238, 8),
65010 => conv_std_logic_vector(239, 8),
65011 => conv_std_logic_vector(240, 8),
65012 => conv_std_logic_vector(241, 8),
65013 => conv_std_logic_vector(242, 8),
65014 => conv_std_logic_vector(243, 8),
65015 => conv_std_logic_vector(244, 8),
65016 => conv_std_logic_vector(245, 8),
65017 => conv_std_logic_vector(246, 8),
65018 => conv_std_logic_vector(247, 8),
65019 => conv_std_logic_vector(248, 8),
65020 => conv_std_logic_vector(249, 8),
65021 => conv_std_logic_vector(250, 8),
65022 => conv_std_logic_vector(251, 8),
65023 => conv_std_logic_vector(252, 8),
65024 => conv_std_logic_vector(0, 8),
65025 => conv_std_logic_vector(0, 8),
65026 => conv_std_logic_vector(1, 8),
65027 => conv_std_logic_vector(2, 8),
65028 => conv_std_logic_vector(3, 8),
65029 => conv_std_logic_vector(4, 8),
65030 => conv_std_logic_vector(5, 8),
65031 => conv_std_logic_vector(6, 8),
65032 => conv_std_logic_vector(7, 8),
65033 => conv_std_logic_vector(8, 8),
65034 => conv_std_logic_vector(9, 8),
65035 => conv_std_logic_vector(10, 8),
65036 => conv_std_logic_vector(11, 8),
65037 => conv_std_logic_vector(12, 8),
65038 => conv_std_logic_vector(13, 8),
65039 => conv_std_logic_vector(14, 8),
65040 => conv_std_logic_vector(15, 8),
65041 => conv_std_logic_vector(16, 8),
65042 => conv_std_logic_vector(17, 8),
65043 => conv_std_logic_vector(18, 8),
65044 => conv_std_logic_vector(19, 8),
65045 => conv_std_logic_vector(20, 8),
65046 => conv_std_logic_vector(21, 8),
65047 => conv_std_logic_vector(22, 8),
65048 => conv_std_logic_vector(23, 8),
65049 => conv_std_logic_vector(24, 8),
65050 => conv_std_logic_vector(25, 8),
65051 => conv_std_logic_vector(26, 8),
65052 => conv_std_logic_vector(27, 8),
65053 => conv_std_logic_vector(28, 8),
65054 => conv_std_logic_vector(29, 8),
65055 => conv_std_logic_vector(30, 8),
65056 => conv_std_logic_vector(31, 8),
65057 => conv_std_logic_vector(32, 8),
65058 => conv_std_logic_vector(33, 8),
65059 => conv_std_logic_vector(34, 8),
65060 => conv_std_logic_vector(35, 8),
65061 => conv_std_logic_vector(36, 8),
65062 => conv_std_logic_vector(37, 8),
65063 => conv_std_logic_vector(38, 8),
65064 => conv_std_logic_vector(39, 8),
65065 => conv_std_logic_vector(40, 8),
65066 => conv_std_logic_vector(41, 8),
65067 => conv_std_logic_vector(42, 8),
65068 => conv_std_logic_vector(43, 8),
65069 => conv_std_logic_vector(44, 8),
65070 => conv_std_logic_vector(45, 8),
65071 => conv_std_logic_vector(46, 8),
65072 => conv_std_logic_vector(47, 8),
65073 => conv_std_logic_vector(48, 8),
65074 => conv_std_logic_vector(49, 8),
65075 => conv_std_logic_vector(50, 8),
65076 => conv_std_logic_vector(51, 8),
65077 => conv_std_logic_vector(52, 8),
65078 => conv_std_logic_vector(53, 8),
65079 => conv_std_logic_vector(54, 8),
65080 => conv_std_logic_vector(55, 8),
65081 => conv_std_logic_vector(56, 8),
65082 => conv_std_logic_vector(57, 8),
65083 => conv_std_logic_vector(58, 8),
65084 => conv_std_logic_vector(59, 8),
65085 => conv_std_logic_vector(60, 8),
65086 => conv_std_logic_vector(61, 8),
65087 => conv_std_logic_vector(62, 8),
65088 => conv_std_logic_vector(63, 8),
65089 => conv_std_logic_vector(64, 8),
65090 => conv_std_logic_vector(65, 8),
65091 => conv_std_logic_vector(66, 8),
65092 => conv_std_logic_vector(67, 8),
65093 => conv_std_logic_vector(68, 8),
65094 => conv_std_logic_vector(69, 8),
65095 => conv_std_logic_vector(70, 8),
65096 => conv_std_logic_vector(71, 8),
65097 => conv_std_logic_vector(72, 8),
65098 => conv_std_logic_vector(73, 8),
65099 => conv_std_logic_vector(74, 8),
65100 => conv_std_logic_vector(75, 8),
65101 => conv_std_logic_vector(76, 8),
65102 => conv_std_logic_vector(77, 8),
65103 => conv_std_logic_vector(78, 8),
65104 => conv_std_logic_vector(79, 8),
65105 => conv_std_logic_vector(80, 8),
65106 => conv_std_logic_vector(81, 8),
65107 => conv_std_logic_vector(82, 8),
65108 => conv_std_logic_vector(83, 8),
65109 => conv_std_logic_vector(84, 8),
65110 => conv_std_logic_vector(85, 8),
65111 => conv_std_logic_vector(86, 8),
65112 => conv_std_logic_vector(87, 8),
65113 => conv_std_logic_vector(88, 8),
65114 => conv_std_logic_vector(89, 8),
65115 => conv_std_logic_vector(90, 8),
65116 => conv_std_logic_vector(91, 8),
65117 => conv_std_logic_vector(92, 8),
65118 => conv_std_logic_vector(93, 8),
65119 => conv_std_logic_vector(94, 8),
65120 => conv_std_logic_vector(95, 8),
65121 => conv_std_logic_vector(96, 8),
65122 => conv_std_logic_vector(97, 8),
65123 => conv_std_logic_vector(98, 8),
65124 => conv_std_logic_vector(99, 8),
65125 => conv_std_logic_vector(100, 8),
65126 => conv_std_logic_vector(101, 8),
65127 => conv_std_logic_vector(102, 8),
65128 => conv_std_logic_vector(103, 8),
65129 => conv_std_logic_vector(104, 8),
65130 => conv_std_logic_vector(105, 8),
65131 => conv_std_logic_vector(106, 8),
65132 => conv_std_logic_vector(107, 8),
65133 => conv_std_logic_vector(108, 8),
65134 => conv_std_logic_vector(109, 8),
65135 => conv_std_logic_vector(110, 8),
65136 => conv_std_logic_vector(111, 8),
65137 => conv_std_logic_vector(112, 8),
65138 => conv_std_logic_vector(113, 8),
65139 => conv_std_logic_vector(114, 8),
65140 => conv_std_logic_vector(115, 8),
65141 => conv_std_logic_vector(116, 8),
65142 => conv_std_logic_vector(117, 8),
65143 => conv_std_logic_vector(118, 8),
65144 => conv_std_logic_vector(119, 8),
65145 => conv_std_logic_vector(120, 8),
65146 => conv_std_logic_vector(121, 8),
65147 => conv_std_logic_vector(122, 8),
65148 => conv_std_logic_vector(123, 8),
65149 => conv_std_logic_vector(124, 8),
65150 => conv_std_logic_vector(125, 8),
65151 => conv_std_logic_vector(126, 8),
65152 => conv_std_logic_vector(127, 8),
65153 => conv_std_logic_vector(127, 8),
65154 => conv_std_logic_vector(128, 8),
65155 => conv_std_logic_vector(129, 8),
65156 => conv_std_logic_vector(130, 8),
65157 => conv_std_logic_vector(131, 8),
65158 => conv_std_logic_vector(132, 8),
65159 => conv_std_logic_vector(133, 8),
65160 => conv_std_logic_vector(134, 8),
65161 => conv_std_logic_vector(135, 8),
65162 => conv_std_logic_vector(136, 8),
65163 => conv_std_logic_vector(137, 8),
65164 => conv_std_logic_vector(138, 8),
65165 => conv_std_logic_vector(139, 8),
65166 => conv_std_logic_vector(140, 8),
65167 => conv_std_logic_vector(141, 8),
65168 => conv_std_logic_vector(142, 8),
65169 => conv_std_logic_vector(143, 8),
65170 => conv_std_logic_vector(144, 8),
65171 => conv_std_logic_vector(145, 8),
65172 => conv_std_logic_vector(146, 8),
65173 => conv_std_logic_vector(147, 8),
65174 => conv_std_logic_vector(148, 8),
65175 => conv_std_logic_vector(149, 8),
65176 => conv_std_logic_vector(150, 8),
65177 => conv_std_logic_vector(151, 8),
65178 => conv_std_logic_vector(152, 8),
65179 => conv_std_logic_vector(153, 8),
65180 => conv_std_logic_vector(154, 8),
65181 => conv_std_logic_vector(155, 8),
65182 => conv_std_logic_vector(156, 8),
65183 => conv_std_logic_vector(157, 8),
65184 => conv_std_logic_vector(158, 8),
65185 => conv_std_logic_vector(159, 8),
65186 => conv_std_logic_vector(160, 8),
65187 => conv_std_logic_vector(161, 8),
65188 => conv_std_logic_vector(162, 8),
65189 => conv_std_logic_vector(163, 8),
65190 => conv_std_logic_vector(164, 8),
65191 => conv_std_logic_vector(165, 8),
65192 => conv_std_logic_vector(166, 8),
65193 => conv_std_logic_vector(167, 8),
65194 => conv_std_logic_vector(168, 8),
65195 => conv_std_logic_vector(169, 8),
65196 => conv_std_logic_vector(170, 8),
65197 => conv_std_logic_vector(171, 8),
65198 => conv_std_logic_vector(172, 8),
65199 => conv_std_logic_vector(173, 8),
65200 => conv_std_logic_vector(174, 8),
65201 => conv_std_logic_vector(175, 8),
65202 => conv_std_logic_vector(176, 8),
65203 => conv_std_logic_vector(177, 8),
65204 => conv_std_logic_vector(178, 8),
65205 => conv_std_logic_vector(179, 8),
65206 => conv_std_logic_vector(180, 8),
65207 => conv_std_logic_vector(181, 8),
65208 => conv_std_logic_vector(182, 8),
65209 => conv_std_logic_vector(183, 8),
65210 => conv_std_logic_vector(184, 8),
65211 => conv_std_logic_vector(185, 8),
65212 => conv_std_logic_vector(186, 8),
65213 => conv_std_logic_vector(187, 8),
65214 => conv_std_logic_vector(188, 8),
65215 => conv_std_logic_vector(189, 8),
65216 => conv_std_logic_vector(190, 8),
65217 => conv_std_logic_vector(191, 8),
65218 => conv_std_logic_vector(192, 8),
65219 => conv_std_logic_vector(193, 8),
65220 => conv_std_logic_vector(194, 8),
65221 => conv_std_logic_vector(195, 8),
65222 => conv_std_logic_vector(196, 8),
65223 => conv_std_logic_vector(197, 8),
65224 => conv_std_logic_vector(198, 8),
65225 => conv_std_logic_vector(199, 8),
65226 => conv_std_logic_vector(200, 8),
65227 => conv_std_logic_vector(201, 8),
65228 => conv_std_logic_vector(202, 8),
65229 => conv_std_logic_vector(203, 8),
65230 => conv_std_logic_vector(204, 8),
65231 => conv_std_logic_vector(205, 8),
65232 => conv_std_logic_vector(206, 8),
65233 => conv_std_logic_vector(207, 8),
65234 => conv_std_logic_vector(208, 8),
65235 => conv_std_logic_vector(209, 8),
65236 => conv_std_logic_vector(210, 8),
65237 => conv_std_logic_vector(211, 8),
65238 => conv_std_logic_vector(212, 8),
65239 => conv_std_logic_vector(213, 8),
65240 => conv_std_logic_vector(214, 8),
65241 => conv_std_logic_vector(215, 8),
65242 => conv_std_logic_vector(216, 8),
65243 => conv_std_logic_vector(217, 8),
65244 => conv_std_logic_vector(218, 8),
65245 => conv_std_logic_vector(219, 8),
65246 => conv_std_logic_vector(220, 8),
65247 => conv_std_logic_vector(221, 8),
65248 => conv_std_logic_vector(222, 8),
65249 => conv_std_logic_vector(223, 8),
65250 => conv_std_logic_vector(224, 8),
65251 => conv_std_logic_vector(225, 8),
65252 => conv_std_logic_vector(226, 8),
65253 => conv_std_logic_vector(227, 8),
65254 => conv_std_logic_vector(228, 8),
65255 => conv_std_logic_vector(229, 8),
65256 => conv_std_logic_vector(230, 8),
65257 => conv_std_logic_vector(231, 8),
65258 => conv_std_logic_vector(232, 8),
65259 => conv_std_logic_vector(233, 8),
65260 => conv_std_logic_vector(234, 8),
65261 => conv_std_logic_vector(235, 8),
65262 => conv_std_logic_vector(236, 8),
65263 => conv_std_logic_vector(237, 8),
65264 => conv_std_logic_vector(238, 8),
65265 => conv_std_logic_vector(239, 8),
65266 => conv_std_logic_vector(240, 8),
65267 => conv_std_logic_vector(241, 8),
65268 => conv_std_logic_vector(242, 8),
65269 => conv_std_logic_vector(243, 8),
65270 => conv_std_logic_vector(244, 8),
65271 => conv_std_logic_vector(245, 8),
65272 => conv_std_logic_vector(246, 8),
65273 => conv_std_logic_vector(247, 8),
65274 => conv_std_logic_vector(248, 8),
65275 => conv_std_logic_vector(249, 8),
65276 => conv_std_logic_vector(250, 8),
65277 => conv_std_logic_vector(251, 8),
65278 => conv_std_logic_vector(252, 8),
65279 => conv_std_logic_vector(253, 8),
65280 => conv_std_logic_vector(0, 8),
65281 => conv_std_logic_vector(0, 8),
65282 => conv_std_logic_vector(1, 8),
65283 => conv_std_logic_vector(2, 8),
65284 => conv_std_logic_vector(3, 8),
65285 => conv_std_logic_vector(4, 8),
65286 => conv_std_logic_vector(5, 8),
65287 => conv_std_logic_vector(6, 8),
65288 => conv_std_logic_vector(7, 8),
65289 => conv_std_logic_vector(8, 8),
65290 => conv_std_logic_vector(9, 8),
65291 => conv_std_logic_vector(10, 8),
65292 => conv_std_logic_vector(11, 8),
65293 => conv_std_logic_vector(12, 8),
65294 => conv_std_logic_vector(13, 8),
65295 => conv_std_logic_vector(14, 8),
65296 => conv_std_logic_vector(15, 8),
65297 => conv_std_logic_vector(16, 8),
65298 => conv_std_logic_vector(17, 8),
65299 => conv_std_logic_vector(18, 8),
65300 => conv_std_logic_vector(19, 8),
65301 => conv_std_logic_vector(20, 8),
65302 => conv_std_logic_vector(21, 8),
65303 => conv_std_logic_vector(22, 8),
65304 => conv_std_logic_vector(23, 8),
65305 => conv_std_logic_vector(24, 8),
65306 => conv_std_logic_vector(25, 8),
65307 => conv_std_logic_vector(26, 8),
65308 => conv_std_logic_vector(27, 8),
65309 => conv_std_logic_vector(28, 8),
65310 => conv_std_logic_vector(29, 8),
65311 => conv_std_logic_vector(30, 8),
65312 => conv_std_logic_vector(31, 8),
65313 => conv_std_logic_vector(32, 8),
65314 => conv_std_logic_vector(33, 8),
65315 => conv_std_logic_vector(34, 8),
65316 => conv_std_logic_vector(35, 8),
65317 => conv_std_logic_vector(36, 8),
65318 => conv_std_logic_vector(37, 8),
65319 => conv_std_logic_vector(38, 8),
65320 => conv_std_logic_vector(39, 8),
65321 => conv_std_logic_vector(40, 8),
65322 => conv_std_logic_vector(41, 8),
65323 => conv_std_logic_vector(42, 8),
65324 => conv_std_logic_vector(43, 8),
65325 => conv_std_logic_vector(44, 8),
65326 => conv_std_logic_vector(45, 8),
65327 => conv_std_logic_vector(46, 8),
65328 => conv_std_logic_vector(47, 8),
65329 => conv_std_logic_vector(48, 8),
65330 => conv_std_logic_vector(49, 8),
65331 => conv_std_logic_vector(50, 8),
65332 => conv_std_logic_vector(51, 8),
65333 => conv_std_logic_vector(52, 8),
65334 => conv_std_logic_vector(53, 8),
65335 => conv_std_logic_vector(54, 8),
65336 => conv_std_logic_vector(55, 8),
65337 => conv_std_logic_vector(56, 8),
65338 => conv_std_logic_vector(57, 8),
65339 => conv_std_logic_vector(58, 8),
65340 => conv_std_logic_vector(59, 8),
65341 => conv_std_logic_vector(60, 8),
65342 => conv_std_logic_vector(61, 8),
65343 => conv_std_logic_vector(62, 8),
65344 => conv_std_logic_vector(63, 8),
65345 => conv_std_logic_vector(64, 8),
65346 => conv_std_logic_vector(65, 8),
65347 => conv_std_logic_vector(66, 8),
65348 => conv_std_logic_vector(67, 8),
65349 => conv_std_logic_vector(68, 8),
65350 => conv_std_logic_vector(69, 8),
65351 => conv_std_logic_vector(70, 8),
65352 => conv_std_logic_vector(71, 8),
65353 => conv_std_logic_vector(72, 8),
65354 => conv_std_logic_vector(73, 8),
65355 => conv_std_logic_vector(74, 8),
65356 => conv_std_logic_vector(75, 8),
65357 => conv_std_logic_vector(76, 8),
65358 => conv_std_logic_vector(77, 8),
65359 => conv_std_logic_vector(78, 8),
65360 => conv_std_logic_vector(79, 8),
65361 => conv_std_logic_vector(80, 8),
65362 => conv_std_logic_vector(81, 8),
65363 => conv_std_logic_vector(82, 8),
65364 => conv_std_logic_vector(83, 8),
65365 => conv_std_logic_vector(84, 8),
65366 => conv_std_logic_vector(85, 8),
65367 => conv_std_logic_vector(86, 8),
65368 => conv_std_logic_vector(87, 8),
65369 => conv_std_logic_vector(88, 8),
65370 => conv_std_logic_vector(89, 8),
65371 => conv_std_logic_vector(90, 8),
65372 => conv_std_logic_vector(91, 8),
65373 => conv_std_logic_vector(92, 8),
65374 => conv_std_logic_vector(93, 8),
65375 => conv_std_logic_vector(94, 8),
65376 => conv_std_logic_vector(95, 8),
65377 => conv_std_logic_vector(96, 8),
65378 => conv_std_logic_vector(97, 8),
65379 => conv_std_logic_vector(98, 8),
65380 => conv_std_logic_vector(99, 8),
65381 => conv_std_logic_vector(100, 8),
65382 => conv_std_logic_vector(101, 8),
65383 => conv_std_logic_vector(102, 8),
65384 => conv_std_logic_vector(103, 8),
65385 => conv_std_logic_vector(104, 8),
65386 => conv_std_logic_vector(105, 8),
65387 => conv_std_logic_vector(106, 8),
65388 => conv_std_logic_vector(107, 8),
65389 => conv_std_logic_vector(108, 8),
65390 => conv_std_logic_vector(109, 8),
65391 => conv_std_logic_vector(110, 8),
65392 => conv_std_logic_vector(111, 8),
65393 => conv_std_logic_vector(112, 8),
65394 => conv_std_logic_vector(113, 8),
65395 => conv_std_logic_vector(114, 8),
65396 => conv_std_logic_vector(115, 8),
65397 => conv_std_logic_vector(116, 8),
65398 => conv_std_logic_vector(117, 8),
65399 => conv_std_logic_vector(118, 8),
65400 => conv_std_logic_vector(119, 8),
65401 => conv_std_logic_vector(120, 8),
65402 => conv_std_logic_vector(121, 8),
65403 => conv_std_logic_vector(122, 8),
65404 => conv_std_logic_vector(123, 8),
65405 => conv_std_logic_vector(124, 8),
65406 => conv_std_logic_vector(125, 8),
65407 => conv_std_logic_vector(126, 8),
65408 => conv_std_logic_vector(127, 8),
65409 => conv_std_logic_vector(128, 8),
65410 => conv_std_logic_vector(129, 8),
65411 => conv_std_logic_vector(130, 8),
65412 => conv_std_logic_vector(131, 8),
65413 => conv_std_logic_vector(132, 8),
65414 => conv_std_logic_vector(133, 8),
65415 => conv_std_logic_vector(134, 8),
65416 => conv_std_logic_vector(135, 8),
65417 => conv_std_logic_vector(136, 8),
65418 => conv_std_logic_vector(137, 8),
65419 => conv_std_logic_vector(138, 8),
65420 => conv_std_logic_vector(139, 8),
65421 => conv_std_logic_vector(140, 8),
65422 => conv_std_logic_vector(141, 8),
65423 => conv_std_logic_vector(142, 8),
65424 => conv_std_logic_vector(143, 8),
65425 => conv_std_logic_vector(144, 8),
65426 => conv_std_logic_vector(145, 8),
65427 => conv_std_logic_vector(146, 8),
65428 => conv_std_logic_vector(147, 8),
65429 => conv_std_logic_vector(148, 8),
65430 => conv_std_logic_vector(149, 8),
65431 => conv_std_logic_vector(150, 8),
65432 => conv_std_logic_vector(151, 8),
65433 => conv_std_logic_vector(152, 8),
65434 => conv_std_logic_vector(153, 8),
65435 => conv_std_logic_vector(154, 8),
65436 => conv_std_logic_vector(155, 8),
65437 => conv_std_logic_vector(156, 8),
65438 => conv_std_logic_vector(157, 8),
65439 => conv_std_logic_vector(158, 8),
65440 => conv_std_logic_vector(159, 8),
65441 => conv_std_logic_vector(160, 8),
65442 => conv_std_logic_vector(161, 8),
65443 => conv_std_logic_vector(162, 8),
65444 => conv_std_logic_vector(163, 8),
65445 => conv_std_logic_vector(164, 8),
65446 => conv_std_logic_vector(165, 8),
65447 => conv_std_logic_vector(166, 8),
65448 => conv_std_logic_vector(167, 8),
65449 => conv_std_logic_vector(168, 8),
65450 => conv_std_logic_vector(169, 8),
65451 => conv_std_logic_vector(170, 8),
65452 => conv_std_logic_vector(171, 8),
65453 => conv_std_logic_vector(172, 8),
65454 => conv_std_logic_vector(173, 8),
65455 => conv_std_logic_vector(174, 8),
65456 => conv_std_logic_vector(175, 8),
65457 => conv_std_logic_vector(176, 8),
65458 => conv_std_logic_vector(177, 8),
65459 => conv_std_logic_vector(178, 8),
65460 => conv_std_logic_vector(179, 8),
65461 => conv_std_logic_vector(180, 8),
65462 => conv_std_logic_vector(181, 8),
65463 => conv_std_logic_vector(182, 8),
65464 => conv_std_logic_vector(183, 8),
65465 => conv_std_logic_vector(184, 8),
65466 => conv_std_logic_vector(185, 8),
65467 => conv_std_logic_vector(186, 8),
65468 => conv_std_logic_vector(187, 8),
65469 => conv_std_logic_vector(188, 8),
65470 => conv_std_logic_vector(189, 8),
65471 => conv_std_logic_vector(190, 8),
65472 => conv_std_logic_vector(191, 8),
65473 => conv_std_logic_vector(192, 8),
65474 => conv_std_logic_vector(193, 8),
65475 => conv_std_logic_vector(194, 8),
65476 => conv_std_logic_vector(195, 8),
65477 => conv_std_logic_vector(196, 8),
65478 => conv_std_logic_vector(197, 8),
65479 => conv_std_logic_vector(198, 8),
65480 => conv_std_logic_vector(199, 8),
65481 => conv_std_logic_vector(200, 8),
65482 => conv_std_logic_vector(201, 8),
65483 => conv_std_logic_vector(202, 8),
65484 => conv_std_logic_vector(203, 8),
65485 => conv_std_logic_vector(204, 8),
65486 => conv_std_logic_vector(205, 8),
65487 => conv_std_logic_vector(206, 8),
65488 => conv_std_logic_vector(207, 8),
65489 => conv_std_logic_vector(208, 8),
65490 => conv_std_logic_vector(209, 8),
65491 => conv_std_logic_vector(210, 8),
65492 => conv_std_logic_vector(211, 8),
65493 => conv_std_logic_vector(212, 8),
65494 => conv_std_logic_vector(213, 8),
65495 => conv_std_logic_vector(214, 8),
65496 => conv_std_logic_vector(215, 8),
65497 => conv_std_logic_vector(216, 8),
65498 => conv_std_logic_vector(217, 8),
65499 => conv_std_logic_vector(218, 8),
65500 => conv_std_logic_vector(219, 8),
65501 => conv_std_logic_vector(220, 8),
65502 => conv_std_logic_vector(221, 8),
65503 => conv_std_logic_vector(222, 8),
65504 => conv_std_logic_vector(223, 8),
65505 => conv_std_logic_vector(224, 8),
65506 => conv_std_logic_vector(225, 8),
65507 => conv_std_logic_vector(226, 8),
65508 => conv_std_logic_vector(227, 8),
65509 => conv_std_logic_vector(228, 8),
65510 => conv_std_logic_vector(229, 8),
65511 => conv_std_logic_vector(230, 8),
65512 => conv_std_logic_vector(231, 8),
65513 => conv_std_logic_vector(232, 8),
65514 => conv_std_logic_vector(233, 8),
65515 => conv_std_logic_vector(234, 8),
65516 => conv_std_logic_vector(235, 8),
65517 => conv_std_logic_vector(236, 8),
65518 => conv_std_logic_vector(237, 8),
65519 => conv_std_logic_vector(238, 8),
65520 => conv_std_logic_vector(239, 8),
65521 => conv_std_logic_vector(240, 8),
65522 => conv_std_logic_vector(241, 8),
65523 => conv_std_logic_vector(242, 8),
65524 => conv_std_logic_vector(243, 8),
65525 => conv_std_logic_vector(244, 8),
65526 => conv_std_logic_vector(245, 8),
65527 => conv_std_logic_vector(246, 8),
65528 => conv_std_logic_vector(247, 8),
65529 => conv_std_logic_vector(248, 8),
65530 => conv_std_logic_vector(249, 8),
65531 => conv_std_logic_vector(250, 8),
65532 => conv_std_logic_vector(251, 8),
65533 => conv_std_logic_vector(252, 8),
65534 => conv_std_logic_vector(253, 8),
65535 => conv_std_logic_vector(254, 8),
OTHERS => conv_std_logic_vector( 0, 8)
  );       

begin
    process(clk)
    begin
       if( clk'event and clk = '1' ) then
          ROM_data <= Content(conv_integer(ROM_addr));
       end if;
    end process;
end a;
