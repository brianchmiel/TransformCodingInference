library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_SIGNED.ALL;

entity ConvLayer1_256 is
  generic (
  	       mult_sum      : string := "sum";
           N             : integer := 8; -- input data width
           M             : integer := 8; -- input weight width
           W             : integer := 8; -- output data width      (Note, W+SR <= N+M+4)
           SR            : integer := 2 -- data shift right before output
  	       );
  port    (
           clk     : in std_logic;
           rst     : in std_logic;
  	       d01_in, d65_in , d129_in, d193_in   : in std_logic_vector (9*N-1 downto 0);
           d02_in, d66_in , d130_in, d194_in   : in std_logic_vector (9*N-1 downto 0);
           d03_in, d67_in , d131_in, d195_in   : in std_logic_vector (9*N-1 downto 0);
           d04_in, d68_in , d132_in, d196_in   : in std_logic_vector (9*N-1 downto 0);
           d05_in, d69_in , d133_in, d197_in   : in std_logic_vector (9*N-1 downto 0);
           d06_in, d70_in , d134_in, d198_in   : in std_logic_vector (9*N-1 downto 0);
           d07_in, d71_in , d135_in, d199_in   : in std_logic_vector (9*N-1 downto 0);
           d08_in, d72_in , d136_in, d200_in   : in std_logic_vector (9*N-1 downto 0);
           d09_in, d73_in , d137_in, d201_in   : in std_logic_vector (9*N-1 downto 0);
           d10_in, d74_in , d138_in, d202_in   : in std_logic_vector (9*N-1 downto 0);
           d11_in, d75_in , d139_in, d203_in   : in std_logic_vector (9*N-1 downto 0);
           d12_in, d76_in , d140_in, d204_in   : in std_logic_vector (9*N-1 downto 0);
           d13_in, d77_in , d141_in, d205_in   : in std_logic_vector (9*N-1 downto 0);
           d14_in, d78_in , d142_in, d206_in   : in std_logic_vector (9*N-1 downto 0);
           d15_in, d79_in , d143_in, d207_in   : in std_logic_vector (9*N-1 downto 0);
           d16_in, d80_in , d144_in, d208_in   : in std_logic_vector (9*N-1 downto 0);
           d17_in, d81_in , d145_in, d209_in   : in std_logic_vector (9*N-1 downto 0);
           d18_in, d82_in , d146_in, d210_in   : in std_logic_vector (9*N-1 downto 0);
           d19_in, d83_in , d147_in, d211_in   : in std_logic_vector (9*N-1 downto 0);
           d20_in, d84_in , d148_in, d212_in   : in std_logic_vector (9*N-1 downto 0);
           d21_in, d85_in , d149_in, d213_in   : in std_logic_vector (9*N-1 downto 0);
           d22_in, d86_in , d150_in, d214_in   : in std_logic_vector (9*N-1 downto 0);
           d23_in, d87_in , d151_in, d215_in   : in std_logic_vector (9*N-1 downto 0);
           d24_in, d88_in , d152_in, d216_in   : in std_logic_vector (9*N-1 downto 0);
           d25_in, d89_in , d153_in, d217_in   : in std_logic_vector (9*N-1 downto 0);
           d26_in, d90_in , d154_in, d218_in   : in std_logic_vector (9*N-1 downto 0);
           d27_in, d91_in , d155_in, d219_in   : in std_logic_vector (9*N-1 downto 0);
           d28_in, d92_in , d156_in, d220_in   : in std_logic_vector (9*N-1 downto 0);
           d29_in, d93_in , d157_in, d221_in   : in std_logic_vector (9*N-1 downto 0);
           d30_in, d94_in , d158_in, d222_in   : in std_logic_vector (9*N-1 downto 0);
           d31_in, d95_in , d159_in, d223_in   : in std_logic_vector (9*N-1 downto 0);
           d32_in, d96_in , d160_in, d224_in   : in std_logic_vector (9*N-1 downto 0);
           d33_in, d97_in , d161_in, d225_in   : in std_logic_vector (9*N-1 downto 0);
           d34_in, d98_in , d162_in, d226_in   : in std_logic_vector (9*N-1 downto 0);
           d35_in, d99_in , d163_in, d227_in   : in std_logic_vector (9*N-1 downto 0);
           d36_in, d100_in, d164_in, d228_in   : in std_logic_vector (9*N-1 downto 0);
           d37_in, d101_in, d165_in, d229_in   : in std_logic_vector (9*N-1 downto 0);
           d38_in, d102_in, d166_in, d230_in   : in std_logic_vector (9*N-1 downto 0);
           d39_in, d103_in, d167_in, d231_in   : in std_logic_vector (9*N-1 downto 0);
           d40_in, d104_in, d168_in, d232_in   : in std_logic_vector (9*N-1 downto 0);
           d41_in, d105_in, d169_in, d233_in   : in std_logic_vector (9*N-1 downto 0);
           d42_in, d106_in, d170_in, d234_in   : in std_logic_vector (9*N-1 downto 0);
           d43_in, d107_in, d171_in, d235_in   : in std_logic_vector (9*N-1 downto 0);
           d44_in, d108_in, d172_in, d236_in   : in std_logic_vector (9*N-1 downto 0);
           d45_in, d109_in, d173_in, d237_in   : in std_logic_vector (9*N-1 downto 0);
           d46_in, d110_in, d174_in, d238_in   : in std_logic_vector (9*N-1 downto 0);
           d47_in, d111_in, d175_in, d239_in   : in std_logic_vector (9*N-1 downto 0);
           d48_in, d112_in, d176_in, d240_in   : in std_logic_vector (9*N-1 downto 0);
           d49_in, d113_in, d177_in, d241_in   : in std_logic_vector (9*N-1 downto 0);
           d50_in, d114_in, d178_in, d242_in   : in std_logic_vector (9*N-1 downto 0);
           d51_in, d115_in, d179_in, d243_in   : in std_logic_vector (9*N-1 downto 0);
           d52_in, d116_in, d180_in, d244_in   : in std_logic_vector (9*N-1 downto 0);
           d53_in, d117_in, d181_in, d245_in   : in std_logic_vector (9*N-1 downto 0);
           d54_in, d118_in, d182_in, d246_in   : in std_logic_vector (9*N-1 downto 0);
           d55_in, d119_in, d183_in, d247_in   : in std_logic_vector (9*N-1 downto 0);
           d56_in, d120_in, d184_in, d248_in   : in std_logic_vector (9*N-1 downto 0);
           d57_in, d121_in, d185_in, d249_in   : in std_logic_vector (9*N-1 downto 0);
           d58_in, d122_in, d186_in, d250_in   : in std_logic_vector (9*N-1 downto 0);
           d59_in, d123_in, d187_in, d251_in   : in std_logic_vector (9*N-1 downto 0);
           d60_in, d124_in, d188_in, d252_in   : in std_logic_vector (9*N-1 downto 0);
           d61_in, d125_in, d189_in, d253_in   : in std_logic_vector (9*N-1 downto 0);
           d62_in, d126_in, d190_in, d254_in   : in std_logic_vector (9*N-1 downto 0);
           d63_in, d127_in, d191_in, d255_in   : in std_logic_vector (9*N-1 downto 0);
           d64_in, d128_in, d192_in, d256_in   : in std_logic_vector (9*N-1 downto 0);
  	       en_in     : in std_logic;
  	       sof_in    : in std_logic; -- start of frame
  	       --sol     : in std_logic; -- start of line
  	       --eof     : in std_logic; -- end of frame

           w01_in, w65_in , w129_in, w193_in   : in std_logic_vector(9*M-1 downto 0);
           w02_in, w66_in , w130_in, w194_in   : in std_logic_vector(9*M-1 downto 0);
           w03_in, w67_in , w131_in, w195_in   : in std_logic_vector(9*M-1 downto 0);
           w04_in, w68_in , w132_in, w196_in   : in std_logic_vector(9*M-1 downto 0);
           w05_in, w69_in , w133_in, w197_in   : in std_logic_vector(9*M-1 downto 0);
           w06_in, w70_in , w134_in, w198_in   : in std_logic_vector(9*M-1 downto 0);
           w07_in, w71_in , w135_in, w199_in   : in std_logic_vector(9*M-1 downto 0);
           w08_in, w72_in , w136_in, w200_in   : in std_logic_vector(9*M-1 downto 0);
           w09_in, w73_in , w137_in, w201_in   : in std_logic_vector(9*M-1 downto 0);
           w10_in, w74_in , w138_in, w202_in   : in std_logic_vector(9*M-1 downto 0);
           w11_in, w75_in , w139_in, w203_in   : in std_logic_vector(9*M-1 downto 0);
           w12_in, w76_in , w140_in, w204_in   : in std_logic_vector(9*M-1 downto 0);
           w13_in, w77_in , w141_in, w205_in   : in std_logic_vector(9*M-1 downto 0);
           w14_in, w78_in , w142_in, w206_in   : in std_logic_vector(9*M-1 downto 0);
           w15_in, w79_in , w143_in, w207_in   : in std_logic_vector(9*M-1 downto 0);
           w16_in, w80_in , w144_in, w208_in   : in std_logic_vector(9*M-1 downto 0);
           w17_in, w81_in , w145_in, w209_in   : in std_logic_vector(9*M-1 downto 0);
           w18_in, w82_in , w146_in, w210_in   : in std_logic_vector(9*M-1 downto 0);
           w19_in, w83_in , w147_in, w211_in   : in std_logic_vector(9*M-1 downto 0);
           w20_in, w84_in , w148_in, w212_in   : in std_logic_vector(9*M-1 downto 0);
           w21_in, w85_in , w149_in, w213_in   : in std_logic_vector(9*M-1 downto 0);
           w22_in, w86_in , w150_in, w214_in   : in std_logic_vector(9*M-1 downto 0);
           w23_in, w87_in , w151_in, w215_in   : in std_logic_vector(9*M-1 downto 0);
           w24_in, w88_in , w152_in, w216_in   : in std_logic_vector(9*M-1 downto 0);
           w25_in, w89_in , w153_in, w217_in   : in std_logic_vector(9*M-1 downto 0);
           w26_in, w90_in , w154_in, w218_in   : in std_logic_vector(9*M-1 downto 0);
           w27_in, w91_in , w155_in, w219_in   : in std_logic_vector(9*M-1 downto 0);
           w28_in, w92_in , w156_in, w220_in   : in std_logic_vector(9*M-1 downto 0);
           w29_in, w93_in , w157_in, w221_in   : in std_logic_vector(9*M-1 downto 0);
           w30_in, w94_in , w158_in, w222_in   : in std_logic_vector(9*M-1 downto 0);
           w31_in, w95_in , w159_in, w223_in   : in std_logic_vector(9*M-1 downto 0);
           w32_in, w96_in , w160_in, w224_in   : in std_logic_vector(9*M-1 downto 0);
           w33_in, w97_in , w161_in, w225_in   : in std_logic_vector(9*M-1 downto 0);
           w34_in, w98_in , w162_in, w226_in   : in std_logic_vector(9*M-1 downto 0);
           w35_in, w99_in , w163_in, w227_in   : in std_logic_vector(9*M-1 downto 0);
           w36_in, w100_in, w164_in, w228_in   : in std_logic_vector(9*M-1 downto 0);
           w37_in, w101_in, w165_in, w229_in   : in std_logic_vector(9*M-1 downto 0);
           w38_in, w102_in, w166_in, w230_in   : in std_logic_vector(9*M-1 downto 0);
           w39_in, w103_in, w167_in, w231_in   : in std_logic_vector(9*M-1 downto 0);
           w40_in, w104_in, w168_in, w232_in   : in std_logic_vector(9*M-1 downto 0);
           w41_in, w105_in, w169_in, w233_in   : in std_logic_vector(9*M-1 downto 0);
           w42_in, w106_in, w170_in, w234_in   : in std_logic_vector(9*M-1 downto 0);
           w43_in, w107_in, w171_in, w235_in   : in std_logic_vector(9*M-1 downto 0);
           w44_in, w108_in, w172_in, w236_in   : in std_logic_vector(9*M-1 downto 0);
           w45_in, w109_in, w173_in, w237_in   : in std_logic_vector(9*M-1 downto 0);
           w46_in, w110_in, w174_in, w238_in   : in std_logic_vector(9*M-1 downto 0);
           w47_in, w111_in, w175_in, w239_in   : in std_logic_vector(9*M-1 downto 0);
           w48_in, w112_in, w176_in, w240_in   : in std_logic_vector(9*M-1 downto 0);
           w49_in, w113_in, w177_in, w241_in   : in std_logic_vector(9*M-1 downto 0);
           w50_in, w114_in, w178_in, w242_in   : in std_logic_vector(9*M-1 downto 0);
           w51_in, w115_in, w179_in, w243_in   : in std_logic_vector(9*M-1 downto 0);
           w52_in, w116_in, w180_in, w244_in   : in std_logic_vector(9*M-1 downto 0);
           w53_in, w117_in, w181_in, w245_in   : in std_logic_vector(9*M-1 downto 0);
           w54_in, w118_in, w182_in, w246_in   : in std_logic_vector(9*M-1 downto 0);
           w55_in, w119_in, w183_in, w247_in   : in std_logic_vector(9*M-1 downto 0);
           w56_in, w120_in, w184_in, w248_in   : in std_logic_vector(9*M-1 downto 0);
           w57_in, w121_in, w185_in, w249_in   : in std_logic_vector(9*M-1 downto 0);
           w58_in, w122_in, w186_in, w250_in   : in std_logic_vector(9*M-1 downto 0);
           w59_in, w123_in, w187_in, w251_in   : in std_logic_vector(9*M-1 downto 0);
           w60_in, w124_in, w188_in, w252_in   : in std_logic_vector(9*M-1 downto 0);
           w61_in, w125_in, w189_in, w253_in   : in std_logic_vector(9*M-1 downto 0);
           w62_in, w126_in, w190_in, w254_in   : in std_logic_vector(9*M-1 downto 0);
           w63_in, w127_in, w191_in, w255_in   : in std_logic_vector(9*M-1 downto 0);
           w64_in, w128_in, w192_in, w256_in   : in std_logic_vector(9*M-1 downto 0);

           d_out   : out std_logic_vector (W-1 downto 0);
           en_out    : out std_logic;
           sof_out   : out std_logic);
end ConvLayer1_256;

architecture a of ConvLayer1_256 is

constant EN_BIT  : integer range 0 to 1 := 0;
constant SOF_BIT : integer range 0 to 1 := 1;

component Binary_adder8 is
  generic (
           N             : integer := 8;                  -- input #1 data width, positive
           M             : integer := 8
           );
  port    (
           clk           : in  std_logic;
           rst           : in  std_logic; 

           en_in         : in  std_logic;                         
           Multiplier    : in  std_logic_vector(N-1 downto 0);    -- positive
           Multiplicand  : in  std_logic_vector(8-1 downto 0);    -- signed

           d_out         : out std_logic_vector (N + M - 1 downto 0);
           en_out        : out std_logic);                        
end component;

component ConvLayer1 is
  generic (
           mult_sum      : string := "sum";
           N             : integer := 8; -- input data width
           M             : integer := 8; -- input weight width
           W             : integer := 8; -- output data width      (Note, W+SR <= N+M+4)
           SR            : integer := 2 -- data shift right before output
           );
  port    (
           clk         : in std_logic;
           rst         : in std_logic;
           data2conv1  : in std_logic_vector (N-1 downto 0);
           data2conv2  : in std_logic_vector (N-1 downto 0);
           data2conv3  : in std_logic_vector (N-1 downto 0);
           data2conv4  : in std_logic_vector (N-1 downto 0);
           data2conv5  : in std_logic_vector (N-1 downto 0);
           data2conv6  : in std_logic_vector (N-1 downto 0);
           data2conv7  : in std_logic_vector (N-1 downto 0);
           data2conv8  : in std_logic_vector (N-1 downto 0);
           data2conv9  : in std_logic_vector (N-1 downto 0);
           en_in       : in std_logic;
           sof_in      : in std_logic; -- start of frame
           --sol     : in std_logic; -- start of line
           --eof     : in std_logic; -- end of frame

          w1           : in std_logic_vector(M-1 downto 0); -- weight matrix
          w2           : in std_logic_vector(M-1 downto 0); -- weight matrix
          w3           : in std_logic_vector(M-1 downto 0); -- weight matrix
          w4           : in std_logic_vector(M-1 downto 0); -- weight matrix
          w5           : in std_logic_vector(M-1 downto 0); -- weight matrix
          w6           : in std_logic_vector(M-1 downto 0); -- weight matrix
          w7           : in std_logic_vector(M-1 downto 0); -- weight matrix
          w8           : in std_logic_vector(M-1 downto 0); -- weight matrix
          w9           : in std_logic_vector(M-1 downto 0); -- weight matrix

           d_out       : out std_logic_vector (W-1 downto 0);
           en_out      : out std_logic;
           sof_out     : out std_logic);
end component;

signal    d01_out, d65_out , d129_out, d193_out   : std_logic_vector (W-1 downto 0);
signal    d02_out, d66_out , d130_out, d194_out   : std_logic_vector (W-1 downto 0);
signal    d03_out, d67_out , d131_out, d195_out   : std_logic_vector (W-1 downto 0);
signal    d04_out, d68_out , d132_out, d196_out   : std_logic_vector (W-1 downto 0);
signal    d05_out, d69_out , d133_out, d197_out   : std_logic_vector (W-1 downto 0);
signal    d06_out, d70_out , d134_out, d198_out   : std_logic_vector (W-1 downto 0);
signal    d07_out, d71_out , d135_out, d199_out   : std_logic_vector (W-1 downto 0);
signal    d08_out, d72_out , d136_out, d200_out   : std_logic_vector (W-1 downto 0);
signal    d09_out, d73_out , d137_out, d201_out   : std_logic_vector (W-1 downto 0);
signal    d10_out, d74_out , d138_out, d202_out   : std_logic_vector (W-1 downto 0);
signal    d11_out, d75_out , d139_out, d203_out   : std_logic_vector (W-1 downto 0);
signal    d12_out, d76_out , d140_out, d204_out   : std_logic_vector (W-1 downto 0);
signal    d13_out, d77_out , d141_out, d205_out   : std_logic_vector (W-1 downto 0);
signal    d14_out, d78_out , d142_out, d206_out   : std_logic_vector (W-1 downto 0);
signal    d15_out, d79_out , d143_out, d207_out   : std_logic_vector (W-1 downto 0);
signal    d16_out, d80_out , d144_out, d208_out   : std_logic_vector (W-1 downto 0);
signal    d17_out, d81_out , d145_out, d209_out   : std_logic_vector (W-1 downto 0);
signal    d18_out, d82_out , d146_out, d210_out   : std_logic_vector (W-1 downto 0);
signal    d19_out, d83_out , d147_out, d211_out   : std_logic_vector (W-1 downto 0);
signal    d20_out, d84_out , d148_out, d212_out   : std_logic_vector (W-1 downto 0);
signal    d21_out, d85_out , d149_out, d213_out   : std_logic_vector (W-1 downto 0);
signal    d22_out, d86_out , d150_out, d214_out   : std_logic_vector (W-1 downto 0);
signal    d23_out, d87_out , d151_out, d215_out   : std_logic_vector (W-1 downto 0);
signal    d24_out, d88_out , d152_out, d216_out   : std_logic_vector (W-1 downto 0);
signal    d25_out, d89_out , d153_out, d217_out   : std_logic_vector (W-1 downto 0);
signal    d26_out, d90_out , d154_out, d218_out   : std_logic_vector (W-1 downto 0);
signal    d27_out, d91_out , d155_out, d219_out   : std_logic_vector (W-1 downto 0);
signal    d28_out, d92_out , d156_out, d220_out   : std_logic_vector (W-1 downto 0);
signal    d29_out, d93_out , d157_out, d221_out   : std_logic_vector (W-1 downto 0);
signal    d30_out, d94_out , d158_out, d222_out   : std_logic_vector (W-1 downto 0);
signal    d31_out, d95_out , d159_out, d223_out   : std_logic_vector (W-1 downto 0);
signal    d32_out, d96_out , d160_out, d224_out   : std_logic_vector (W-1 downto 0);
signal    d33_out, d97_out , d161_out, d225_out   : std_logic_vector (W-1 downto 0);
signal    d34_out, d98_out , d162_out, d226_out   : std_logic_vector (W-1 downto 0);
signal    d35_out, d99_out , d163_out, d227_out   : std_logic_vector (W-1 downto 0);
signal    d36_out, d100_out, d164_out, d228_out   : std_logic_vector (W-1 downto 0);
signal    d37_out, d101_out, d165_out, d229_out   : std_logic_vector (W-1 downto 0);
signal    d38_out, d102_out, d166_out, d230_out   : std_logic_vector (W-1 downto 0);
signal    d39_out, d103_out, d167_out, d231_out   : std_logic_vector (W-1 downto 0);
signal    d40_out, d104_out, d168_out, d232_out   : std_logic_vector (W-1 downto 0);
signal    d41_out, d105_out, d169_out, d233_out   : std_logic_vector (W-1 downto 0);
signal    d42_out, d106_out, d170_out, d234_out   : std_logic_vector (W-1 downto 0);
signal    d43_out, d107_out, d171_out, d235_out   : std_logic_vector (W-1 downto 0);
signal    d44_out, d108_out, d172_out, d236_out   : std_logic_vector (W-1 downto 0);
signal    d45_out, d109_out, d173_out, d237_out   : std_logic_vector (W-1 downto 0);
signal    d46_out, d110_out, d174_out, d238_out   : std_logic_vector (W-1 downto 0);
signal    d47_out, d111_out, d175_out, d239_out   : std_logic_vector (W-1 downto 0);
signal    d48_out, d112_out, d176_out, d240_out   : std_logic_vector (W-1 downto 0);
signal    d49_out, d113_out, d177_out, d241_out   : std_logic_vector (W-1 downto 0);
signal    d50_out, d114_out, d178_out, d242_out   : std_logic_vector (W-1 downto 0);
signal    d51_out, d115_out, d179_out, d243_out   : std_logic_vector (W-1 downto 0);
signal    d52_out, d116_out, d180_out, d244_out   : std_logic_vector (W-1 downto 0);
signal    d53_out, d117_out, d181_out, d245_out   : std_logic_vector (W-1 downto 0);
signal    d54_out, d118_out, d182_out, d246_out   : std_logic_vector (W-1 downto 0);
signal    d55_out, d119_out, d183_out, d247_out   : std_logic_vector (W-1 downto 0);
signal    d56_out, d120_out, d184_out, d248_out   : std_logic_vector (W-1 downto 0);
signal    d57_out, d121_out, d185_out, d249_out   : std_logic_vector (W-1 downto 0);
signal    d58_out, d122_out, d186_out, d250_out   : std_logic_vector (W-1 downto 0);
signal    d59_out, d123_out, d187_out, d251_out   : std_logic_vector (W-1 downto 0);
signal    d60_out, d124_out, d188_out, d252_out   : std_logic_vector (W-1 downto 0);
signal    d61_out, d125_out, d189_out, d253_out   : std_logic_vector (W-1 downto 0);
signal    d62_out, d126_out, d190_out, d254_out   : std_logic_vector (W-1 downto 0);
signal    d63_out, d127_out, d191_out, d255_out   : std_logic_vector (W-1 downto 0);
signal    d64_out, d128_out, d192_out, d256_out   : std_logic_vector (W-1 downto 0);

signal    sum1 , sum22, sum44, sum60     : std_logic_vector (W+1 downto 0); 
signal    sum2 , sum23, sum45, sum61     : std_logic_vector (W+1 downto 0); 
signal    sum3 , sum24, sum46, sum62     : std_logic_vector (W+1 downto 0); 
signal    sum4 , sum25, sum47, sum63     : std_logic_vector (W+1 downto 0); 
signal    sum5 , sum26, sum48, sum64     : std_logic_vector (W+1 downto 0); 
signal    sum6 , sum27, sum49, sum65     : std_logic_vector (W+1 downto 0); 
signal    sum7 , sum28, sum50, sum66     : std_logic_vector (W+1 downto 0); 
signal    sum8 , sum29, sum51, sum67     : std_logic_vector (W+1 downto 0); 
signal    sum9 , sum30, sum52, sum68     : std_logic_vector (W+1 downto 0); 
signal    sum10, sum31, sum53, sum69     : std_logic_vector (W+1 downto 0); 
signal    sum11, sum32, sum54, sum70     : std_logic_vector (W+1 downto 0); 
signal    sum12, sum33, sum55, sum71     : std_logic_vector (W+1 downto 0); 
signal    sum13, sum34, sum56, sum72     : std_logic_vector (W+1 downto 0); 
signal    sum14, sum35, sum57, sum73     : std_logic_vector (W+1 downto 0); 
signal    sum15, sum36, sum58, sum74     : std_logic_vector (W+1 downto 0); 
signal    sum16, sum37, sum59, sum75     : std_logic_vector (W+1 downto 0); 
       
signal    sum17, sum38, sum76, sum80     : std_logic_vector (W+3 downto 0);   
signal    sum18, sum39, sum77, sum81     : std_logic_vector (W+3 downto 0);   
signal    sum19, sum40, sum78, sum82     : std_logic_vector (W+3 downto 0); 
signal    sum20, sum41, sum79, sum83     : std_logic_vector (W+3 downto 0); 
       
signal    sum21, sum42, sum84, sum85     : std_logic_vector (W+5 downto 0); 

signal    sum43            : std_logic_vector (W+7 downto 0); 

begin


CL01: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d01_in(9*N-1 downto 8*N),data2conv2 =>d01_in(8*N-1 downto 7*N),data2conv3 =>d01_in(7*N-1 downto 6*N),data2conv4 =>d01_in(6*N-1 downto 5*N),data2conv5 =>d01_in(5*N-1 downto 4*N),data2conv6 =>d01_in(4*N-1 downto 3*N),data2conv7 =>d01_in(3*N-1 downto 2*N),data2conv8 =>d01_in(2*N-1 downto N),data2conv9 =>d01_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d01_in(9*N-1 downto 8*N),w2 => d01_in(8*N-1 downto 7*N),w3 => d01_in(7*N-1 downto 6*N),w4 => d01_in(6*N-1 downto 5*N),w5 => d01_in(5*N-1 downto 4*N),w6 => d01_in(4*N-1 downto 3*N),w7 => d01_in(3*N-1 downto 2*N),w8 => d01_in(2*N-1 downto N),w9 => d01_in(N-1 downto 0 ),d_out => d01_out,en_out =>en_out,sof_out=>sof_out);
CL02: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d02_in(9*N-1 downto 8*N),data2conv2 =>d02_in(8*N-1 downto 7*N),data2conv3 =>d02_in(7*N-1 downto 6*N),data2conv4 =>d02_in(6*N-1 downto 5*N),data2conv5 =>d02_in(5*N-1 downto 4*N),data2conv6 =>d02_in(4*N-1 downto 3*N),data2conv7 =>d02_in(3*N-1 downto 2*N),data2conv8 =>d02_in(2*N-1 downto N),data2conv9 =>d02_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d02_in(9*N-1 downto 8*N),w2 => d02_in(8*N-1 downto 7*N),w3 => d02_in(7*N-1 downto 6*N),w4 => d02_in(6*N-1 downto 5*N),w5 => d02_in(5*N-1 downto 4*N),w6 => d02_in(4*N-1 downto 3*N),w7 => d02_in(3*N-1 downto 2*N),w8 => d02_in(2*N-1 downto N),w9 => d02_in(N-1 downto 0 ),d_out => d02_out,en_out =>open  ,sof_out=>open   );
CL03: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d03_in(9*N-1 downto 8*N),data2conv2 =>d03_in(8*N-1 downto 7*N),data2conv3 =>d03_in(7*N-1 downto 6*N),data2conv4 =>d03_in(6*N-1 downto 5*N),data2conv5 =>d03_in(5*N-1 downto 4*N),data2conv6 =>d03_in(4*N-1 downto 3*N),data2conv7 =>d03_in(3*N-1 downto 2*N),data2conv8 =>d03_in(2*N-1 downto N),data2conv9 =>d03_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d03_in(9*N-1 downto 8*N),w2 => d03_in(8*N-1 downto 7*N),w3 => d03_in(7*N-1 downto 6*N),w4 => d03_in(6*N-1 downto 5*N),w5 => d03_in(5*N-1 downto 4*N),w6 => d03_in(4*N-1 downto 3*N),w7 => d03_in(3*N-1 downto 2*N),w8 => d03_in(2*N-1 downto N),w9 => d03_in(N-1 downto 0 ),d_out => d03_out,en_out =>open  ,sof_out=>open   );
CL04: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d04_in(9*N-1 downto 8*N),data2conv2 =>d04_in(8*N-1 downto 7*N),data2conv3 =>d04_in(7*N-1 downto 6*N),data2conv4 =>d04_in(6*N-1 downto 5*N),data2conv5 =>d04_in(5*N-1 downto 4*N),data2conv6 =>d04_in(4*N-1 downto 3*N),data2conv7 =>d04_in(3*N-1 downto 2*N),data2conv8 =>d04_in(2*N-1 downto N),data2conv9 =>d04_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d04_in(9*N-1 downto 8*N),w2 => d04_in(8*N-1 downto 7*N),w3 => d04_in(7*N-1 downto 6*N),w4 => d04_in(6*N-1 downto 5*N),w5 => d04_in(5*N-1 downto 4*N),w6 => d04_in(4*N-1 downto 3*N),w7 => d04_in(3*N-1 downto 2*N),w8 => d04_in(2*N-1 downto N),w9 => d04_in(N-1 downto 0 ),d_out => d04_out,en_out =>open  ,sof_out=>open   );
CL05: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d05_in(9*N-1 downto 8*N),data2conv2 =>d05_in(8*N-1 downto 7*N),data2conv3 =>d05_in(7*N-1 downto 6*N),data2conv4 =>d05_in(6*N-1 downto 5*N),data2conv5 =>d05_in(5*N-1 downto 4*N),data2conv6 =>d05_in(4*N-1 downto 3*N),data2conv7 =>d05_in(3*N-1 downto 2*N),data2conv8 =>d05_in(2*N-1 downto N),data2conv9 =>d05_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d05_in(9*N-1 downto 8*N),w2 => d05_in(8*N-1 downto 7*N),w3 => d05_in(7*N-1 downto 6*N),w4 => d05_in(6*N-1 downto 5*N),w5 => d05_in(5*N-1 downto 4*N),w6 => d05_in(4*N-1 downto 3*N),w7 => d05_in(3*N-1 downto 2*N),w8 => d05_in(2*N-1 downto N),w9 => d05_in(N-1 downto 0 ),d_out => d05_out,en_out =>open  ,sof_out=>open   );
CL06: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d06_in(9*N-1 downto 8*N),data2conv2 =>d06_in(8*N-1 downto 7*N),data2conv3 =>d06_in(7*N-1 downto 6*N),data2conv4 =>d06_in(6*N-1 downto 5*N),data2conv5 =>d06_in(5*N-1 downto 4*N),data2conv6 =>d06_in(4*N-1 downto 3*N),data2conv7 =>d06_in(3*N-1 downto 2*N),data2conv8 =>d06_in(2*N-1 downto N),data2conv9 =>d06_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d06_in(9*N-1 downto 8*N),w2 => d06_in(8*N-1 downto 7*N),w3 => d06_in(7*N-1 downto 6*N),w4 => d06_in(6*N-1 downto 5*N),w5 => d06_in(5*N-1 downto 4*N),w6 => d06_in(4*N-1 downto 3*N),w7 => d06_in(3*N-1 downto 2*N),w8 => d06_in(2*N-1 downto N),w9 => d06_in(N-1 downto 0 ),d_out => d06_out,en_out =>open  ,sof_out=>open   );
CL07: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d07_in(9*N-1 downto 8*N),data2conv2 =>d07_in(8*N-1 downto 7*N),data2conv3 =>d07_in(7*N-1 downto 6*N),data2conv4 =>d07_in(6*N-1 downto 5*N),data2conv5 =>d07_in(5*N-1 downto 4*N),data2conv6 =>d07_in(4*N-1 downto 3*N),data2conv7 =>d07_in(3*N-1 downto 2*N),data2conv8 =>d07_in(2*N-1 downto N),data2conv9 =>d07_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d07_in(9*N-1 downto 8*N),w2 => d07_in(8*N-1 downto 7*N),w3 => d07_in(7*N-1 downto 6*N),w4 => d07_in(6*N-1 downto 5*N),w5 => d07_in(5*N-1 downto 4*N),w6 => d07_in(4*N-1 downto 3*N),w7 => d07_in(3*N-1 downto 2*N),w8 => d07_in(2*N-1 downto N),w9 => d07_in(N-1 downto 0 ),d_out => d07_out,en_out =>open  ,sof_out=>open   );
CL08: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d08_in(9*N-1 downto 8*N),data2conv2 =>d08_in(8*N-1 downto 7*N),data2conv3 =>d08_in(7*N-1 downto 6*N),data2conv4 =>d08_in(6*N-1 downto 5*N),data2conv5 =>d08_in(5*N-1 downto 4*N),data2conv6 =>d08_in(4*N-1 downto 3*N),data2conv7 =>d08_in(3*N-1 downto 2*N),data2conv8 =>d08_in(2*N-1 downto N),data2conv9 =>d08_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d08_in(9*N-1 downto 8*N),w2 => d08_in(8*N-1 downto 7*N),w3 => d08_in(7*N-1 downto 6*N),w4 => d08_in(6*N-1 downto 5*N),w5 => d08_in(5*N-1 downto 4*N),w6 => d08_in(4*N-1 downto 3*N),w7 => d08_in(3*N-1 downto 2*N),w8 => d08_in(2*N-1 downto N),w9 => d08_in(N-1 downto 0 ),d_out => d08_out,en_out =>open  ,sof_out=>open   );
CL09: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d09_in(9*N-1 downto 8*N),data2conv2 =>d09_in(8*N-1 downto 7*N),data2conv3 =>d09_in(7*N-1 downto 6*N),data2conv4 =>d09_in(6*N-1 downto 5*N),data2conv5 =>d09_in(5*N-1 downto 4*N),data2conv6 =>d09_in(4*N-1 downto 3*N),data2conv7 =>d09_in(3*N-1 downto 2*N),data2conv8 =>d09_in(2*N-1 downto N),data2conv9 =>d09_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d09_in(9*N-1 downto 8*N),w2 => d09_in(8*N-1 downto 7*N),w3 => d09_in(7*N-1 downto 6*N),w4 => d09_in(6*N-1 downto 5*N),w5 => d09_in(5*N-1 downto 4*N),w6 => d09_in(4*N-1 downto 3*N),w7 => d09_in(3*N-1 downto 2*N),w8 => d09_in(2*N-1 downto N),w9 => d09_in(N-1 downto 0 ),d_out => d09_out,en_out =>open  ,sof_out=>open   );
CL10: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d10_in(9*N-1 downto 8*N),data2conv2 =>d10_in(8*N-1 downto 7*N),data2conv3 =>d10_in(7*N-1 downto 6*N),data2conv4 =>d10_in(6*N-1 downto 5*N),data2conv5 =>d10_in(5*N-1 downto 4*N),data2conv6 =>d10_in(4*N-1 downto 3*N),data2conv7 =>d10_in(3*N-1 downto 2*N),data2conv8 =>d10_in(2*N-1 downto N),data2conv9 =>d10_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d10_in(9*N-1 downto 8*N),w2 => d10_in(8*N-1 downto 7*N),w3 => d10_in(7*N-1 downto 6*N),w4 => d10_in(6*N-1 downto 5*N),w5 => d10_in(5*N-1 downto 4*N),w6 => d10_in(4*N-1 downto 3*N),w7 => d10_in(3*N-1 downto 2*N),w8 => d10_in(2*N-1 downto N),w9 => d10_in(N-1 downto 0 ),d_out => d10_out,en_out =>open  ,sof_out=>open   );
CL11: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d11_in(9*N-1 downto 8*N),data2conv2 =>d11_in(8*N-1 downto 7*N),data2conv3 =>d11_in(7*N-1 downto 6*N),data2conv4 =>d11_in(6*N-1 downto 5*N),data2conv5 =>d11_in(5*N-1 downto 4*N),data2conv6 =>d11_in(4*N-1 downto 3*N),data2conv7 =>d11_in(3*N-1 downto 2*N),data2conv8 =>d11_in(2*N-1 downto N),data2conv9 =>d11_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d11_in(9*N-1 downto 8*N),w2 => d11_in(8*N-1 downto 7*N),w3 => d11_in(7*N-1 downto 6*N),w4 => d11_in(6*N-1 downto 5*N),w5 => d11_in(5*N-1 downto 4*N),w6 => d11_in(4*N-1 downto 3*N),w7 => d11_in(3*N-1 downto 2*N),w8 => d11_in(2*N-1 downto N),w9 => d11_in(N-1 downto 0 ),d_out => d11_out,en_out =>open  ,sof_out=>open   );
CL12: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d12_in(9*N-1 downto 8*N),data2conv2 =>d12_in(8*N-1 downto 7*N),data2conv3 =>d12_in(7*N-1 downto 6*N),data2conv4 =>d12_in(6*N-1 downto 5*N),data2conv5 =>d12_in(5*N-1 downto 4*N),data2conv6 =>d12_in(4*N-1 downto 3*N),data2conv7 =>d12_in(3*N-1 downto 2*N),data2conv8 =>d12_in(2*N-1 downto N),data2conv9 =>d12_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d12_in(9*N-1 downto 8*N),w2 => d12_in(8*N-1 downto 7*N),w3 => d12_in(7*N-1 downto 6*N),w4 => d12_in(6*N-1 downto 5*N),w5 => d12_in(5*N-1 downto 4*N),w6 => d12_in(4*N-1 downto 3*N),w7 => d12_in(3*N-1 downto 2*N),w8 => d12_in(2*N-1 downto N),w9 => d12_in(N-1 downto 0 ),d_out => d12_out,en_out =>open  ,sof_out=>open   );
CL13: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d13_in(9*N-1 downto 8*N),data2conv2 =>d13_in(8*N-1 downto 7*N),data2conv3 =>d13_in(7*N-1 downto 6*N),data2conv4 =>d13_in(6*N-1 downto 5*N),data2conv5 =>d13_in(5*N-1 downto 4*N),data2conv6 =>d13_in(4*N-1 downto 3*N),data2conv7 =>d13_in(3*N-1 downto 2*N),data2conv8 =>d13_in(2*N-1 downto N),data2conv9 =>d13_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d13_in(9*N-1 downto 8*N),w2 => d13_in(8*N-1 downto 7*N),w3 => d13_in(7*N-1 downto 6*N),w4 => d13_in(6*N-1 downto 5*N),w5 => d13_in(5*N-1 downto 4*N),w6 => d13_in(4*N-1 downto 3*N),w7 => d13_in(3*N-1 downto 2*N),w8 => d13_in(2*N-1 downto N),w9 => d13_in(N-1 downto 0 ),d_out => d13_out,en_out =>open  ,sof_out=>open   );
CL14: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d14_in(9*N-1 downto 8*N),data2conv2 =>d14_in(8*N-1 downto 7*N),data2conv3 =>d14_in(7*N-1 downto 6*N),data2conv4 =>d14_in(6*N-1 downto 5*N),data2conv5 =>d14_in(5*N-1 downto 4*N),data2conv6 =>d14_in(4*N-1 downto 3*N),data2conv7 =>d14_in(3*N-1 downto 2*N),data2conv8 =>d14_in(2*N-1 downto N),data2conv9 =>d14_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d14_in(9*N-1 downto 8*N),w2 => d14_in(8*N-1 downto 7*N),w3 => d14_in(7*N-1 downto 6*N),w4 => d14_in(6*N-1 downto 5*N),w5 => d14_in(5*N-1 downto 4*N),w6 => d14_in(4*N-1 downto 3*N),w7 => d14_in(3*N-1 downto 2*N),w8 => d14_in(2*N-1 downto N),w9 => d14_in(N-1 downto 0 ),d_out => d14_out,en_out =>open  ,sof_out=>open   );
CL15: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d15_in(9*N-1 downto 8*N),data2conv2 =>d15_in(8*N-1 downto 7*N),data2conv3 =>d15_in(7*N-1 downto 6*N),data2conv4 =>d15_in(6*N-1 downto 5*N),data2conv5 =>d15_in(5*N-1 downto 4*N),data2conv6 =>d15_in(4*N-1 downto 3*N),data2conv7 =>d15_in(3*N-1 downto 2*N),data2conv8 =>d15_in(2*N-1 downto N),data2conv9 =>d15_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d15_in(9*N-1 downto 8*N),w2 => d15_in(8*N-1 downto 7*N),w3 => d15_in(7*N-1 downto 6*N),w4 => d15_in(6*N-1 downto 5*N),w5 => d15_in(5*N-1 downto 4*N),w6 => d15_in(4*N-1 downto 3*N),w7 => d15_in(3*N-1 downto 2*N),w8 => d15_in(2*N-1 downto N),w9 => d15_in(N-1 downto 0 ),d_out => d15_out,en_out =>open  ,sof_out=>open   );
CL16: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d16_in(9*N-1 downto 8*N),data2conv2 =>d16_in(8*N-1 downto 7*N),data2conv3 =>d16_in(7*N-1 downto 6*N),data2conv4 =>d16_in(6*N-1 downto 5*N),data2conv5 =>d16_in(5*N-1 downto 4*N),data2conv6 =>d16_in(4*N-1 downto 3*N),data2conv7 =>d16_in(3*N-1 downto 2*N),data2conv8 =>d16_in(2*N-1 downto N),data2conv9 =>d16_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d16_in(9*N-1 downto 8*N),w2 => d16_in(8*N-1 downto 7*N),w3 => d16_in(7*N-1 downto 6*N),w4 => d16_in(6*N-1 downto 5*N),w5 => d16_in(5*N-1 downto 4*N),w6 => d16_in(4*N-1 downto 3*N),w7 => d16_in(3*N-1 downto 2*N),w8 => d16_in(2*N-1 downto N),w9 => d16_in(N-1 downto 0 ),d_out => d16_out,en_out =>open  ,sof_out=>open   );
CL17: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d17_in(9*N-1 downto 8*N),data2conv2 =>d17_in(8*N-1 downto 7*N),data2conv3 =>d17_in(7*N-1 downto 6*N),data2conv4 =>d17_in(6*N-1 downto 5*N),data2conv5 =>d17_in(5*N-1 downto 4*N),data2conv6 =>d17_in(4*N-1 downto 3*N),data2conv7 =>d17_in(3*N-1 downto 2*N),data2conv8 =>d17_in(2*N-1 downto N),data2conv9 =>d17_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d17_in(9*N-1 downto 8*N),w2 => d17_in(8*N-1 downto 7*N),w3 => d17_in(7*N-1 downto 6*N),w4 => d17_in(6*N-1 downto 5*N),w5 => d17_in(5*N-1 downto 4*N),w6 => d17_in(4*N-1 downto 3*N),w7 => d17_in(3*N-1 downto 2*N),w8 => d17_in(2*N-1 downto N),w9 => d17_in(N-1 downto 0 ),d_out => d17_out,en_out =>open  ,sof_out=>open   );
CL18: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d18_in(9*N-1 downto 8*N),data2conv2 =>d18_in(8*N-1 downto 7*N),data2conv3 =>d18_in(7*N-1 downto 6*N),data2conv4 =>d18_in(6*N-1 downto 5*N),data2conv5 =>d18_in(5*N-1 downto 4*N),data2conv6 =>d18_in(4*N-1 downto 3*N),data2conv7 =>d18_in(3*N-1 downto 2*N),data2conv8 =>d18_in(2*N-1 downto N),data2conv9 =>d18_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d18_in(9*N-1 downto 8*N),w2 => d18_in(8*N-1 downto 7*N),w3 => d18_in(7*N-1 downto 6*N),w4 => d18_in(6*N-1 downto 5*N),w5 => d18_in(5*N-1 downto 4*N),w6 => d18_in(4*N-1 downto 3*N),w7 => d18_in(3*N-1 downto 2*N),w8 => d18_in(2*N-1 downto N),w9 => d18_in(N-1 downto 0 ),d_out => d18_out,en_out =>open  ,sof_out=>open   );
CL19: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d19_in(9*N-1 downto 8*N),data2conv2 =>d19_in(8*N-1 downto 7*N),data2conv3 =>d19_in(7*N-1 downto 6*N),data2conv4 =>d19_in(6*N-1 downto 5*N),data2conv5 =>d19_in(5*N-1 downto 4*N),data2conv6 =>d19_in(4*N-1 downto 3*N),data2conv7 =>d19_in(3*N-1 downto 2*N),data2conv8 =>d19_in(2*N-1 downto N),data2conv9 =>d19_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d19_in(9*N-1 downto 8*N),w2 => d19_in(8*N-1 downto 7*N),w3 => d19_in(7*N-1 downto 6*N),w4 => d19_in(6*N-1 downto 5*N),w5 => d19_in(5*N-1 downto 4*N),w6 => d19_in(4*N-1 downto 3*N),w7 => d19_in(3*N-1 downto 2*N),w8 => d19_in(2*N-1 downto N),w9 => d19_in(N-1 downto 0 ),d_out => d19_out,en_out =>open  ,sof_out=>open   );
CL20: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d20_in(9*N-1 downto 8*N),data2conv2 =>d20_in(8*N-1 downto 7*N),data2conv3 =>d20_in(7*N-1 downto 6*N),data2conv4 =>d20_in(6*N-1 downto 5*N),data2conv5 =>d20_in(5*N-1 downto 4*N),data2conv6 =>d20_in(4*N-1 downto 3*N),data2conv7 =>d20_in(3*N-1 downto 2*N),data2conv8 =>d20_in(2*N-1 downto N),data2conv9 =>d20_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d20_in(9*N-1 downto 8*N),w2 => d20_in(8*N-1 downto 7*N),w3 => d20_in(7*N-1 downto 6*N),w4 => d20_in(6*N-1 downto 5*N),w5 => d20_in(5*N-1 downto 4*N),w6 => d20_in(4*N-1 downto 3*N),w7 => d20_in(3*N-1 downto 2*N),w8 => d20_in(2*N-1 downto N),w9 => d20_in(N-1 downto 0 ),d_out => d20_out,en_out =>open  ,sof_out=>open   );
CL21: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d21_in(9*N-1 downto 8*N),data2conv2 =>d21_in(8*N-1 downto 7*N),data2conv3 =>d21_in(7*N-1 downto 6*N),data2conv4 =>d21_in(6*N-1 downto 5*N),data2conv5 =>d21_in(5*N-1 downto 4*N),data2conv6 =>d21_in(4*N-1 downto 3*N),data2conv7 =>d21_in(3*N-1 downto 2*N),data2conv8 =>d21_in(2*N-1 downto N),data2conv9 =>d21_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d21_in(9*N-1 downto 8*N),w2 => d21_in(8*N-1 downto 7*N),w3 => d21_in(7*N-1 downto 6*N),w4 => d21_in(6*N-1 downto 5*N),w5 => d21_in(5*N-1 downto 4*N),w6 => d21_in(4*N-1 downto 3*N),w7 => d21_in(3*N-1 downto 2*N),w8 => d21_in(2*N-1 downto N),w9 => d21_in(N-1 downto 0 ),d_out => d21_out,en_out =>open  ,sof_out=>open   );
CL22: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d22_in(9*N-1 downto 8*N),data2conv2 =>d22_in(8*N-1 downto 7*N),data2conv3 =>d22_in(7*N-1 downto 6*N),data2conv4 =>d22_in(6*N-1 downto 5*N),data2conv5 =>d22_in(5*N-1 downto 4*N),data2conv6 =>d22_in(4*N-1 downto 3*N),data2conv7 =>d22_in(3*N-1 downto 2*N),data2conv8 =>d22_in(2*N-1 downto N),data2conv9 =>d22_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d22_in(9*N-1 downto 8*N),w2 => d22_in(8*N-1 downto 7*N),w3 => d22_in(7*N-1 downto 6*N),w4 => d22_in(6*N-1 downto 5*N),w5 => d22_in(5*N-1 downto 4*N),w6 => d22_in(4*N-1 downto 3*N),w7 => d22_in(3*N-1 downto 2*N),w8 => d22_in(2*N-1 downto N),w9 => d22_in(N-1 downto 0 ),d_out => d22_out,en_out =>open  ,sof_out=>open   );
CL23: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d23_in(9*N-1 downto 8*N),data2conv2 =>d23_in(8*N-1 downto 7*N),data2conv3 =>d23_in(7*N-1 downto 6*N),data2conv4 =>d23_in(6*N-1 downto 5*N),data2conv5 =>d23_in(5*N-1 downto 4*N),data2conv6 =>d23_in(4*N-1 downto 3*N),data2conv7 =>d23_in(3*N-1 downto 2*N),data2conv8 =>d23_in(2*N-1 downto N),data2conv9 =>d23_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d23_in(9*N-1 downto 8*N),w2 => d23_in(8*N-1 downto 7*N),w3 => d23_in(7*N-1 downto 6*N),w4 => d23_in(6*N-1 downto 5*N),w5 => d23_in(5*N-1 downto 4*N),w6 => d23_in(4*N-1 downto 3*N),w7 => d23_in(3*N-1 downto 2*N),w8 => d23_in(2*N-1 downto N),w9 => d23_in(N-1 downto 0 ),d_out => d23_out,en_out =>open  ,sof_out=>open   );
CL24: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d24_in(9*N-1 downto 8*N),data2conv2 =>d24_in(8*N-1 downto 7*N),data2conv3 =>d24_in(7*N-1 downto 6*N),data2conv4 =>d24_in(6*N-1 downto 5*N),data2conv5 =>d24_in(5*N-1 downto 4*N),data2conv6 =>d24_in(4*N-1 downto 3*N),data2conv7 =>d24_in(3*N-1 downto 2*N),data2conv8 =>d24_in(2*N-1 downto N),data2conv9 =>d24_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d24_in(9*N-1 downto 8*N),w2 => d24_in(8*N-1 downto 7*N),w3 => d24_in(7*N-1 downto 6*N),w4 => d24_in(6*N-1 downto 5*N),w5 => d24_in(5*N-1 downto 4*N),w6 => d24_in(4*N-1 downto 3*N),w7 => d24_in(3*N-1 downto 2*N),w8 => d24_in(2*N-1 downto N),w9 => d24_in(N-1 downto 0 ),d_out => d24_out,en_out =>open  ,sof_out=>open   );
CL25: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d25_in(9*N-1 downto 8*N),data2conv2 =>d25_in(8*N-1 downto 7*N),data2conv3 =>d25_in(7*N-1 downto 6*N),data2conv4 =>d25_in(6*N-1 downto 5*N),data2conv5 =>d25_in(5*N-1 downto 4*N),data2conv6 =>d25_in(4*N-1 downto 3*N),data2conv7 =>d25_in(3*N-1 downto 2*N),data2conv8 =>d25_in(2*N-1 downto N),data2conv9 =>d25_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d25_in(9*N-1 downto 8*N),w2 => d25_in(8*N-1 downto 7*N),w3 => d25_in(7*N-1 downto 6*N),w4 => d25_in(6*N-1 downto 5*N),w5 => d25_in(5*N-1 downto 4*N),w6 => d25_in(4*N-1 downto 3*N),w7 => d25_in(3*N-1 downto 2*N),w8 => d25_in(2*N-1 downto N),w9 => d25_in(N-1 downto 0 ),d_out => d25_out,en_out =>open  ,sof_out=>open   );
CL26: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d26_in(9*N-1 downto 8*N),data2conv2 =>d26_in(8*N-1 downto 7*N),data2conv3 =>d26_in(7*N-1 downto 6*N),data2conv4 =>d26_in(6*N-1 downto 5*N),data2conv5 =>d26_in(5*N-1 downto 4*N),data2conv6 =>d26_in(4*N-1 downto 3*N),data2conv7 =>d26_in(3*N-1 downto 2*N),data2conv8 =>d26_in(2*N-1 downto N),data2conv9 =>d26_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d26_in(9*N-1 downto 8*N),w2 => d26_in(8*N-1 downto 7*N),w3 => d26_in(7*N-1 downto 6*N),w4 => d26_in(6*N-1 downto 5*N),w5 => d26_in(5*N-1 downto 4*N),w6 => d26_in(4*N-1 downto 3*N),w7 => d26_in(3*N-1 downto 2*N),w8 => d26_in(2*N-1 downto N),w9 => d26_in(N-1 downto 0 ),d_out => d26_out,en_out =>open  ,sof_out=>open   );
CL27: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d27_in(9*N-1 downto 8*N),data2conv2 =>d27_in(8*N-1 downto 7*N),data2conv3 =>d27_in(7*N-1 downto 6*N),data2conv4 =>d27_in(6*N-1 downto 5*N),data2conv5 =>d27_in(5*N-1 downto 4*N),data2conv6 =>d27_in(4*N-1 downto 3*N),data2conv7 =>d27_in(3*N-1 downto 2*N),data2conv8 =>d27_in(2*N-1 downto N),data2conv9 =>d27_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d27_in(9*N-1 downto 8*N),w2 => d27_in(8*N-1 downto 7*N),w3 => d27_in(7*N-1 downto 6*N),w4 => d27_in(6*N-1 downto 5*N),w5 => d27_in(5*N-1 downto 4*N),w6 => d27_in(4*N-1 downto 3*N),w7 => d27_in(3*N-1 downto 2*N),w8 => d27_in(2*N-1 downto N),w9 => d27_in(N-1 downto 0 ),d_out => d27_out,en_out =>open  ,sof_out=>open   );
CL28: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d28_in(9*N-1 downto 8*N),data2conv2 =>d28_in(8*N-1 downto 7*N),data2conv3 =>d28_in(7*N-1 downto 6*N),data2conv4 =>d28_in(6*N-1 downto 5*N),data2conv5 =>d28_in(5*N-1 downto 4*N),data2conv6 =>d28_in(4*N-1 downto 3*N),data2conv7 =>d28_in(3*N-1 downto 2*N),data2conv8 =>d28_in(2*N-1 downto N),data2conv9 =>d28_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d28_in(9*N-1 downto 8*N),w2 => d28_in(8*N-1 downto 7*N),w3 => d28_in(7*N-1 downto 6*N),w4 => d28_in(6*N-1 downto 5*N),w5 => d28_in(5*N-1 downto 4*N),w6 => d28_in(4*N-1 downto 3*N),w7 => d28_in(3*N-1 downto 2*N),w8 => d28_in(2*N-1 downto N),w9 => d28_in(N-1 downto 0 ),d_out => d28_out,en_out =>open  ,sof_out=>open   );
CL29: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d29_in(9*N-1 downto 8*N),data2conv2 =>d29_in(8*N-1 downto 7*N),data2conv3 =>d29_in(7*N-1 downto 6*N),data2conv4 =>d29_in(6*N-1 downto 5*N),data2conv5 =>d29_in(5*N-1 downto 4*N),data2conv6 =>d29_in(4*N-1 downto 3*N),data2conv7 =>d29_in(3*N-1 downto 2*N),data2conv8 =>d29_in(2*N-1 downto N),data2conv9 =>d29_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d29_in(9*N-1 downto 8*N),w2 => d29_in(8*N-1 downto 7*N),w3 => d29_in(7*N-1 downto 6*N),w4 => d29_in(6*N-1 downto 5*N),w5 => d29_in(5*N-1 downto 4*N),w6 => d29_in(4*N-1 downto 3*N),w7 => d29_in(3*N-1 downto 2*N),w8 => d29_in(2*N-1 downto N),w9 => d29_in(N-1 downto 0 ),d_out => d29_out,en_out =>open  ,sof_out=>open   );
CL30: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d30_in(9*N-1 downto 8*N),data2conv2 =>d30_in(8*N-1 downto 7*N),data2conv3 =>d30_in(7*N-1 downto 6*N),data2conv4 =>d30_in(6*N-1 downto 5*N),data2conv5 =>d30_in(5*N-1 downto 4*N),data2conv6 =>d30_in(4*N-1 downto 3*N),data2conv7 =>d30_in(3*N-1 downto 2*N),data2conv8 =>d30_in(2*N-1 downto N),data2conv9 =>d30_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d30_in(9*N-1 downto 8*N),w2 => d30_in(8*N-1 downto 7*N),w3 => d30_in(7*N-1 downto 6*N),w4 => d30_in(6*N-1 downto 5*N),w5 => d30_in(5*N-1 downto 4*N),w6 => d30_in(4*N-1 downto 3*N),w7 => d30_in(3*N-1 downto 2*N),w8 => d30_in(2*N-1 downto N),w9 => d30_in(N-1 downto 0 ),d_out => d30_out,en_out =>open  ,sof_out=>open   );
CL31: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d31_in(9*N-1 downto 8*N),data2conv2 =>d31_in(8*N-1 downto 7*N),data2conv3 =>d31_in(7*N-1 downto 6*N),data2conv4 =>d31_in(6*N-1 downto 5*N),data2conv5 =>d31_in(5*N-1 downto 4*N),data2conv6 =>d31_in(4*N-1 downto 3*N),data2conv7 =>d31_in(3*N-1 downto 2*N),data2conv8 =>d31_in(2*N-1 downto N),data2conv9 =>d31_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d31_in(9*N-1 downto 8*N),w2 => d31_in(8*N-1 downto 7*N),w3 => d31_in(7*N-1 downto 6*N),w4 => d31_in(6*N-1 downto 5*N),w5 => d31_in(5*N-1 downto 4*N),w6 => d31_in(4*N-1 downto 3*N),w7 => d31_in(3*N-1 downto 2*N),w8 => d31_in(2*N-1 downto N),w9 => d31_in(N-1 downto 0 ),d_out => d31_out,en_out =>open  ,sof_out=>open   );
CL32: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d32_in(9*N-1 downto 8*N),data2conv2 =>d32_in(8*N-1 downto 7*N),data2conv3 =>d32_in(7*N-1 downto 6*N),data2conv4 =>d32_in(6*N-1 downto 5*N),data2conv5 =>d32_in(5*N-1 downto 4*N),data2conv6 =>d32_in(4*N-1 downto 3*N),data2conv7 =>d32_in(3*N-1 downto 2*N),data2conv8 =>d32_in(2*N-1 downto N),data2conv9 =>d32_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d32_in(9*N-1 downto 8*N),w2 => d32_in(8*N-1 downto 7*N),w3 => d32_in(7*N-1 downto 6*N),w4 => d32_in(6*N-1 downto 5*N),w5 => d32_in(5*N-1 downto 4*N),w6 => d32_in(4*N-1 downto 3*N),w7 => d32_in(3*N-1 downto 2*N),w8 => d32_in(2*N-1 downto N),w9 => d32_in(N-1 downto 0 ),d_out => d32_out,en_out =>open  ,sof_out=>open   );
CL33: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d33_in(9*N-1 downto 8*N),data2conv2 =>d33_in(8*N-1 downto 7*N),data2conv3 =>d33_in(7*N-1 downto 6*N),data2conv4 =>d33_in(6*N-1 downto 5*N),data2conv5 =>d33_in(5*N-1 downto 4*N),data2conv6 =>d33_in(4*N-1 downto 3*N),data2conv7 =>d33_in(3*N-1 downto 2*N),data2conv8 =>d33_in(2*N-1 downto N),data2conv9 =>d33_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d33_in(9*N-1 downto 8*N),w2 => d33_in(8*N-1 downto 7*N),w3 => d33_in(7*N-1 downto 6*N),w4 => d33_in(6*N-1 downto 5*N),w5 => d33_in(5*N-1 downto 4*N),w6 => d33_in(4*N-1 downto 3*N),w7 => d33_in(3*N-1 downto 2*N),w8 => d33_in(2*N-1 downto N),w9 => d33_in(N-1 downto 0 ),d_out => d33_out,en_out =>open  ,sof_out=>open   );
CL34: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d34_in(9*N-1 downto 8*N),data2conv2 =>d34_in(8*N-1 downto 7*N),data2conv3 =>d34_in(7*N-1 downto 6*N),data2conv4 =>d34_in(6*N-1 downto 5*N),data2conv5 =>d34_in(5*N-1 downto 4*N),data2conv6 =>d34_in(4*N-1 downto 3*N),data2conv7 =>d34_in(3*N-1 downto 2*N),data2conv8 =>d34_in(2*N-1 downto N),data2conv9 =>d34_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d34_in(9*N-1 downto 8*N),w2 => d34_in(8*N-1 downto 7*N),w3 => d34_in(7*N-1 downto 6*N),w4 => d34_in(6*N-1 downto 5*N),w5 => d34_in(5*N-1 downto 4*N),w6 => d34_in(4*N-1 downto 3*N),w7 => d34_in(3*N-1 downto 2*N),w8 => d34_in(2*N-1 downto N),w9 => d34_in(N-1 downto 0 ),d_out => d34_out,en_out =>open  ,sof_out=>open   );
CL35: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d35_in(9*N-1 downto 8*N),data2conv2 =>d35_in(8*N-1 downto 7*N),data2conv3 =>d35_in(7*N-1 downto 6*N),data2conv4 =>d35_in(6*N-1 downto 5*N),data2conv5 =>d35_in(5*N-1 downto 4*N),data2conv6 =>d35_in(4*N-1 downto 3*N),data2conv7 =>d35_in(3*N-1 downto 2*N),data2conv8 =>d35_in(2*N-1 downto N),data2conv9 =>d35_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d35_in(9*N-1 downto 8*N),w2 => d35_in(8*N-1 downto 7*N),w3 => d35_in(7*N-1 downto 6*N),w4 => d35_in(6*N-1 downto 5*N),w5 => d35_in(5*N-1 downto 4*N),w6 => d35_in(4*N-1 downto 3*N),w7 => d35_in(3*N-1 downto 2*N),w8 => d35_in(2*N-1 downto N),w9 => d35_in(N-1 downto 0 ),d_out => d35_out,en_out =>open  ,sof_out=>open   );
CL36: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d36_in(9*N-1 downto 8*N),data2conv2 =>d36_in(8*N-1 downto 7*N),data2conv3 =>d36_in(7*N-1 downto 6*N),data2conv4 =>d36_in(6*N-1 downto 5*N),data2conv5 =>d36_in(5*N-1 downto 4*N),data2conv6 =>d36_in(4*N-1 downto 3*N),data2conv7 =>d36_in(3*N-1 downto 2*N),data2conv8 =>d36_in(2*N-1 downto N),data2conv9 =>d36_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d36_in(9*N-1 downto 8*N),w2 => d36_in(8*N-1 downto 7*N),w3 => d36_in(7*N-1 downto 6*N),w4 => d36_in(6*N-1 downto 5*N),w5 => d36_in(5*N-1 downto 4*N),w6 => d36_in(4*N-1 downto 3*N),w7 => d36_in(3*N-1 downto 2*N),w8 => d36_in(2*N-1 downto N),w9 => d36_in(N-1 downto 0 ),d_out => d36_out,en_out =>open  ,sof_out=>open   );
CL37: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d37_in(9*N-1 downto 8*N),data2conv2 =>d37_in(8*N-1 downto 7*N),data2conv3 =>d37_in(7*N-1 downto 6*N),data2conv4 =>d37_in(6*N-1 downto 5*N),data2conv5 =>d37_in(5*N-1 downto 4*N),data2conv6 =>d37_in(4*N-1 downto 3*N),data2conv7 =>d37_in(3*N-1 downto 2*N),data2conv8 =>d37_in(2*N-1 downto N),data2conv9 =>d37_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d37_in(9*N-1 downto 8*N),w2 => d37_in(8*N-1 downto 7*N),w3 => d37_in(7*N-1 downto 6*N),w4 => d37_in(6*N-1 downto 5*N),w5 => d37_in(5*N-1 downto 4*N),w6 => d37_in(4*N-1 downto 3*N),w7 => d37_in(3*N-1 downto 2*N),w8 => d37_in(2*N-1 downto N),w9 => d37_in(N-1 downto 0 ),d_out => d37_out,en_out =>open  ,sof_out=>open   );
CL38: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d38_in(9*N-1 downto 8*N),data2conv2 =>d38_in(8*N-1 downto 7*N),data2conv3 =>d38_in(7*N-1 downto 6*N),data2conv4 =>d38_in(6*N-1 downto 5*N),data2conv5 =>d38_in(5*N-1 downto 4*N),data2conv6 =>d38_in(4*N-1 downto 3*N),data2conv7 =>d38_in(3*N-1 downto 2*N),data2conv8 =>d38_in(2*N-1 downto N),data2conv9 =>d38_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d38_in(9*N-1 downto 8*N),w2 => d38_in(8*N-1 downto 7*N),w3 => d38_in(7*N-1 downto 6*N),w4 => d38_in(6*N-1 downto 5*N),w5 => d38_in(5*N-1 downto 4*N),w6 => d38_in(4*N-1 downto 3*N),w7 => d38_in(3*N-1 downto 2*N),w8 => d38_in(2*N-1 downto N),w9 => d38_in(N-1 downto 0 ),d_out => d38_out,en_out =>open  ,sof_out=>open   );
CL39: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d39_in(9*N-1 downto 8*N),data2conv2 =>d39_in(8*N-1 downto 7*N),data2conv3 =>d39_in(7*N-1 downto 6*N),data2conv4 =>d39_in(6*N-1 downto 5*N),data2conv5 =>d39_in(5*N-1 downto 4*N),data2conv6 =>d39_in(4*N-1 downto 3*N),data2conv7 =>d39_in(3*N-1 downto 2*N),data2conv8 =>d39_in(2*N-1 downto N),data2conv9 =>d39_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d39_in(9*N-1 downto 8*N),w2 => d39_in(8*N-1 downto 7*N),w3 => d39_in(7*N-1 downto 6*N),w4 => d39_in(6*N-1 downto 5*N),w5 => d39_in(5*N-1 downto 4*N),w6 => d39_in(4*N-1 downto 3*N),w7 => d39_in(3*N-1 downto 2*N),w8 => d39_in(2*N-1 downto N),w9 => d39_in(N-1 downto 0 ),d_out => d39_out,en_out =>open  ,sof_out=>open   );
CL40: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d40_in(9*N-1 downto 8*N),data2conv2 =>d40_in(8*N-1 downto 7*N),data2conv3 =>d40_in(7*N-1 downto 6*N),data2conv4 =>d40_in(6*N-1 downto 5*N),data2conv5 =>d40_in(5*N-1 downto 4*N),data2conv6 =>d40_in(4*N-1 downto 3*N),data2conv7 =>d40_in(3*N-1 downto 2*N),data2conv8 =>d40_in(2*N-1 downto N),data2conv9 =>d40_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d40_in(9*N-1 downto 8*N),w2 => d40_in(8*N-1 downto 7*N),w3 => d40_in(7*N-1 downto 6*N),w4 => d40_in(6*N-1 downto 5*N),w5 => d40_in(5*N-1 downto 4*N),w6 => d40_in(4*N-1 downto 3*N),w7 => d40_in(3*N-1 downto 2*N),w8 => d40_in(2*N-1 downto N),w9 => d40_in(N-1 downto 0 ),d_out => d40_out,en_out =>open  ,sof_out=>open   );
CL41: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d41_in(9*N-1 downto 8*N),data2conv2 =>d41_in(8*N-1 downto 7*N),data2conv3 =>d41_in(7*N-1 downto 6*N),data2conv4 =>d41_in(6*N-1 downto 5*N),data2conv5 =>d41_in(5*N-1 downto 4*N),data2conv6 =>d41_in(4*N-1 downto 3*N),data2conv7 =>d41_in(3*N-1 downto 2*N),data2conv8 =>d41_in(2*N-1 downto N),data2conv9 =>d41_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d41_in(9*N-1 downto 8*N),w2 => d41_in(8*N-1 downto 7*N),w3 => d41_in(7*N-1 downto 6*N),w4 => d41_in(6*N-1 downto 5*N),w5 => d41_in(5*N-1 downto 4*N),w6 => d41_in(4*N-1 downto 3*N),w7 => d41_in(3*N-1 downto 2*N),w8 => d41_in(2*N-1 downto N),w9 => d41_in(N-1 downto 0 ),d_out => d41_out,en_out =>open  ,sof_out=>open   );
CL42: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d42_in(9*N-1 downto 8*N),data2conv2 =>d42_in(8*N-1 downto 7*N),data2conv3 =>d42_in(7*N-1 downto 6*N),data2conv4 =>d42_in(6*N-1 downto 5*N),data2conv5 =>d42_in(5*N-1 downto 4*N),data2conv6 =>d42_in(4*N-1 downto 3*N),data2conv7 =>d42_in(3*N-1 downto 2*N),data2conv8 =>d42_in(2*N-1 downto N),data2conv9 =>d42_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d42_in(9*N-1 downto 8*N),w2 => d42_in(8*N-1 downto 7*N),w3 => d42_in(7*N-1 downto 6*N),w4 => d42_in(6*N-1 downto 5*N),w5 => d42_in(5*N-1 downto 4*N),w6 => d42_in(4*N-1 downto 3*N),w7 => d42_in(3*N-1 downto 2*N),w8 => d42_in(2*N-1 downto N),w9 => d42_in(N-1 downto 0 ),d_out => d42_out,en_out =>open  ,sof_out=>open   );
CL43: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d43_in(9*N-1 downto 8*N),data2conv2 =>d43_in(8*N-1 downto 7*N),data2conv3 =>d43_in(7*N-1 downto 6*N),data2conv4 =>d43_in(6*N-1 downto 5*N),data2conv5 =>d43_in(5*N-1 downto 4*N),data2conv6 =>d43_in(4*N-1 downto 3*N),data2conv7 =>d43_in(3*N-1 downto 2*N),data2conv8 =>d43_in(2*N-1 downto N),data2conv9 =>d43_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d43_in(9*N-1 downto 8*N),w2 => d43_in(8*N-1 downto 7*N),w3 => d43_in(7*N-1 downto 6*N),w4 => d43_in(6*N-1 downto 5*N),w5 => d43_in(5*N-1 downto 4*N),w6 => d43_in(4*N-1 downto 3*N),w7 => d43_in(3*N-1 downto 2*N),w8 => d43_in(2*N-1 downto N),w9 => d43_in(N-1 downto 0 ),d_out => d43_out,en_out =>open  ,sof_out=>open   );
CL44: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d44_in(9*N-1 downto 8*N),data2conv2 =>d44_in(8*N-1 downto 7*N),data2conv3 =>d44_in(7*N-1 downto 6*N),data2conv4 =>d44_in(6*N-1 downto 5*N),data2conv5 =>d44_in(5*N-1 downto 4*N),data2conv6 =>d44_in(4*N-1 downto 3*N),data2conv7 =>d44_in(3*N-1 downto 2*N),data2conv8 =>d44_in(2*N-1 downto N),data2conv9 =>d44_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d44_in(9*N-1 downto 8*N),w2 => d44_in(8*N-1 downto 7*N),w3 => d44_in(7*N-1 downto 6*N),w4 => d44_in(6*N-1 downto 5*N),w5 => d44_in(5*N-1 downto 4*N),w6 => d44_in(4*N-1 downto 3*N),w7 => d44_in(3*N-1 downto 2*N),w8 => d44_in(2*N-1 downto N),w9 => d44_in(N-1 downto 0 ),d_out => d44_out,en_out =>open  ,sof_out=>open   );
CL45: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d45_in(9*N-1 downto 8*N),data2conv2 =>d45_in(8*N-1 downto 7*N),data2conv3 =>d45_in(7*N-1 downto 6*N),data2conv4 =>d45_in(6*N-1 downto 5*N),data2conv5 =>d45_in(5*N-1 downto 4*N),data2conv6 =>d45_in(4*N-1 downto 3*N),data2conv7 =>d45_in(3*N-1 downto 2*N),data2conv8 =>d45_in(2*N-1 downto N),data2conv9 =>d45_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d45_in(9*N-1 downto 8*N),w2 => d45_in(8*N-1 downto 7*N),w3 => d45_in(7*N-1 downto 6*N),w4 => d45_in(6*N-1 downto 5*N),w5 => d45_in(5*N-1 downto 4*N),w6 => d45_in(4*N-1 downto 3*N),w7 => d45_in(3*N-1 downto 2*N),w8 => d45_in(2*N-1 downto N),w9 => d45_in(N-1 downto 0 ),d_out => d45_out,en_out =>open  ,sof_out=>open   );
CL46: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d46_in(9*N-1 downto 8*N),data2conv2 =>d46_in(8*N-1 downto 7*N),data2conv3 =>d46_in(7*N-1 downto 6*N),data2conv4 =>d46_in(6*N-1 downto 5*N),data2conv5 =>d46_in(5*N-1 downto 4*N),data2conv6 =>d46_in(4*N-1 downto 3*N),data2conv7 =>d46_in(3*N-1 downto 2*N),data2conv8 =>d46_in(2*N-1 downto N),data2conv9 =>d46_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d46_in(9*N-1 downto 8*N),w2 => d46_in(8*N-1 downto 7*N),w3 => d46_in(7*N-1 downto 6*N),w4 => d46_in(6*N-1 downto 5*N),w5 => d46_in(5*N-1 downto 4*N),w6 => d46_in(4*N-1 downto 3*N),w7 => d46_in(3*N-1 downto 2*N),w8 => d46_in(2*N-1 downto N),w9 => d46_in(N-1 downto 0 ),d_out => d46_out,en_out =>open  ,sof_out=>open   );
CL47: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d47_in(9*N-1 downto 8*N),data2conv2 =>d47_in(8*N-1 downto 7*N),data2conv3 =>d47_in(7*N-1 downto 6*N),data2conv4 =>d47_in(6*N-1 downto 5*N),data2conv5 =>d47_in(5*N-1 downto 4*N),data2conv6 =>d47_in(4*N-1 downto 3*N),data2conv7 =>d47_in(3*N-1 downto 2*N),data2conv8 =>d47_in(2*N-1 downto N),data2conv9 =>d47_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d47_in(9*N-1 downto 8*N),w2 => d47_in(8*N-1 downto 7*N),w3 => d47_in(7*N-1 downto 6*N),w4 => d47_in(6*N-1 downto 5*N),w5 => d47_in(5*N-1 downto 4*N),w6 => d47_in(4*N-1 downto 3*N),w7 => d47_in(3*N-1 downto 2*N),w8 => d47_in(2*N-1 downto N),w9 => d47_in(N-1 downto 0 ),d_out => d47_out,en_out =>open  ,sof_out=>open   );
CL48: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d48_in(9*N-1 downto 8*N),data2conv2 =>d48_in(8*N-1 downto 7*N),data2conv3 =>d48_in(7*N-1 downto 6*N),data2conv4 =>d48_in(6*N-1 downto 5*N),data2conv5 =>d48_in(5*N-1 downto 4*N),data2conv6 =>d48_in(4*N-1 downto 3*N),data2conv7 =>d48_in(3*N-1 downto 2*N),data2conv8 =>d48_in(2*N-1 downto N),data2conv9 =>d48_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d48_in(9*N-1 downto 8*N),w2 => d48_in(8*N-1 downto 7*N),w3 => d48_in(7*N-1 downto 6*N),w4 => d48_in(6*N-1 downto 5*N),w5 => d48_in(5*N-1 downto 4*N),w6 => d48_in(4*N-1 downto 3*N),w7 => d48_in(3*N-1 downto 2*N),w8 => d48_in(2*N-1 downto N),w9 => d48_in(N-1 downto 0 ),d_out => d48_out,en_out =>open  ,sof_out=>open   );
CL49: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d49_in(9*N-1 downto 8*N),data2conv2 =>d49_in(8*N-1 downto 7*N),data2conv3 =>d49_in(7*N-1 downto 6*N),data2conv4 =>d49_in(6*N-1 downto 5*N),data2conv5 =>d49_in(5*N-1 downto 4*N),data2conv6 =>d49_in(4*N-1 downto 3*N),data2conv7 =>d49_in(3*N-1 downto 2*N),data2conv8 =>d49_in(2*N-1 downto N),data2conv9 =>d49_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d49_in(9*N-1 downto 8*N),w2 => d49_in(8*N-1 downto 7*N),w3 => d49_in(7*N-1 downto 6*N),w4 => d49_in(6*N-1 downto 5*N),w5 => d49_in(5*N-1 downto 4*N),w6 => d49_in(4*N-1 downto 3*N),w7 => d49_in(3*N-1 downto 2*N),w8 => d49_in(2*N-1 downto N),w9 => d49_in(N-1 downto 0 ),d_out => d49_out,en_out =>open  ,sof_out=>open   );
CL50: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d50_in(9*N-1 downto 8*N),data2conv2 =>d50_in(8*N-1 downto 7*N),data2conv3 =>d50_in(7*N-1 downto 6*N),data2conv4 =>d50_in(6*N-1 downto 5*N),data2conv5 =>d50_in(5*N-1 downto 4*N),data2conv6 =>d50_in(4*N-1 downto 3*N),data2conv7 =>d50_in(3*N-1 downto 2*N),data2conv8 =>d50_in(2*N-1 downto N),data2conv9 =>d50_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d50_in(9*N-1 downto 8*N),w2 => d50_in(8*N-1 downto 7*N),w3 => d50_in(7*N-1 downto 6*N),w4 => d50_in(6*N-1 downto 5*N),w5 => d50_in(5*N-1 downto 4*N),w6 => d50_in(4*N-1 downto 3*N),w7 => d50_in(3*N-1 downto 2*N),w8 => d50_in(2*N-1 downto N),w9 => d50_in(N-1 downto 0 ),d_out => d50_out,en_out =>open  ,sof_out=>open   );
CL51: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d51_in(9*N-1 downto 8*N),data2conv2 =>d51_in(8*N-1 downto 7*N),data2conv3 =>d51_in(7*N-1 downto 6*N),data2conv4 =>d51_in(6*N-1 downto 5*N),data2conv5 =>d51_in(5*N-1 downto 4*N),data2conv6 =>d51_in(4*N-1 downto 3*N),data2conv7 =>d51_in(3*N-1 downto 2*N),data2conv8 =>d51_in(2*N-1 downto N),data2conv9 =>d51_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d51_in(9*N-1 downto 8*N),w2 => d51_in(8*N-1 downto 7*N),w3 => d51_in(7*N-1 downto 6*N),w4 => d51_in(6*N-1 downto 5*N),w5 => d51_in(5*N-1 downto 4*N),w6 => d51_in(4*N-1 downto 3*N),w7 => d51_in(3*N-1 downto 2*N),w8 => d51_in(2*N-1 downto N),w9 => d51_in(N-1 downto 0 ),d_out => d51_out,en_out =>open  ,sof_out=>open   );
CL52: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d52_in(9*N-1 downto 8*N),data2conv2 =>d52_in(8*N-1 downto 7*N),data2conv3 =>d52_in(7*N-1 downto 6*N),data2conv4 =>d52_in(6*N-1 downto 5*N),data2conv5 =>d52_in(5*N-1 downto 4*N),data2conv6 =>d52_in(4*N-1 downto 3*N),data2conv7 =>d52_in(3*N-1 downto 2*N),data2conv8 =>d52_in(2*N-1 downto N),data2conv9 =>d52_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d52_in(9*N-1 downto 8*N),w2 => d52_in(8*N-1 downto 7*N),w3 => d52_in(7*N-1 downto 6*N),w4 => d52_in(6*N-1 downto 5*N),w5 => d52_in(5*N-1 downto 4*N),w6 => d52_in(4*N-1 downto 3*N),w7 => d52_in(3*N-1 downto 2*N),w8 => d52_in(2*N-1 downto N),w9 => d52_in(N-1 downto 0 ),d_out => d52_out,en_out =>open  ,sof_out=>open   );
CL53: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d53_in(9*N-1 downto 8*N),data2conv2 =>d53_in(8*N-1 downto 7*N),data2conv3 =>d53_in(7*N-1 downto 6*N),data2conv4 =>d53_in(6*N-1 downto 5*N),data2conv5 =>d53_in(5*N-1 downto 4*N),data2conv6 =>d53_in(4*N-1 downto 3*N),data2conv7 =>d53_in(3*N-1 downto 2*N),data2conv8 =>d53_in(2*N-1 downto N),data2conv9 =>d53_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d53_in(9*N-1 downto 8*N),w2 => d53_in(8*N-1 downto 7*N),w3 => d53_in(7*N-1 downto 6*N),w4 => d53_in(6*N-1 downto 5*N),w5 => d53_in(5*N-1 downto 4*N),w6 => d53_in(4*N-1 downto 3*N),w7 => d53_in(3*N-1 downto 2*N),w8 => d53_in(2*N-1 downto N),w9 => d53_in(N-1 downto 0 ),d_out => d53_out,en_out =>open  ,sof_out=>open   );
CL54: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d54_in(9*N-1 downto 8*N),data2conv2 =>d54_in(8*N-1 downto 7*N),data2conv3 =>d54_in(7*N-1 downto 6*N),data2conv4 =>d54_in(6*N-1 downto 5*N),data2conv5 =>d54_in(5*N-1 downto 4*N),data2conv6 =>d54_in(4*N-1 downto 3*N),data2conv7 =>d54_in(3*N-1 downto 2*N),data2conv8 =>d54_in(2*N-1 downto N),data2conv9 =>d54_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d54_in(9*N-1 downto 8*N),w2 => d54_in(8*N-1 downto 7*N),w3 => d54_in(7*N-1 downto 6*N),w4 => d54_in(6*N-1 downto 5*N),w5 => d54_in(5*N-1 downto 4*N),w6 => d54_in(4*N-1 downto 3*N),w7 => d54_in(3*N-1 downto 2*N),w8 => d54_in(2*N-1 downto N),w9 => d54_in(N-1 downto 0 ),d_out => d54_out,en_out =>open  ,sof_out=>open   );
CL55: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d55_in(9*N-1 downto 8*N),data2conv2 =>d55_in(8*N-1 downto 7*N),data2conv3 =>d55_in(7*N-1 downto 6*N),data2conv4 =>d55_in(6*N-1 downto 5*N),data2conv5 =>d55_in(5*N-1 downto 4*N),data2conv6 =>d55_in(4*N-1 downto 3*N),data2conv7 =>d55_in(3*N-1 downto 2*N),data2conv8 =>d55_in(2*N-1 downto N),data2conv9 =>d55_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d55_in(9*N-1 downto 8*N),w2 => d55_in(8*N-1 downto 7*N),w3 => d55_in(7*N-1 downto 6*N),w4 => d55_in(6*N-1 downto 5*N),w5 => d55_in(5*N-1 downto 4*N),w6 => d55_in(4*N-1 downto 3*N),w7 => d55_in(3*N-1 downto 2*N),w8 => d55_in(2*N-1 downto N),w9 => d55_in(N-1 downto 0 ),d_out => d55_out,en_out =>open  ,sof_out=>open   );
CL56: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d56_in(9*N-1 downto 8*N),data2conv2 =>d56_in(8*N-1 downto 7*N),data2conv3 =>d56_in(7*N-1 downto 6*N),data2conv4 =>d56_in(6*N-1 downto 5*N),data2conv5 =>d56_in(5*N-1 downto 4*N),data2conv6 =>d56_in(4*N-1 downto 3*N),data2conv7 =>d56_in(3*N-1 downto 2*N),data2conv8 =>d56_in(2*N-1 downto N),data2conv9 =>d56_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d56_in(9*N-1 downto 8*N),w2 => d56_in(8*N-1 downto 7*N),w3 => d56_in(7*N-1 downto 6*N),w4 => d56_in(6*N-1 downto 5*N),w5 => d56_in(5*N-1 downto 4*N),w6 => d56_in(4*N-1 downto 3*N),w7 => d56_in(3*N-1 downto 2*N),w8 => d56_in(2*N-1 downto N),w9 => d56_in(N-1 downto 0 ),d_out => d56_out,en_out =>open  ,sof_out=>open   );
CL57: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d57_in(9*N-1 downto 8*N),data2conv2 =>d57_in(8*N-1 downto 7*N),data2conv3 =>d57_in(7*N-1 downto 6*N),data2conv4 =>d57_in(6*N-1 downto 5*N),data2conv5 =>d57_in(5*N-1 downto 4*N),data2conv6 =>d57_in(4*N-1 downto 3*N),data2conv7 =>d57_in(3*N-1 downto 2*N),data2conv8 =>d57_in(2*N-1 downto N),data2conv9 =>d57_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d57_in(9*N-1 downto 8*N),w2 => d57_in(8*N-1 downto 7*N),w3 => d57_in(7*N-1 downto 6*N),w4 => d57_in(6*N-1 downto 5*N),w5 => d57_in(5*N-1 downto 4*N),w6 => d57_in(4*N-1 downto 3*N),w7 => d57_in(3*N-1 downto 2*N),w8 => d57_in(2*N-1 downto N),w9 => d57_in(N-1 downto 0 ),d_out => d57_out,en_out =>open  ,sof_out=>open   );
CL58: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d58_in(9*N-1 downto 8*N),data2conv2 =>d58_in(8*N-1 downto 7*N),data2conv3 =>d58_in(7*N-1 downto 6*N),data2conv4 =>d58_in(6*N-1 downto 5*N),data2conv5 =>d58_in(5*N-1 downto 4*N),data2conv6 =>d58_in(4*N-1 downto 3*N),data2conv7 =>d58_in(3*N-1 downto 2*N),data2conv8 =>d58_in(2*N-1 downto N),data2conv9 =>d58_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d58_in(9*N-1 downto 8*N),w2 => d58_in(8*N-1 downto 7*N),w3 => d58_in(7*N-1 downto 6*N),w4 => d58_in(6*N-1 downto 5*N),w5 => d58_in(5*N-1 downto 4*N),w6 => d58_in(4*N-1 downto 3*N),w7 => d58_in(3*N-1 downto 2*N),w8 => d58_in(2*N-1 downto N),w9 => d58_in(N-1 downto 0 ),d_out => d58_out,en_out =>open  ,sof_out=>open   );
CL59: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d59_in(9*N-1 downto 8*N),data2conv2 =>d59_in(8*N-1 downto 7*N),data2conv3 =>d59_in(7*N-1 downto 6*N),data2conv4 =>d59_in(6*N-1 downto 5*N),data2conv5 =>d59_in(5*N-1 downto 4*N),data2conv6 =>d59_in(4*N-1 downto 3*N),data2conv7 =>d59_in(3*N-1 downto 2*N),data2conv8 =>d59_in(2*N-1 downto N),data2conv9 =>d59_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d59_in(9*N-1 downto 8*N),w2 => d59_in(8*N-1 downto 7*N),w3 => d59_in(7*N-1 downto 6*N),w4 => d59_in(6*N-1 downto 5*N),w5 => d59_in(5*N-1 downto 4*N),w6 => d59_in(4*N-1 downto 3*N),w7 => d59_in(3*N-1 downto 2*N),w8 => d59_in(2*N-1 downto N),w9 => d59_in(N-1 downto 0 ),d_out => d59_out,en_out =>open  ,sof_out=>open   );
CL60: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d60_in(9*N-1 downto 8*N),data2conv2 =>d60_in(8*N-1 downto 7*N),data2conv3 =>d60_in(7*N-1 downto 6*N),data2conv4 =>d60_in(6*N-1 downto 5*N),data2conv5 =>d60_in(5*N-1 downto 4*N),data2conv6 =>d60_in(4*N-1 downto 3*N),data2conv7 =>d60_in(3*N-1 downto 2*N),data2conv8 =>d60_in(2*N-1 downto N),data2conv9 =>d60_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d60_in(9*N-1 downto 8*N),w2 => d60_in(8*N-1 downto 7*N),w3 => d60_in(7*N-1 downto 6*N),w4 => d60_in(6*N-1 downto 5*N),w5 => d60_in(5*N-1 downto 4*N),w6 => d60_in(4*N-1 downto 3*N),w7 => d60_in(3*N-1 downto 2*N),w8 => d60_in(2*N-1 downto N),w9 => d60_in(N-1 downto 0 ),d_out => d60_out,en_out =>open  ,sof_out=>open   );
CL61: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d61_in(9*N-1 downto 8*N),data2conv2 =>d61_in(8*N-1 downto 7*N),data2conv3 =>d61_in(7*N-1 downto 6*N),data2conv4 =>d61_in(6*N-1 downto 5*N),data2conv5 =>d61_in(5*N-1 downto 4*N),data2conv6 =>d61_in(4*N-1 downto 3*N),data2conv7 =>d61_in(3*N-1 downto 2*N),data2conv8 =>d61_in(2*N-1 downto N),data2conv9 =>d61_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d61_in(9*N-1 downto 8*N),w2 => d61_in(8*N-1 downto 7*N),w3 => d61_in(7*N-1 downto 6*N),w4 => d61_in(6*N-1 downto 5*N),w5 => d61_in(5*N-1 downto 4*N),w6 => d61_in(4*N-1 downto 3*N),w7 => d61_in(3*N-1 downto 2*N),w8 => d61_in(2*N-1 downto N),w9 => d61_in(N-1 downto 0 ),d_out => d61_out,en_out =>open  ,sof_out=>open   );
CL62: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d62_in(9*N-1 downto 8*N),data2conv2 =>d62_in(8*N-1 downto 7*N),data2conv3 =>d62_in(7*N-1 downto 6*N),data2conv4 =>d62_in(6*N-1 downto 5*N),data2conv5 =>d62_in(5*N-1 downto 4*N),data2conv6 =>d62_in(4*N-1 downto 3*N),data2conv7 =>d62_in(3*N-1 downto 2*N),data2conv8 =>d62_in(2*N-1 downto N),data2conv9 =>d62_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d62_in(9*N-1 downto 8*N),w2 => d62_in(8*N-1 downto 7*N),w3 => d62_in(7*N-1 downto 6*N),w4 => d62_in(6*N-1 downto 5*N),w5 => d62_in(5*N-1 downto 4*N),w6 => d62_in(4*N-1 downto 3*N),w7 => d62_in(3*N-1 downto 2*N),w8 => d62_in(2*N-1 downto N),w9 => d62_in(N-1 downto 0 ),d_out => d62_out,en_out =>open  ,sof_out=>open   );
CL63: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d63_in(9*N-1 downto 8*N),data2conv2 =>d63_in(8*N-1 downto 7*N),data2conv3 =>d63_in(7*N-1 downto 6*N),data2conv4 =>d63_in(6*N-1 downto 5*N),data2conv5 =>d63_in(5*N-1 downto 4*N),data2conv6 =>d63_in(4*N-1 downto 3*N),data2conv7 =>d63_in(3*N-1 downto 2*N),data2conv8 =>d63_in(2*N-1 downto N),data2conv9 =>d63_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d63_in(9*N-1 downto 8*N),w2 => d63_in(8*N-1 downto 7*N),w3 => d63_in(7*N-1 downto 6*N),w4 => d63_in(6*N-1 downto 5*N),w5 => d63_in(5*N-1 downto 4*N),w6 => d63_in(4*N-1 downto 3*N),w7 => d63_in(3*N-1 downto 2*N),w8 => d63_in(2*N-1 downto N),w9 => d63_in(N-1 downto 0 ),d_out => d63_out,en_out =>open  ,sof_out=>open   );
CL64: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d64_in(9*N-1 downto 8*N),data2conv2 =>d64_in(8*N-1 downto 7*N),data2conv3 =>d64_in(7*N-1 downto 6*N),data2conv4 =>d64_in(6*N-1 downto 5*N),data2conv5 =>d64_in(5*N-1 downto 4*N),data2conv6 =>d64_in(4*N-1 downto 3*N),data2conv7 =>d64_in(3*N-1 downto 2*N),data2conv8 =>d64_in(2*N-1 downto N),data2conv9 =>d64_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d64_in(9*N-1 downto 8*N),w2 => d64_in(8*N-1 downto 7*N),w3 => d64_in(7*N-1 downto 6*N),w4 => d64_in(6*N-1 downto 5*N),w5 => d64_in(5*N-1 downto 4*N),w6 => d64_in(4*N-1 downto 3*N),w7 => d64_in(3*N-1 downto 2*N),w8 => d64_in(2*N-1 downto N),w9 => d64_in(N-1 downto 0 ),d_out => d64_out,en_out =>open  ,sof_out=>open   );

CL65 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d65_in (9*N-1 downto 8*N),data2conv2 =>d65_in (8*N-1 downto 7*N),data2conv3 =>d65_in (7*N-1 downto 6*N),data2conv4 =>d65_in (6*N-1 downto 5*N),data2conv5 =>d65_in (5*N-1 downto 4*N),data2conv6 =>d65_in (4*N-1 downto 3*N),data2conv7 =>d65_in (3*N-1 downto 2*N),data2conv8 =>d65_in (2*N-1 downto N),data2conv9 =>d65_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d65_in (9*N-1 downto 8*N),w2 => d65_in (8*N-1 downto 7*N),w3 => d65_in (7*N-1 downto 6*N),w4 => d65_in (6*N-1 downto 5*N),w5 => d65_in (5*N-1 downto 4*N),w6 => d65_in (4*N-1 downto 3*N),w7 => d65_in (3*N-1 downto 2*N),w8 => d65_in (2*N-1 downto N),w9 => d65_in (N-1 downto 0 ),d_out => d65_out ,en_out =>open  ,sof_out=>open   );
CL66 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d66_in (9*N-1 downto 8*N),data2conv2 =>d66_in (8*N-1 downto 7*N),data2conv3 =>d66_in (7*N-1 downto 6*N),data2conv4 =>d66_in (6*N-1 downto 5*N),data2conv5 =>d66_in (5*N-1 downto 4*N),data2conv6 =>d66_in (4*N-1 downto 3*N),data2conv7 =>d66_in (3*N-1 downto 2*N),data2conv8 =>d66_in (2*N-1 downto N),data2conv9 =>d66_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d66_in (9*N-1 downto 8*N),w2 => d66_in (8*N-1 downto 7*N),w3 => d66_in (7*N-1 downto 6*N),w4 => d66_in (6*N-1 downto 5*N),w5 => d66_in (5*N-1 downto 4*N),w6 => d66_in (4*N-1 downto 3*N),w7 => d66_in (3*N-1 downto 2*N),w8 => d66_in (2*N-1 downto N),w9 => d66_in (N-1 downto 0 ),d_out => d66_out ,en_out =>open  ,sof_out=>open   );
CL67 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d67_in (9*N-1 downto 8*N),data2conv2 =>d67_in (8*N-1 downto 7*N),data2conv3 =>d67_in (7*N-1 downto 6*N),data2conv4 =>d67_in (6*N-1 downto 5*N),data2conv5 =>d67_in (5*N-1 downto 4*N),data2conv6 =>d67_in (4*N-1 downto 3*N),data2conv7 =>d67_in (3*N-1 downto 2*N),data2conv8 =>d67_in (2*N-1 downto N),data2conv9 =>d67_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d67_in (9*N-1 downto 8*N),w2 => d67_in (8*N-1 downto 7*N),w3 => d67_in (7*N-1 downto 6*N),w4 => d67_in (6*N-1 downto 5*N),w5 => d67_in (5*N-1 downto 4*N),w6 => d67_in (4*N-1 downto 3*N),w7 => d67_in (3*N-1 downto 2*N),w8 => d67_in (2*N-1 downto N),w9 => d67_in (N-1 downto 0 ),d_out => d67_out ,en_out =>open  ,sof_out=>open   );
CL68 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d68_in (9*N-1 downto 8*N),data2conv2 =>d68_in (8*N-1 downto 7*N),data2conv3 =>d68_in (7*N-1 downto 6*N),data2conv4 =>d68_in (6*N-1 downto 5*N),data2conv5 =>d68_in (5*N-1 downto 4*N),data2conv6 =>d68_in (4*N-1 downto 3*N),data2conv7 =>d68_in (3*N-1 downto 2*N),data2conv8 =>d68_in (2*N-1 downto N),data2conv9 =>d68_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d68_in (9*N-1 downto 8*N),w2 => d68_in (8*N-1 downto 7*N),w3 => d68_in (7*N-1 downto 6*N),w4 => d68_in (6*N-1 downto 5*N),w5 => d68_in (5*N-1 downto 4*N),w6 => d68_in (4*N-1 downto 3*N),w7 => d68_in (3*N-1 downto 2*N),w8 => d68_in (2*N-1 downto N),w9 => d68_in (N-1 downto 0 ),d_out => d68_out ,en_out =>open  ,sof_out=>open   );
CL69 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d69_in (9*N-1 downto 8*N),data2conv2 =>d69_in (8*N-1 downto 7*N),data2conv3 =>d69_in (7*N-1 downto 6*N),data2conv4 =>d69_in (6*N-1 downto 5*N),data2conv5 =>d69_in (5*N-1 downto 4*N),data2conv6 =>d69_in (4*N-1 downto 3*N),data2conv7 =>d69_in (3*N-1 downto 2*N),data2conv8 =>d69_in (2*N-1 downto N),data2conv9 =>d69_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d69_in (9*N-1 downto 8*N),w2 => d69_in (8*N-1 downto 7*N),w3 => d69_in (7*N-1 downto 6*N),w4 => d69_in (6*N-1 downto 5*N),w5 => d69_in (5*N-1 downto 4*N),w6 => d69_in (4*N-1 downto 3*N),w7 => d69_in (3*N-1 downto 2*N),w8 => d69_in (2*N-1 downto N),w9 => d69_in (N-1 downto 0 ),d_out => d69_out ,en_out =>open  ,sof_out=>open   );
CL70 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d70_in (9*N-1 downto 8*N),data2conv2 =>d70_in (8*N-1 downto 7*N),data2conv3 =>d70_in (7*N-1 downto 6*N),data2conv4 =>d70_in (6*N-1 downto 5*N),data2conv5 =>d70_in (5*N-1 downto 4*N),data2conv6 =>d70_in (4*N-1 downto 3*N),data2conv7 =>d70_in (3*N-1 downto 2*N),data2conv8 =>d70_in (2*N-1 downto N),data2conv9 =>d70_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d70_in (9*N-1 downto 8*N),w2 => d70_in (8*N-1 downto 7*N),w3 => d70_in (7*N-1 downto 6*N),w4 => d70_in (6*N-1 downto 5*N),w5 => d70_in (5*N-1 downto 4*N),w6 => d70_in (4*N-1 downto 3*N),w7 => d70_in (3*N-1 downto 2*N),w8 => d70_in (2*N-1 downto N),w9 => d70_in (N-1 downto 0 ),d_out => d70_out ,en_out =>open  ,sof_out=>open   );
CL71 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d71_in (9*N-1 downto 8*N),data2conv2 =>d71_in (8*N-1 downto 7*N),data2conv3 =>d71_in (7*N-1 downto 6*N),data2conv4 =>d71_in (6*N-1 downto 5*N),data2conv5 =>d71_in (5*N-1 downto 4*N),data2conv6 =>d71_in (4*N-1 downto 3*N),data2conv7 =>d71_in (3*N-1 downto 2*N),data2conv8 =>d71_in (2*N-1 downto N),data2conv9 =>d71_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d71_in (9*N-1 downto 8*N),w2 => d71_in (8*N-1 downto 7*N),w3 => d71_in (7*N-1 downto 6*N),w4 => d71_in (6*N-1 downto 5*N),w5 => d71_in (5*N-1 downto 4*N),w6 => d71_in (4*N-1 downto 3*N),w7 => d71_in (3*N-1 downto 2*N),w8 => d71_in (2*N-1 downto N),w9 => d71_in (N-1 downto 0 ),d_out => d71_out ,en_out =>open  ,sof_out=>open   );
CL72 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d72_in (9*N-1 downto 8*N),data2conv2 =>d72_in (8*N-1 downto 7*N),data2conv3 =>d72_in (7*N-1 downto 6*N),data2conv4 =>d72_in (6*N-1 downto 5*N),data2conv5 =>d72_in (5*N-1 downto 4*N),data2conv6 =>d72_in (4*N-1 downto 3*N),data2conv7 =>d72_in (3*N-1 downto 2*N),data2conv8 =>d72_in (2*N-1 downto N),data2conv9 =>d72_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d72_in (9*N-1 downto 8*N),w2 => d72_in (8*N-1 downto 7*N),w3 => d72_in (7*N-1 downto 6*N),w4 => d72_in (6*N-1 downto 5*N),w5 => d72_in (5*N-1 downto 4*N),w6 => d72_in (4*N-1 downto 3*N),w7 => d72_in (3*N-1 downto 2*N),w8 => d72_in (2*N-1 downto N),w9 => d72_in (N-1 downto 0 ),d_out => d72_out ,en_out =>open  ,sof_out=>open   );
CL73 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d73_in (9*N-1 downto 8*N),data2conv2 =>d73_in (8*N-1 downto 7*N),data2conv3 =>d73_in (7*N-1 downto 6*N),data2conv4 =>d73_in (6*N-1 downto 5*N),data2conv5 =>d73_in (5*N-1 downto 4*N),data2conv6 =>d73_in (4*N-1 downto 3*N),data2conv7 =>d73_in (3*N-1 downto 2*N),data2conv8 =>d73_in (2*N-1 downto N),data2conv9 =>d73_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d73_in (9*N-1 downto 8*N),w2 => d73_in (8*N-1 downto 7*N),w3 => d73_in (7*N-1 downto 6*N),w4 => d73_in (6*N-1 downto 5*N),w5 => d73_in (5*N-1 downto 4*N),w6 => d73_in (4*N-1 downto 3*N),w7 => d73_in (3*N-1 downto 2*N),w8 => d73_in (2*N-1 downto N),w9 => d73_in (N-1 downto 0 ),d_out => d73_out ,en_out =>open  ,sof_out=>open   );
CL74 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d74_in (9*N-1 downto 8*N),data2conv2 =>d74_in (8*N-1 downto 7*N),data2conv3 =>d74_in (7*N-1 downto 6*N),data2conv4 =>d74_in (6*N-1 downto 5*N),data2conv5 =>d74_in (5*N-1 downto 4*N),data2conv6 =>d74_in (4*N-1 downto 3*N),data2conv7 =>d74_in (3*N-1 downto 2*N),data2conv8 =>d74_in (2*N-1 downto N),data2conv9 =>d74_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d74_in (9*N-1 downto 8*N),w2 => d74_in (8*N-1 downto 7*N),w3 => d74_in (7*N-1 downto 6*N),w4 => d74_in (6*N-1 downto 5*N),w5 => d74_in (5*N-1 downto 4*N),w6 => d74_in (4*N-1 downto 3*N),w7 => d74_in (3*N-1 downto 2*N),w8 => d74_in (2*N-1 downto N),w9 => d74_in (N-1 downto 0 ),d_out => d74_out ,en_out =>open  ,sof_out=>open   );
CL75 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d75_in (9*N-1 downto 8*N),data2conv2 =>d75_in (8*N-1 downto 7*N),data2conv3 =>d75_in (7*N-1 downto 6*N),data2conv4 =>d75_in (6*N-1 downto 5*N),data2conv5 =>d75_in (5*N-1 downto 4*N),data2conv6 =>d75_in (4*N-1 downto 3*N),data2conv7 =>d75_in (3*N-1 downto 2*N),data2conv8 =>d75_in (2*N-1 downto N),data2conv9 =>d75_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d75_in (9*N-1 downto 8*N),w2 => d75_in (8*N-1 downto 7*N),w3 => d75_in (7*N-1 downto 6*N),w4 => d75_in (6*N-1 downto 5*N),w5 => d75_in (5*N-1 downto 4*N),w6 => d75_in (4*N-1 downto 3*N),w7 => d75_in (3*N-1 downto 2*N),w8 => d75_in (2*N-1 downto N),w9 => d75_in (N-1 downto 0 ),d_out => d75_out ,en_out =>open  ,sof_out=>open   );
CL76 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d76_in (9*N-1 downto 8*N),data2conv2 =>d76_in (8*N-1 downto 7*N),data2conv3 =>d76_in (7*N-1 downto 6*N),data2conv4 =>d76_in (6*N-1 downto 5*N),data2conv5 =>d76_in (5*N-1 downto 4*N),data2conv6 =>d76_in (4*N-1 downto 3*N),data2conv7 =>d76_in (3*N-1 downto 2*N),data2conv8 =>d76_in (2*N-1 downto N),data2conv9 =>d76_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d76_in (9*N-1 downto 8*N),w2 => d76_in (8*N-1 downto 7*N),w3 => d76_in (7*N-1 downto 6*N),w4 => d76_in (6*N-1 downto 5*N),w5 => d76_in (5*N-1 downto 4*N),w6 => d76_in (4*N-1 downto 3*N),w7 => d76_in (3*N-1 downto 2*N),w8 => d76_in (2*N-1 downto N),w9 => d76_in (N-1 downto 0 ),d_out => d76_out ,en_out =>open  ,sof_out=>open   );
CL77 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d77_in (9*N-1 downto 8*N),data2conv2 =>d77_in (8*N-1 downto 7*N),data2conv3 =>d77_in (7*N-1 downto 6*N),data2conv4 =>d77_in (6*N-1 downto 5*N),data2conv5 =>d77_in (5*N-1 downto 4*N),data2conv6 =>d77_in (4*N-1 downto 3*N),data2conv7 =>d77_in (3*N-1 downto 2*N),data2conv8 =>d77_in (2*N-1 downto N),data2conv9 =>d77_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d77_in (9*N-1 downto 8*N),w2 => d77_in (8*N-1 downto 7*N),w3 => d77_in (7*N-1 downto 6*N),w4 => d77_in (6*N-1 downto 5*N),w5 => d77_in (5*N-1 downto 4*N),w6 => d77_in (4*N-1 downto 3*N),w7 => d77_in (3*N-1 downto 2*N),w8 => d77_in (2*N-1 downto N),w9 => d77_in (N-1 downto 0 ),d_out => d77_out ,en_out =>open  ,sof_out=>open   );
CL78 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d78_in (9*N-1 downto 8*N),data2conv2 =>d78_in (8*N-1 downto 7*N),data2conv3 =>d78_in (7*N-1 downto 6*N),data2conv4 =>d78_in (6*N-1 downto 5*N),data2conv5 =>d78_in (5*N-1 downto 4*N),data2conv6 =>d78_in (4*N-1 downto 3*N),data2conv7 =>d78_in (3*N-1 downto 2*N),data2conv8 =>d78_in (2*N-1 downto N),data2conv9 =>d78_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d78_in (9*N-1 downto 8*N),w2 => d78_in (8*N-1 downto 7*N),w3 => d78_in (7*N-1 downto 6*N),w4 => d78_in (6*N-1 downto 5*N),w5 => d78_in (5*N-1 downto 4*N),w6 => d78_in (4*N-1 downto 3*N),w7 => d78_in (3*N-1 downto 2*N),w8 => d78_in (2*N-1 downto N),w9 => d78_in (N-1 downto 0 ),d_out => d78_out ,en_out =>open  ,sof_out=>open   );
CL79 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d79_in (9*N-1 downto 8*N),data2conv2 =>d79_in (8*N-1 downto 7*N),data2conv3 =>d79_in (7*N-1 downto 6*N),data2conv4 =>d79_in (6*N-1 downto 5*N),data2conv5 =>d79_in (5*N-1 downto 4*N),data2conv6 =>d79_in (4*N-1 downto 3*N),data2conv7 =>d79_in (3*N-1 downto 2*N),data2conv8 =>d79_in (2*N-1 downto N),data2conv9 =>d79_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d79_in (9*N-1 downto 8*N),w2 => d79_in (8*N-1 downto 7*N),w3 => d79_in (7*N-1 downto 6*N),w4 => d79_in (6*N-1 downto 5*N),w5 => d79_in (5*N-1 downto 4*N),w6 => d79_in (4*N-1 downto 3*N),w7 => d79_in (3*N-1 downto 2*N),w8 => d79_in (2*N-1 downto N),w9 => d79_in (N-1 downto 0 ),d_out => d79_out ,en_out =>open  ,sof_out=>open   );
CL80 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d80_in (9*N-1 downto 8*N),data2conv2 =>d80_in (8*N-1 downto 7*N),data2conv3 =>d80_in (7*N-1 downto 6*N),data2conv4 =>d80_in (6*N-1 downto 5*N),data2conv5 =>d80_in (5*N-1 downto 4*N),data2conv6 =>d80_in (4*N-1 downto 3*N),data2conv7 =>d80_in (3*N-1 downto 2*N),data2conv8 =>d80_in (2*N-1 downto N),data2conv9 =>d80_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d80_in (9*N-1 downto 8*N),w2 => d80_in (8*N-1 downto 7*N),w3 => d80_in (7*N-1 downto 6*N),w4 => d80_in (6*N-1 downto 5*N),w5 => d80_in (5*N-1 downto 4*N),w6 => d80_in (4*N-1 downto 3*N),w7 => d80_in (3*N-1 downto 2*N),w8 => d80_in (2*N-1 downto N),w9 => d80_in (N-1 downto 0 ),d_out => d80_out ,en_out =>open  ,sof_out=>open   );
CL81 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d81_in (9*N-1 downto 8*N),data2conv2 =>d81_in (8*N-1 downto 7*N),data2conv3 =>d81_in (7*N-1 downto 6*N),data2conv4 =>d81_in (6*N-1 downto 5*N),data2conv5 =>d81_in (5*N-1 downto 4*N),data2conv6 =>d81_in (4*N-1 downto 3*N),data2conv7 =>d81_in (3*N-1 downto 2*N),data2conv8 =>d81_in (2*N-1 downto N),data2conv9 =>d81_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d81_in (9*N-1 downto 8*N),w2 => d81_in (8*N-1 downto 7*N),w3 => d81_in (7*N-1 downto 6*N),w4 => d81_in (6*N-1 downto 5*N),w5 => d81_in (5*N-1 downto 4*N),w6 => d81_in (4*N-1 downto 3*N),w7 => d81_in (3*N-1 downto 2*N),w8 => d81_in (2*N-1 downto N),w9 => d81_in (N-1 downto 0 ),d_out => d81_out ,en_out =>open  ,sof_out=>open   );
CL82 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d82_in (9*N-1 downto 8*N),data2conv2 =>d82_in (8*N-1 downto 7*N),data2conv3 =>d82_in (7*N-1 downto 6*N),data2conv4 =>d82_in (6*N-1 downto 5*N),data2conv5 =>d82_in (5*N-1 downto 4*N),data2conv6 =>d82_in (4*N-1 downto 3*N),data2conv7 =>d82_in (3*N-1 downto 2*N),data2conv8 =>d82_in (2*N-1 downto N),data2conv9 =>d82_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d82_in (9*N-1 downto 8*N),w2 => d82_in (8*N-1 downto 7*N),w3 => d82_in (7*N-1 downto 6*N),w4 => d82_in (6*N-1 downto 5*N),w5 => d82_in (5*N-1 downto 4*N),w6 => d82_in (4*N-1 downto 3*N),w7 => d82_in (3*N-1 downto 2*N),w8 => d82_in (2*N-1 downto N),w9 => d82_in (N-1 downto 0 ),d_out => d82_out ,en_out =>open  ,sof_out=>open   );
CL83 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d83_in (9*N-1 downto 8*N),data2conv2 =>d83_in (8*N-1 downto 7*N),data2conv3 =>d83_in (7*N-1 downto 6*N),data2conv4 =>d83_in (6*N-1 downto 5*N),data2conv5 =>d83_in (5*N-1 downto 4*N),data2conv6 =>d83_in (4*N-1 downto 3*N),data2conv7 =>d83_in (3*N-1 downto 2*N),data2conv8 =>d83_in (2*N-1 downto N),data2conv9 =>d83_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d83_in (9*N-1 downto 8*N),w2 => d83_in (8*N-1 downto 7*N),w3 => d83_in (7*N-1 downto 6*N),w4 => d83_in (6*N-1 downto 5*N),w5 => d83_in (5*N-1 downto 4*N),w6 => d83_in (4*N-1 downto 3*N),w7 => d83_in (3*N-1 downto 2*N),w8 => d83_in (2*N-1 downto N),w9 => d83_in (N-1 downto 0 ),d_out => d83_out ,en_out =>open  ,sof_out=>open   );
CL84 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d84_in (9*N-1 downto 8*N),data2conv2 =>d84_in (8*N-1 downto 7*N),data2conv3 =>d84_in (7*N-1 downto 6*N),data2conv4 =>d84_in (6*N-1 downto 5*N),data2conv5 =>d84_in (5*N-1 downto 4*N),data2conv6 =>d84_in (4*N-1 downto 3*N),data2conv7 =>d84_in (3*N-1 downto 2*N),data2conv8 =>d84_in (2*N-1 downto N),data2conv9 =>d84_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d84_in (9*N-1 downto 8*N),w2 => d84_in (8*N-1 downto 7*N),w3 => d84_in (7*N-1 downto 6*N),w4 => d84_in (6*N-1 downto 5*N),w5 => d84_in (5*N-1 downto 4*N),w6 => d84_in (4*N-1 downto 3*N),w7 => d84_in (3*N-1 downto 2*N),w8 => d84_in (2*N-1 downto N),w9 => d84_in (N-1 downto 0 ),d_out => d84_out ,en_out =>open  ,sof_out=>open   );
CL85 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d85_in (9*N-1 downto 8*N),data2conv2 =>d85_in (8*N-1 downto 7*N),data2conv3 =>d85_in (7*N-1 downto 6*N),data2conv4 =>d85_in (6*N-1 downto 5*N),data2conv5 =>d85_in (5*N-1 downto 4*N),data2conv6 =>d85_in (4*N-1 downto 3*N),data2conv7 =>d85_in (3*N-1 downto 2*N),data2conv8 =>d85_in (2*N-1 downto N),data2conv9 =>d85_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d85_in (9*N-1 downto 8*N),w2 => d85_in (8*N-1 downto 7*N),w3 => d85_in (7*N-1 downto 6*N),w4 => d85_in (6*N-1 downto 5*N),w5 => d85_in (5*N-1 downto 4*N),w6 => d85_in (4*N-1 downto 3*N),w7 => d85_in (3*N-1 downto 2*N),w8 => d85_in (2*N-1 downto N),w9 => d85_in (N-1 downto 0 ),d_out => d85_out ,en_out =>open  ,sof_out=>open   );
CL86 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d86_in (9*N-1 downto 8*N),data2conv2 =>d86_in (8*N-1 downto 7*N),data2conv3 =>d86_in (7*N-1 downto 6*N),data2conv4 =>d86_in (6*N-1 downto 5*N),data2conv5 =>d86_in (5*N-1 downto 4*N),data2conv6 =>d86_in (4*N-1 downto 3*N),data2conv7 =>d86_in (3*N-1 downto 2*N),data2conv8 =>d86_in (2*N-1 downto N),data2conv9 =>d86_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d86_in (9*N-1 downto 8*N),w2 => d86_in (8*N-1 downto 7*N),w3 => d86_in (7*N-1 downto 6*N),w4 => d86_in (6*N-1 downto 5*N),w5 => d86_in (5*N-1 downto 4*N),w6 => d86_in (4*N-1 downto 3*N),w7 => d86_in (3*N-1 downto 2*N),w8 => d86_in (2*N-1 downto N),w9 => d86_in (N-1 downto 0 ),d_out => d86_out ,en_out =>open  ,sof_out=>open   );
CL87 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d87_in (9*N-1 downto 8*N),data2conv2 =>d87_in (8*N-1 downto 7*N),data2conv3 =>d87_in (7*N-1 downto 6*N),data2conv4 =>d87_in (6*N-1 downto 5*N),data2conv5 =>d87_in (5*N-1 downto 4*N),data2conv6 =>d87_in (4*N-1 downto 3*N),data2conv7 =>d87_in (3*N-1 downto 2*N),data2conv8 =>d87_in (2*N-1 downto N),data2conv9 =>d87_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d87_in (9*N-1 downto 8*N),w2 => d87_in (8*N-1 downto 7*N),w3 => d87_in (7*N-1 downto 6*N),w4 => d87_in (6*N-1 downto 5*N),w5 => d87_in (5*N-1 downto 4*N),w6 => d87_in (4*N-1 downto 3*N),w7 => d87_in (3*N-1 downto 2*N),w8 => d87_in (2*N-1 downto N),w9 => d87_in (N-1 downto 0 ),d_out => d87_out ,en_out =>open  ,sof_out=>open   );
CL88 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d88_in (9*N-1 downto 8*N),data2conv2 =>d88_in (8*N-1 downto 7*N),data2conv3 =>d88_in (7*N-1 downto 6*N),data2conv4 =>d88_in (6*N-1 downto 5*N),data2conv5 =>d88_in (5*N-1 downto 4*N),data2conv6 =>d88_in (4*N-1 downto 3*N),data2conv7 =>d88_in (3*N-1 downto 2*N),data2conv8 =>d88_in (2*N-1 downto N),data2conv9 =>d88_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d88_in (9*N-1 downto 8*N),w2 => d88_in (8*N-1 downto 7*N),w3 => d88_in (7*N-1 downto 6*N),w4 => d88_in (6*N-1 downto 5*N),w5 => d88_in (5*N-1 downto 4*N),w6 => d88_in (4*N-1 downto 3*N),w7 => d88_in (3*N-1 downto 2*N),w8 => d88_in (2*N-1 downto N),w9 => d88_in (N-1 downto 0 ),d_out => d88_out ,en_out =>open  ,sof_out=>open   );
CL89 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d89_in (9*N-1 downto 8*N),data2conv2 =>d89_in (8*N-1 downto 7*N),data2conv3 =>d89_in (7*N-1 downto 6*N),data2conv4 =>d89_in (6*N-1 downto 5*N),data2conv5 =>d89_in (5*N-1 downto 4*N),data2conv6 =>d89_in (4*N-1 downto 3*N),data2conv7 =>d89_in (3*N-1 downto 2*N),data2conv8 =>d89_in (2*N-1 downto N),data2conv9 =>d89_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d89_in (9*N-1 downto 8*N),w2 => d89_in (8*N-1 downto 7*N),w3 => d89_in (7*N-1 downto 6*N),w4 => d89_in (6*N-1 downto 5*N),w5 => d89_in (5*N-1 downto 4*N),w6 => d89_in (4*N-1 downto 3*N),w7 => d89_in (3*N-1 downto 2*N),w8 => d89_in (2*N-1 downto N),w9 => d89_in (N-1 downto 0 ),d_out => d89_out ,en_out =>open  ,sof_out=>open   );
CL90 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d90_in (9*N-1 downto 8*N),data2conv2 =>d90_in (8*N-1 downto 7*N),data2conv3 =>d90_in (7*N-1 downto 6*N),data2conv4 =>d90_in (6*N-1 downto 5*N),data2conv5 =>d90_in (5*N-1 downto 4*N),data2conv6 =>d90_in (4*N-1 downto 3*N),data2conv7 =>d90_in (3*N-1 downto 2*N),data2conv8 =>d90_in (2*N-1 downto N),data2conv9 =>d90_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d90_in (9*N-1 downto 8*N),w2 => d90_in (8*N-1 downto 7*N),w3 => d90_in (7*N-1 downto 6*N),w4 => d90_in (6*N-1 downto 5*N),w5 => d90_in (5*N-1 downto 4*N),w6 => d90_in (4*N-1 downto 3*N),w7 => d90_in (3*N-1 downto 2*N),w8 => d90_in (2*N-1 downto N),w9 => d90_in (N-1 downto 0 ),d_out => d90_out ,en_out =>open  ,sof_out=>open   );
CL91 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d91_in (9*N-1 downto 8*N),data2conv2 =>d91_in (8*N-1 downto 7*N),data2conv3 =>d91_in (7*N-1 downto 6*N),data2conv4 =>d91_in (6*N-1 downto 5*N),data2conv5 =>d91_in (5*N-1 downto 4*N),data2conv6 =>d91_in (4*N-1 downto 3*N),data2conv7 =>d91_in (3*N-1 downto 2*N),data2conv8 =>d91_in (2*N-1 downto N),data2conv9 =>d91_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d91_in (9*N-1 downto 8*N),w2 => d91_in (8*N-1 downto 7*N),w3 => d91_in (7*N-1 downto 6*N),w4 => d91_in (6*N-1 downto 5*N),w5 => d91_in (5*N-1 downto 4*N),w6 => d91_in (4*N-1 downto 3*N),w7 => d91_in (3*N-1 downto 2*N),w8 => d91_in (2*N-1 downto N),w9 => d91_in (N-1 downto 0 ),d_out => d91_out ,en_out =>open  ,sof_out=>open   );
CL92 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d92_in (9*N-1 downto 8*N),data2conv2 =>d92_in (8*N-1 downto 7*N),data2conv3 =>d92_in (7*N-1 downto 6*N),data2conv4 =>d92_in (6*N-1 downto 5*N),data2conv5 =>d92_in (5*N-1 downto 4*N),data2conv6 =>d92_in (4*N-1 downto 3*N),data2conv7 =>d92_in (3*N-1 downto 2*N),data2conv8 =>d92_in (2*N-1 downto N),data2conv9 =>d92_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d92_in (9*N-1 downto 8*N),w2 => d92_in (8*N-1 downto 7*N),w3 => d92_in (7*N-1 downto 6*N),w4 => d92_in (6*N-1 downto 5*N),w5 => d92_in (5*N-1 downto 4*N),w6 => d92_in (4*N-1 downto 3*N),w7 => d92_in (3*N-1 downto 2*N),w8 => d92_in (2*N-1 downto N),w9 => d92_in (N-1 downto 0 ),d_out => d92_out ,en_out =>open  ,sof_out=>open   );
CL93 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d93_in (9*N-1 downto 8*N),data2conv2 =>d93_in (8*N-1 downto 7*N),data2conv3 =>d93_in (7*N-1 downto 6*N),data2conv4 =>d93_in (6*N-1 downto 5*N),data2conv5 =>d93_in (5*N-1 downto 4*N),data2conv6 =>d93_in (4*N-1 downto 3*N),data2conv7 =>d93_in (3*N-1 downto 2*N),data2conv8 =>d93_in (2*N-1 downto N),data2conv9 =>d93_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d93_in (9*N-1 downto 8*N),w2 => d93_in (8*N-1 downto 7*N),w3 => d93_in (7*N-1 downto 6*N),w4 => d93_in (6*N-1 downto 5*N),w5 => d93_in (5*N-1 downto 4*N),w6 => d93_in (4*N-1 downto 3*N),w7 => d93_in (3*N-1 downto 2*N),w8 => d93_in (2*N-1 downto N),w9 => d93_in (N-1 downto 0 ),d_out => d93_out ,en_out =>open  ,sof_out=>open   );
CL94 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d94_in (9*N-1 downto 8*N),data2conv2 =>d94_in (8*N-1 downto 7*N),data2conv3 =>d94_in (7*N-1 downto 6*N),data2conv4 =>d94_in (6*N-1 downto 5*N),data2conv5 =>d94_in (5*N-1 downto 4*N),data2conv6 =>d94_in (4*N-1 downto 3*N),data2conv7 =>d94_in (3*N-1 downto 2*N),data2conv8 =>d94_in (2*N-1 downto N),data2conv9 =>d94_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d94_in (9*N-1 downto 8*N),w2 => d94_in (8*N-1 downto 7*N),w3 => d94_in (7*N-1 downto 6*N),w4 => d94_in (6*N-1 downto 5*N),w5 => d94_in (5*N-1 downto 4*N),w6 => d94_in (4*N-1 downto 3*N),w7 => d94_in (3*N-1 downto 2*N),w8 => d94_in (2*N-1 downto N),w9 => d94_in (N-1 downto 0 ),d_out => d94_out ,en_out =>open  ,sof_out=>open   );
CL95 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d95_in (9*N-1 downto 8*N),data2conv2 =>d95_in (8*N-1 downto 7*N),data2conv3 =>d95_in (7*N-1 downto 6*N),data2conv4 =>d95_in (6*N-1 downto 5*N),data2conv5 =>d95_in (5*N-1 downto 4*N),data2conv6 =>d95_in (4*N-1 downto 3*N),data2conv7 =>d95_in (3*N-1 downto 2*N),data2conv8 =>d95_in (2*N-1 downto N),data2conv9 =>d95_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d95_in (9*N-1 downto 8*N),w2 => d95_in (8*N-1 downto 7*N),w3 => d95_in (7*N-1 downto 6*N),w4 => d95_in (6*N-1 downto 5*N),w5 => d95_in (5*N-1 downto 4*N),w6 => d95_in (4*N-1 downto 3*N),w7 => d95_in (3*N-1 downto 2*N),w8 => d95_in (2*N-1 downto N),w9 => d95_in (N-1 downto 0 ),d_out => d95_out ,en_out =>open  ,sof_out=>open   );
CL96 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d96_in (9*N-1 downto 8*N),data2conv2 =>d96_in (8*N-1 downto 7*N),data2conv3 =>d96_in (7*N-1 downto 6*N),data2conv4 =>d96_in (6*N-1 downto 5*N),data2conv5 =>d96_in (5*N-1 downto 4*N),data2conv6 =>d96_in (4*N-1 downto 3*N),data2conv7 =>d96_in (3*N-1 downto 2*N),data2conv8 =>d96_in (2*N-1 downto N),data2conv9 =>d96_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d96_in (9*N-1 downto 8*N),w2 => d96_in (8*N-1 downto 7*N),w3 => d96_in (7*N-1 downto 6*N),w4 => d96_in (6*N-1 downto 5*N),w5 => d96_in (5*N-1 downto 4*N),w6 => d96_in (4*N-1 downto 3*N),w7 => d96_in (3*N-1 downto 2*N),w8 => d96_in (2*N-1 downto N),w9 => d96_in (N-1 downto 0 ),d_out => d96_out ,en_out =>open  ,sof_out=>open   );
CL97 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d97_in (9*N-1 downto 8*N),data2conv2 =>d97_in (8*N-1 downto 7*N),data2conv3 =>d97_in (7*N-1 downto 6*N),data2conv4 =>d97_in (6*N-1 downto 5*N),data2conv5 =>d97_in (5*N-1 downto 4*N),data2conv6 =>d97_in (4*N-1 downto 3*N),data2conv7 =>d97_in (3*N-1 downto 2*N),data2conv8 =>d97_in (2*N-1 downto N),data2conv9 =>d97_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d97_in (9*N-1 downto 8*N),w2 => d97_in (8*N-1 downto 7*N),w3 => d97_in (7*N-1 downto 6*N),w4 => d97_in (6*N-1 downto 5*N),w5 => d97_in (5*N-1 downto 4*N),w6 => d97_in (4*N-1 downto 3*N),w7 => d97_in (3*N-1 downto 2*N),w8 => d97_in (2*N-1 downto N),w9 => d97_in (N-1 downto 0 ),d_out => d97_out ,en_out =>open  ,sof_out=>open   );
CL98 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d98_in (9*N-1 downto 8*N),data2conv2 =>d98_in (8*N-1 downto 7*N),data2conv3 =>d98_in (7*N-1 downto 6*N),data2conv4 =>d98_in (6*N-1 downto 5*N),data2conv5 =>d98_in (5*N-1 downto 4*N),data2conv6 =>d98_in (4*N-1 downto 3*N),data2conv7 =>d98_in (3*N-1 downto 2*N),data2conv8 =>d98_in (2*N-1 downto N),data2conv9 =>d98_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d98_in (9*N-1 downto 8*N),w2 => d98_in (8*N-1 downto 7*N),w3 => d98_in (7*N-1 downto 6*N),w4 => d98_in (6*N-1 downto 5*N),w5 => d98_in (5*N-1 downto 4*N),w6 => d98_in (4*N-1 downto 3*N),w7 => d98_in (3*N-1 downto 2*N),w8 => d98_in (2*N-1 downto N),w9 => d98_in (N-1 downto 0 ),d_out => d98_out ,en_out =>open  ,sof_out=>open   );
CL99 : ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d99_in (9*N-1 downto 8*N),data2conv2 =>d99_in (8*N-1 downto 7*N),data2conv3 =>d99_in (7*N-1 downto 6*N),data2conv4 =>d99_in (6*N-1 downto 5*N),data2conv5 =>d99_in (5*N-1 downto 4*N),data2conv6 =>d99_in (4*N-1 downto 3*N),data2conv7 =>d99_in (3*N-1 downto 2*N),data2conv8 =>d99_in (2*N-1 downto N),data2conv9 =>d99_in (N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d99_in (9*N-1 downto 8*N),w2 => d99_in (8*N-1 downto 7*N),w3 => d99_in (7*N-1 downto 6*N),w4 => d99_in (6*N-1 downto 5*N),w5 => d99_in (5*N-1 downto 4*N),w6 => d99_in (4*N-1 downto 3*N),w7 => d99_in (3*N-1 downto 2*N),w8 => d99_in (2*N-1 downto N),w9 => d99_in (N-1 downto 0 ),d_out => d99_out ,en_out =>open  ,sof_out=>open   );
CL100: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d100_in(9*N-1 downto 8*N),data2conv2 =>d100_in(8*N-1 downto 7*N),data2conv3 =>d100_in(7*N-1 downto 6*N),data2conv4 =>d100_in(6*N-1 downto 5*N),data2conv5 =>d100_in(5*N-1 downto 4*N),data2conv6 =>d100_in(4*N-1 downto 3*N),data2conv7 =>d100_in(3*N-1 downto 2*N),data2conv8 =>d100_in(2*N-1 downto N),data2conv9 =>d100_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d100_in(9*N-1 downto 8*N),w2 => d100_in(8*N-1 downto 7*N),w3 => d100_in(7*N-1 downto 6*N),w4 => d100_in(6*N-1 downto 5*N),w5 => d100_in(5*N-1 downto 4*N),w6 => d100_in(4*N-1 downto 3*N),w7 => d100_in(3*N-1 downto 2*N),w8 => d100_in(2*N-1 downto N),w9 => d100_in(N-1 downto 0 ),d_out => d100_out,en_out =>open  ,sof_out=>open   );
CL101: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d101_in(9*N-1 downto 8*N),data2conv2 =>d101_in(8*N-1 downto 7*N),data2conv3 =>d101_in(7*N-1 downto 6*N),data2conv4 =>d101_in(6*N-1 downto 5*N),data2conv5 =>d101_in(5*N-1 downto 4*N),data2conv6 =>d101_in(4*N-1 downto 3*N),data2conv7 =>d101_in(3*N-1 downto 2*N),data2conv8 =>d101_in(2*N-1 downto N),data2conv9 =>d101_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d101_in(9*N-1 downto 8*N),w2 => d101_in(8*N-1 downto 7*N),w3 => d101_in(7*N-1 downto 6*N),w4 => d101_in(6*N-1 downto 5*N),w5 => d101_in(5*N-1 downto 4*N),w6 => d101_in(4*N-1 downto 3*N),w7 => d101_in(3*N-1 downto 2*N),w8 => d101_in(2*N-1 downto N),w9 => d101_in(N-1 downto 0 ),d_out => d101_out,en_out =>open  ,sof_out=>open   );
CL102: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d102_in(9*N-1 downto 8*N),data2conv2 =>d102_in(8*N-1 downto 7*N),data2conv3 =>d102_in(7*N-1 downto 6*N),data2conv4 =>d102_in(6*N-1 downto 5*N),data2conv5 =>d102_in(5*N-1 downto 4*N),data2conv6 =>d102_in(4*N-1 downto 3*N),data2conv7 =>d102_in(3*N-1 downto 2*N),data2conv8 =>d102_in(2*N-1 downto N),data2conv9 =>d102_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d102_in(9*N-1 downto 8*N),w2 => d102_in(8*N-1 downto 7*N),w3 => d102_in(7*N-1 downto 6*N),w4 => d102_in(6*N-1 downto 5*N),w5 => d102_in(5*N-1 downto 4*N),w6 => d102_in(4*N-1 downto 3*N),w7 => d102_in(3*N-1 downto 2*N),w8 => d102_in(2*N-1 downto N),w9 => d102_in(N-1 downto 0 ),d_out => d102_out,en_out =>open  ,sof_out=>open   );
CL103: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d103_in(9*N-1 downto 8*N),data2conv2 =>d103_in(8*N-1 downto 7*N),data2conv3 =>d103_in(7*N-1 downto 6*N),data2conv4 =>d103_in(6*N-1 downto 5*N),data2conv5 =>d103_in(5*N-1 downto 4*N),data2conv6 =>d103_in(4*N-1 downto 3*N),data2conv7 =>d103_in(3*N-1 downto 2*N),data2conv8 =>d103_in(2*N-1 downto N),data2conv9 =>d103_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d103_in(9*N-1 downto 8*N),w2 => d103_in(8*N-1 downto 7*N),w3 => d103_in(7*N-1 downto 6*N),w4 => d103_in(6*N-1 downto 5*N),w5 => d103_in(5*N-1 downto 4*N),w6 => d103_in(4*N-1 downto 3*N),w7 => d103_in(3*N-1 downto 2*N),w8 => d103_in(2*N-1 downto N),w9 => d103_in(N-1 downto 0 ),d_out => d103_out,en_out =>open  ,sof_out=>open   );
CL104: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d104_in(9*N-1 downto 8*N),data2conv2 =>d104_in(8*N-1 downto 7*N),data2conv3 =>d104_in(7*N-1 downto 6*N),data2conv4 =>d104_in(6*N-1 downto 5*N),data2conv5 =>d104_in(5*N-1 downto 4*N),data2conv6 =>d104_in(4*N-1 downto 3*N),data2conv7 =>d104_in(3*N-1 downto 2*N),data2conv8 =>d104_in(2*N-1 downto N),data2conv9 =>d104_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d104_in(9*N-1 downto 8*N),w2 => d104_in(8*N-1 downto 7*N),w3 => d104_in(7*N-1 downto 6*N),w4 => d104_in(6*N-1 downto 5*N),w5 => d104_in(5*N-1 downto 4*N),w6 => d104_in(4*N-1 downto 3*N),w7 => d104_in(3*N-1 downto 2*N),w8 => d104_in(2*N-1 downto N),w9 => d104_in(N-1 downto 0 ),d_out => d104_out,en_out =>open  ,sof_out=>open   );
CL105: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d105_in(9*N-1 downto 8*N),data2conv2 =>d105_in(8*N-1 downto 7*N),data2conv3 =>d105_in(7*N-1 downto 6*N),data2conv4 =>d105_in(6*N-1 downto 5*N),data2conv5 =>d105_in(5*N-1 downto 4*N),data2conv6 =>d105_in(4*N-1 downto 3*N),data2conv7 =>d105_in(3*N-1 downto 2*N),data2conv8 =>d105_in(2*N-1 downto N),data2conv9 =>d105_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d105_in(9*N-1 downto 8*N),w2 => d105_in(8*N-1 downto 7*N),w3 => d105_in(7*N-1 downto 6*N),w4 => d105_in(6*N-1 downto 5*N),w5 => d105_in(5*N-1 downto 4*N),w6 => d105_in(4*N-1 downto 3*N),w7 => d105_in(3*N-1 downto 2*N),w8 => d105_in(2*N-1 downto N),w9 => d105_in(N-1 downto 0 ),d_out => d105_out,en_out =>open  ,sof_out=>open   );
CL106: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d106_in(9*N-1 downto 8*N),data2conv2 =>d106_in(8*N-1 downto 7*N),data2conv3 =>d106_in(7*N-1 downto 6*N),data2conv4 =>d106_in(6*N-1 downto 5*N),data2conv5 =>d106_in(5*N-1 downto 4*N),data2conv6 =>d106_in(4*N-1 downto 3*N),data2conv7 =>d106_in(3*N-1 downto 2*N),data2conv8 =>d106_in(2*N-1 downto N),data2conv9 =>d106_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d106_in(9*N-1 downto 8*N),w2 => d106_in(8*N-1 downto 7*N),w3 => d106_in(7*N-1 downto 6*N),w4 => d106_in(6*N-1 downto 5*N),w5 => d106_in(5*N-1 downto 4*N),w6 => d106_in(4*N-1 downto 3*N),w7 => d106_in(3*N-1 downto 2*N),w8 => d106_in(2*N-1 downto N),w9 => d106_in(N-1 downto 0 ),d_out => d106_out,en_out =>open  ,sof_out=>open   );
CL107: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d107_in(9*N-1 downto 8*N),data2conv2 =>d107_in(8*N-1 downto 7*N),data2conv3 =>d107_in(7*N-1 downto 6*N),data2conv4 =>d107_in(6*N-1 downto 5*N),data2conv5 =>d107_in(5*N-1 downto 4*N),data2conv6 =>d107_in(4*N-1 downto 3*N),data2conv7 =>d107_in(3*N-1 downto 2*N),data2conv8 =>d107_in(2*N-1 downto N),data2conv9 =>d107_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d107_in(9*N-1 downto 8*N),w2 => d107_in(8*N-1 downto 7*N),w3 => d107_in(7*N-1 downto 6*N),w4 => d107_in(6*N-1 downto 5*N),w5 => d107_in(5*N-1 downto 4*N),w6 => d107_in(4*N-1 downto 3*N),w7 => d107_in(3*N-1 downto 2*N),w8 => d107_in(2*N-1 downto N),w9 => d107_in(N-1 downto 0 ),d_out => d107_out,en_out =>open  ,sof_out=>open   );
CL108: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d108_in(9*N-1 downto 8*N),data2conv2 =>d108_in(8*N-1 downto 7*N),data2conv3 =>d108_in(7*N-1 downto 6*N),data2conv4 =>d108_in(6*N-1 downto 5*N),data2conv5 =>d108_in(5*N-1 downto 4*N),data2conv6 =>d108_in(4*N-1 downto 3*N),data2conv7 =>d108_in(3*N-1 downto 2*N),data2conv8 =>d108_in(2*N-1 downto N),data2conv9 =>d108_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d108_in(9*N-1 downto 8*N),w2 => d108_in(8*N-1 downto 7*N),w3 => d108_in(7*N-1 downto 6*N),w4 => d108_in(6*N-1 downto 5*N),w5 => d108_in(5*N-1 downto 4*N),w6 => d108_in(4*N-1 downto 3*N),w7 => d108_in(3*N-1 downto 2*N),w8 => d108_in(2*N-1 downto N),w9 => d108_in(N-1 downto 0 ),d_out => d108_out,en_out =>open  ,sof_out=>open   );
CL109: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d109_in(9*N-1 downto 8*N),data2conv2 =>d109_in(8*N-1 downto 7*N),data2conv3 =>d109_in(7*N-1 downto 6*N),data2conv4 =>d109_in(6*N-1 downto 5*N),data2conv5 =>d109_in(5*N-1 downto 4*N),data2conv6 =>d109_in(4*N-1 downto 3*N),data2conv7 =>d109_in(3*N-1 downto 2*N),data2conv8 =>d109_in(2*N-1 downto N),data2conv9 =>d109_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d109_in(9*N-1 downto 8*N),w2 => d109_in(8*N-1 downto 7*N),w3 => d109_in(7*N-1 downto 6*N),w4 => d109_in(6*N-1 downto 5*N),w5 => d109_in(5*N-1 downto 4*N),w6 => d109_in(4*N-1 downto 3*N),w7 => d109_in(3*N-1 downto 2*N),w8 => d109_in(2*N-1 downto N),w9 => d109_in(N-1 downto 0 ),d_out => d109_out,en_out =>open  ,sof_out=>open   );
CL110: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d110_in(9*N-1 downto 8*N),data2conv2 =>d110_in(8*N-1 downto 7*N),data2conv3 =>d110_in(7*N-1 downto 6*N),data2conv4 =>d110_in(6*N-1 downto 5*N),data2conv5 =>d110_in(5*N-1 downto 4*N),data2conv6 =>d110_in(4*N-1 downto 3*N),data2conv7 =>d110_in(3*N-1 downto 2*N),data2conv8 =>d110_in(2*N-1 downto N),data2conv9 =>d110_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d110_in(9*N-1 downto 8*N),w2 => d110_in(8*N-1 downto 7*N),w3 => d110_in(7*N-1 downto 6*N),w4 => d110_in(6*N-1 downto 5*N),w5 => d110_in(5*N-1 downto 4*N),w6 => d110_in(4*N-1 downto 3*N),w7 => d110_in(3*N-1 downto 2*N),w8 => d110_in(2*N-1 downto N),w9 => d110_in(N-1 downto 0 ),d_out => d110_out,en_out =>open  ,sof_out=>open   );
CL111: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d111_in(9*N-1 downto 8*N),data2conv2 =>d111_in(8*N-1 downto 7*N),data2conv3 =>d111_in(7*N-1 downto 6*N),data2conv4 =>d111_in(6*N-1 downto 5*N),data2conv5 =>d111_in(5*N-1 downto 4*N),data2conv6 =>d111_in(4*N-1 downto 3*N),data2conv7 =>d111_in(3*N-1 downto 2*N),data2conv8 =>d111_in(2*N-1 downto N),data2conv9 =>d111_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d111_in(9*N-1 downto 8*N),w2 => d111_in(8*N-1 downto 7*N),w3 => d111_in(7*N-1 downto 6*N),w4 => d111_in(6*N-1 downto 5*N),w5 => d111_in(5*N-1 downto 4*N),w6 => d111_in(4*N-1 downto 3*N),w7 => d111_in(3*N-1 downto 2*N),w8 => d111_in(2*N-1 downto N),w9 => d111_in(N-1 downto 0 ),d_out => d111_out,en_out =>open  ,sof_out=>open   );
CL112: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d112_in(9*N-1 downto 8*N),data2conv2 =>d112_in(8*N-1 downto 7*N),data2conv3 =>d112_in(7*N-1 downto 6*N),data2conv4 =>d112_in(6*N-1 downto 5*N),data2conv5 =>d112_in(5*N-1 downto 4*N),data2conv6 =>d112_in(4*N-1 downto 3*N),data2conv7 =>d112_in(3*N-1 downto 2*N),data2conv8 =>d112_in(2*N-1 downto N),data2conv9 =>d112_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d112_in(9*N-1 downto 8*N),w2 => d112_in(8*N-1 downto 7*N),w3 => d112_in(7*N-1 downto 6*N),w4 => d112_in(6*N-1 downto 5*N),w5 => d112_in(5*N-1 downto 4*N),w6 => d112_in(4*N-1 downto 3*N),w7 => d112_in(3*N-1 downto 2*N),w8 => d112_in(2*N-1 downto N),w9 => d112_in(N-1 downto 0 ),d_out => d112_out,en_out =>open  ,sof_out=>open   );
CL113: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d113_in(9*N-1 downto 8*N),data2conv2 =>d113_in(8*N-1 downto 7*N),data2conv3 =>d113_in(7*N-1 downto 6*N),data2conv4 =>d113_in(6*N-1 downto 5*N),data2conv5 =>d113_in(5*N-1 downto 4*N),data2conv6 =>d113_in(4*N-1 downto 3*N),data2conv7 =>d113_in(3*N-1 downto 2*N),data2conv8 =>d113_in(2*N-1 downto N),data2conv9 =>d113_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d113_in(9*N-1 downto 8*N),w2 => d113_in(8*N-1 downto 7*N),w3 => d113_in(7*N-1 downto 6*N),w4 => d113_in(6*N-1 downto 5*N),w5 => d113_in(5*N-1 downto 4*N),w6 => d113_in(4*N-1 downto 3*N),w7 => d113_in(3*N-1 downto 2*N),w8 => d113_in(2*N-1 downto N),w9 => d113_in(N-1 downto 0 ),d_out => d113_out,en_out =>open  ,sof_out=>open   );
CL114: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d114_in(9*N-1 downto 8*N),data2conv2 =>d114_in(8*N-1 downto 7*N),data2conv3 =>d114_in(7*N-1 downto 6*N),data2conv4 =>d114_in(6*N-1 downto 5*N),data2conv5 =>d114_in(5*N-1 downto 4*N),data2conv6 =>d114_in(4*N-1 downto 3*N),data2conv7 =>d114_in(3*N-1 downto 2*N),data2conv8 =>d114_in(2*N-1 downto N),data2conv9 =>d114_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d114_in(9*N-1 downto 8*N),w2 => d114_in(8*N-1 downto 7*N),w3 => d114_in(7*N-1 downto 6*N),w4 => d114_in(6*N-1 downto 5*N),w5 => d114_in(5*N-1 downto 4*N),w6 => d114_in(4*N-1 downto 3*N),w7 => d114_in(3*N-1 downto 2*N),w8 => d114_in(2*N-1 downto N),w9 => d114_in(N-1 downto 0 ),d_out => d114_out,en_out =>open  ,sof_out=>open   );
CL115: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d115_in(9*N-1 downto 8*N),data2conv2 =>d115_in(8*N-1 downto 7*N),data2conv3 =>d115_in(7*N-1 downto 6*N),data2conv4 =>d115_in(6*N-1 downto 5*N),data2conv5 =>d115_in(5*N-1 downto 4*N),data2conv6 =>d115_in(4*N-1 downto 3*N),data2conv7 =>d115_in(3*N-1 downto 2*N),data2conv8 =>d115_in(2*N-1 downto N),data2conv9 =>d115_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d115_in(9*N-1 downto 8*N),w2 => d115_in(8*N-1 downto 7*N),w3 => d115_in(7*N-1 downto 6*N),w4 => d115_in(6*N-1 downto 5*N),w5 => d115_in(5*N-1 downto 4*N),w6 => d115_in(4*N-1 downto 3*N),w7 => d115_in(3*N-1 downto 2*N),w8 => d115_in(2*N-1 downto N),w9 => d115_in(N-1 downto 0 ),d_out => d115_out,en_out =>open  ,sof_out=>open   );
CL116: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d116_in(9*N-1 downto 8*N),data2conv2 =>d116_in(8*N-1 downto 7*N),data2conv3 =>d116_in(7*N-1 downto 6*N),data2conv4 =>d116_in(6*N-1 downto 5*N),data2conv5 =>d116_in(5*N-1 downto 4*N),data2conv6 =>d116_in(4*N-1 downto 3*N),data2conv7 =>d116_in(3*N-1 downto 2*N),data2conv8 =>d116_in(2*N-1 downto N),data2conv9 =>d116_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d116_in(9*N-1 downto 8*N),w2 => d116_in(8*N-1 downto 7*N),w3 => d116_in(7*N-1 downto 6*N),w4 => d116_in(6*N-1 downto 5*N),w5 => d116_in(5*N-1 downto 4*N),w6 => d116_in(4*N-1 downto 3*N),w7 => d116_in(3*N-1 downto 2*N),w8 => d116_in(2*N-1 downto N),w9 => d116_in(N-1 downto 0 ),d_out => d116_out,en_out =>open  ,sof_out=>open   );
CL117: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d117_in(9*N-1 downto 8*N),data2conv2 =>d117_in(8*N-1 downto 7*N),data2conv3 =>d117_in(7*N-1 downto 6*N),data2conv4 =>d117_in(6*N-1 downto 5*N),data2conv5 =>d117_in(5*N-1 downto 4*N),data2conv6 =>d117_in(4*N-1 downto 3*N),data2conv7 =>d117_in(3*N-1 downto 2*N),data2conv8 =>d117_in(2*N-1 downto N),data2conv9 =>d117_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d117_in(9*N-1 downto 8*N),w2 => d117_in(8*N-1 downto 7*N),w3 => d117_in(7*N-1 downto 6*N),w4 => d117_in(6*N-1 downto 5*N),w5 => d117_in(5*N-1 downto 4*N),w6 => d117_in(4*N-1 downto 3*N),w7 => d117_in(3*N-1 downto 2*N),w8 => d117_in(2*N-1 downto N),w9 => d117_in(N-1 downto 0 ),d_out => d117_out,en_out =>open  ,sof_out=>open   );
CL118: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d118_in(9*N-1 downto 8*N),data2conv2 =>d118_in(8*N-1 downto 7*N),data2conv3 =>d118_in(7*N-1 downto 6*N),data2conv4 =>d118_in(6*N-1 downto 5*N),data2conv5 =>d118_in(5*N-1 downto 4*N),data2conv6 =>d118_in(4*N-1 downto 3*N),data2conv7 =>d118_in(3*N-1 downto 2*N),data2conv8 =>d118_in(2*N-1 downto N),data2conv9 =>d118_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d118_in(9*N-1 downto 8*N),w2 => d118_in(8*N-1 downto 7*N),w3 => d118_in(7*N-1 downto 6*N),w4 => d118_in(6*N-1 downto 5*N),w5 => d118_in(5*N-1 downto 4*N),w6 => d118_in(4*N-1 downto 3*N),w7 => d118_in(3*N-1 downto 2*N),w8 => d118_in(2*N-1 downto N),w9 => d118_in(N-1 downto 0 ),d_out => d118_out,en_out =>open  ,sof_out=>open   );
CL119: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d119_in(9*N-1 downto 8*N),data2conv2 =>d119_in(8*N-1 downto 7*N),data2conv3 =>d119_in(7*N-1 downto 6*N),data2conv4 =>d119_in(6*N-1 downto 5*N),data2conv5 =>d119_in(5*N-1 downto 4*N),data2conv6 =>d119_in(4*N-1 downto 3*N),data2conv7 =>d119_in(3*N-1 downto 2*N),data2conv8 =>d119_in(2*N-1 downto N),data2conv9 =>d119_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d119_in(9*N-1 downto 8*N),w2 => d119_in(8*N-1 downto 7*N),w3 => d119_in(7*N-1 downto 6*N),w4 => d119_in(6*N-1 downto 5*N),w5 => d119_in(5*N-1 downto 4*N),w6 => d119_in(4*N-1 downto 3*N),w7 => d119_in(3*N-1 downto 2*N),w8 => d119_in(2*N-1 downto N),w9 => d119_in(N-1 downto 0 ),d_out => d119_out,en_out =>open  ,sof_out=>open   );
CL120: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d120_in(9*N-1 downto 8*N),data2conv2 =>d120_in(8*N-1 downto 7*N),data2conv3 =>d120_in(7*N-1 downto 6*N),data2conv4 =>d120_in(6*N-1 downto 5*N),data2conv5 =>d120_in(5*N-1 downto 4*N),data2conv6 =>d120_in(4*N-1 downto 3*N),data2conv7 =>d120_in(3*N-1 downto 2*N),data2conv8 =>d120_in(2*N-1 downto N),data2conv9 =>d120_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d120_in(9*N-1 downto 8*N),w2 => d120_in(8*N-1 downto 7*N),w3 => d120_in(7*N-1 downto 6*N),w4 => d120_in(6*N-1 downto 5*N),w5 => d120_in(5*N-1 downto 4*N),w6 => d120_in(4*N-1 downto 3*N),w7 => d120_in(3*N-1 downto 2*N),w8 => d120_in(2*N-1 downto N),w9 => d120_in(N-1 downto 0 ),d_out => d120_out,en_out =>open  ,sof_out=>open   );
CL121: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d121_in(9*N-1 downto 8*N),data2conv2 =>d121_in(8*N-1 downto 7*N),data2conv3 =>d121_in(7*N-1 downto 6*N),data2conv4 =>d121_in(6*N-1 downto 5*N),data2conv5 =>d121_in(5*N-1 downto 4*N),data2conv6 =>d121_in(4*N-1 downto 3*N),data2conv7 =>d121_in(3*N-1 downto 2*N),data2conv8 =>d121_in(2*N-1 downto N),data2conv9 =>d121_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d121_in(9*N-1 downto 8*N),w2 => d121_in(8*N-1 downto 7*N),w3 => d121_in(7*N-1 downto 6*N),w4 => d121_in(6*N-1 downto 5*N),w5 => d121_in(5*N-1 downto 4*N),w6 => d121_in(4*N-1 downto 3*N),w7 => d121_in(3*N-1 downto 2*N),w8 => d121_in(2*N-1 downto N),w9 => d121_in(N-1 downto 0 ),d_out => d121_out,en_out =>open  ,sof_out=>open   );
CL122: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d122_in(9*N-1 downto 8*N),data2conv2 =>d122_in(8*N-1 downto 7*N),data2conv3 =>d122_in(7*N-1 downto 6*N),data2conv4 =>d122_in(6*N-1 downto 5*N),data2conv5 =>d122_in(5*N-1 downto 4*N),data2conv6 =>d122_in(4*N-1 downto 3*N),data2conv7 =>d122_in(3*N-1 downto 2*N),data2conv8 =>d122_in(2*N-1 downto N),data2conv9 =>d122_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d122_in(9*N-1 downto 8*N),w2 => d122_in(8*N-1 downto 7*N),w3 => d122_in(7*N-1 downto 6*N),w4 => d122_in(6*N-1 downto 5*N),w5 => d122_in(5*N-1 downto 4*N),w6 => d122_in(4*N-1 downto 3*N),w7 => d122_in(3*N-1 downto 2*N),w8 => d122_in(2*N-1 downto N),w9 => d122_in(N-1 downto 0 ),d_out => d122_out,en_out =>open  ,sof_out=>open   );
CL123: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d123_in(9*N-1 downto 8*N),data2conv2 =>d123_in(8*N-1 downto 7*N),data2conv3 =>d123_in(7*N-1 downto 6*N),data2conv4 =>d123_in(6*N-1 downto 5*N),data2conv5 =>d123_in(5*N-1 downto 4*N),data2conv6 =>d123_in(4*N-1 downto 3*N),data2conv7 =>d123_in(3*N-1 downto 2*N),data2conv8 =>d123_in(2*N-1 downto N),data2conv9 =>d123_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d123_in(9*N-1 downto 8*N),w2 => d123_in(8*N-1 downto 7*N),w3 => d123_in(7*N-1 downto 6*N),w4 => d123_in(6*N-1 downto 5*N),w5 => d123_in(5*N-1 downto 4*N),w6 => d123_in(4*N-1 downto 3*N),w7 => d123_in(3*N-1 downto 2*N),w8 => d123_in(2*N-1 downto N),w9 => d123_in(N-1 downto 0 ),d_out => d123_out,en_out =>open  ,sof_out=>open   );
CL124: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d124_in(9*N-1 downto 8*N),data2conv2 =>d124_in(8*N-1 downto 7*N),data2conv3 =>d124_in(7*N-1 downto 6*N),data2conv4 =>d124_in(6*N-1 downto 5*N),data2conv5 =>d124_in(5*N-1 downto 4*N),data2conv6 =>d124_in(4*N-1 downto 3*N),data2conv7 =>d124_in(3*N-1 downto 2*N),data2conv8 =>d124_in(2*N-1 downto N),data2conv9 =>d124_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d124_in(9*N-1 downto 8*N),w2 => d124_in(8*N-1 downto 7*N),w3 => d124_in(7*N-1 downto 6*N),w4 => d124_in(6*N-1 downto 5*N),w5 => d124_in(5*N-1 downto 4*N),w6 => d124_in(4*N-1 downto 3*N),w7 => d124_in(3*N-1 downto 2*N),w8 => d124_in(2*N-1 downto N),w9 => d124_in(N-1 downto 0 ),d_out => d124_out,en_out =>open  ,sof_out=>open   );
CL125: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d125_in(9*N-1 downto 8*N),data2conv2 =>d125_in(8*N-1 downto 7*N),data2conv3 =>d125_in(7*N-1 downto 6*N),data2conv4 =>d125_in(6*N-1 downto 5*N),data2conv5 =>d125_in(5*N-1 downto 4*N),data2conv6 =>d125_in(4*N-1 downto 3*N),data2conv7 =>d125_in(3*N-1 downto 2*N),data2conv8 =>d125_in(2*N-1 downto N),data2conv9 =>d125_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d125_in(9*N-1 downto 8*N),w2 => d125_in(8*N-1 downto 7*N),w3 => d125_in(7*N-1 downto 6*N),w4 => d125_in(6*N-1 downto 5*N),w5 => d125_in(5*N-1 downto 4*N),w6 => d125_in(4*N-1 downto 3*N),w7 => d125_in(3*N-1 downto 2*N),w8 => d125_in(2*N-1 downto N),w9 => d125_in(N-1 downto 0 ),d_out => d125_out,en_out =>open  ,sof_out=>open   );
CL126: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d126_in(9*N-1 downto 8*N),data2conv2 =>d126_in(8*N-1 downto 7*N),data2conv3 =>d126_in(7*N-1 downto 6*N),data2conv4 =>d126_in(6*N-1 downto 5*N),data2conv5 =>d126_in(5*N-1 downto 4*N),data2conv6 =>d126_in(4*N-1 downto 3*N),data2conv7 =>d126_in(3*N-1 downto 2*N),data2conv8 =>d126_in(2*N-1 downto N),data2conv9 =>d126_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d126_in(9*N-1 downto 8*N),w2 => d126_in(8*N-1 downto 7*N),w3 => d126_in(7*N-1 downto 6*N),w4 => d126_in(6*N-1 downto 5*N),w5 => d126_in(5*N-1 downto 4*N),w6 => d126_in(4*N-1 downto 3*N),w7 => d126_in(3*N-1 downto 2*N),w8 => d126_in(2*N-1 downto N),w9 => d126_in(N-1 downto 0 ),d_out => d126_out,en_out =>open  ,sof_out=>open   );
CL127: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d127_in(9*N-1 downto 8*N),data2conv2 =>d127_in(8*N-1 downto 7*N),data2conv3 =>d127_in(7*N-1 downto 6*N),data2conv4 =>d127_in(6*N-1 downto 5*N),data2conv5 =>d127_in(5*N-1 downto 4*N),data2conv6 =>d127_in(4*N-1 downto 3*N),data2conv7 =>d127_in(3*N-1 downto 2*N),data2conv8 =>d127_in(2*N-1 downto N),data2conv9 =>d127_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d127_in(9*N-1 downto 8*N),w2 => d127_in(8*N-1 downto 7*N),w3 => d127_in(7*N-1 downto 6*N),w4 => d127_in(6*N-1 downto 5*N),w5 => d127_in(5*N-1 downto 4*N),w6 => d127_in(4*N-1 downto 3*N),w7 => d127_in(3*N-1 downto 2*N),w8 => d127_in(2*N-1 downto N),w9 => d127_in(N-1 downto 0 ),d_out => d127_out,en_out =>open  ,sof_out=>open   );
CL128: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d128_in(9*N-1 downto 8*N),data2conv2 =>d128_in(8*N-1 downto 7*N),data2conv3 =>d128_in(7*N-1 downto 6*N),data2conv4 =>d128_in(6*N-1 downto 5*N),data2conv5 =>d128_in(5*N-1 downto 4*N),data2conv6 =>d128_in(4*N-1 downto 3*N),data2conv7 =>d128_in(3*N-1 downto 2*N),data2conv8 =>d128_in(2*N-1 downto N),data2conv9 =>d128_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d128_in(9*N-1 downto 8*N),w2 => d128_in(8*N-1 downto 7*N),w3 => d128_in(7*N-1 downto 6*N),w4 => d128_in(6*N-1 downto 5*N),w5 => d128_in(5*N-1 downto 4*N),w6 => d128_in(4*N-1 downto 3*N),w7 => d128_in(3*N-1 downto 2*N),w8 => d128_in(2*N-1 downto N),w9 => d128_in(N-1 downto 0 ),d_out => d128_out,en_out =>open  ,sof_out=>open   );


CL129: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d129_in(9*N-1 downto 8*N),data2conv2 =>d129_in(8*N-1 downto 7*N),data2conv3 =>d129_in(7*N-1 downto 6*N),data2conv4 =>d129_in(6*N-1 downto 5*N),data2conv5 =>d129_in(5*N-1 downto 4*N),data2conv6 =>d129_in(4*N-1 downto 3*N),data2conv7 =>d129_in(3*N-1 downto 2*N),data2conv8 =>d129_in(2*N-1 downto N),data2conv9 =>d129_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d129_in(9*N-1 downto 8*N),w2 => d129_in(8*N-1 downto 7*N),w3 => d129_in(7*N-1 downto 6*N),w4 => d129_in(6*N-1 downto 5*N),w5 => d129_in(5*N-1 downto 4*N),w6 => d129_in(4*N-1 downto 3*N),w7 => d129_in(3*N-1 downto 2*N),w8 => d129_in(2*N-1 downto N),w9 => d129_in(N-1 downto 0 ),d_out => d129_out,en_out =>open  ,sof_out=>open   );
CL130: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d130_in(9*N-1 downto 8*N),data2conv2 =>d130_in(8*N-1 downto 7*N),data2conv3 =>d130_in(7*N-1 downto 6*N),data2conv4 =>d130_in(6*N-1 downto 5*N),data2conv5 =>d130_in(5*N-1 downto 4*N),data2conv6 =>d130_in(4*N-1 downto 3*N),data2conv7 =>d130_in(3*N-1 downto 2*N),data2conv8 =>d130_in(2*N-1 downto N),data2conv9 =>d130_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d130_in(9*N-1 downto 8*N),w2 => d130_in(8*N-1 downto 7*N),w3 => d130_in(7*N-1 downto 6*N),w4 => d130_in(6*N-1 downto 5*N),w5 => d130_in(5*N-1 downto 4*N),w6 => d130_in(4*N-1 downto 3*N),w7 => d130_in(3*N-1 downto 2*N),w8 => d130_in(2*N-1 downto N),w9 => d130_in(N-1 downto 0 ),d_out => d130_out,en_out =>open  ,sof_out=>open   );
CL131: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d131_in(9*N-1 downto 8*N),data2conv2 =>d131_in(8*N-1 downto 7*N),data2conv3 =>d131_in(7*N-1 downto 6*N),data2conv4 =>d131_in(6*N-1 downto 5*N),data2conv5 =>d131_in(5*N-1 downto 4*N),data2conv6 =>d131_in(4*N-1 downto 3*N),data2conv7 =>d131_in(3*N-1 downto 2*N),data2conv8 =>d131_in(2*N-1 downto N),data2conv9 =>d131_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d131_in(9*N-1 downto 8*N),w2 => d131_in(8*N-1 downto 7*N),w3 => d131_in(7*N-1 downto 6*N),w4 => d131_in(6*N-1 downto 5*N),w5 => d131_in(5*N-1 downto 4*N),w6 => d131_in(4*N-1 downto 3*N),w7 => d131_in(3*N-1 downto 2*N),w8 => d131_in(2*N-1 downto N),w9 => d131_in(N-1 downto 0 ),d_out => d131_out,en_out =>open  ,sof_out=>open   );
CL132: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d132_in(9*N-1 downto 8*N),data2conv2 =>d132_in(8*N-1 downto 7*N),data2conv3 =>d132_in(7*N-1 downto 6*N),data2conv4 =>d132_in(6*N-1 downto 5*N),data2conv5 =>d132_in(5*N-1 downto 4*N),data2conv6 =>d132_in(4*N-1 downto 3*N),data2conv7 =>d132_in(3*N-1 downto 2*N),data2conv8 =>d132_in(2*N-1 downto N),data2conv9 =>d132_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d132_in(9*N-1 downto 8*N),w2 => d132_in(8*N-1 downto 7*N),w3 => d132_in(7*N-1 downto 6*N),w4 => d132_in(6*N-1 downto 5*N),w5 => d132_in(5*N-1 downto 4*N),w6 => d132_in(4*N-1 downto 3*N),w7 => d132_in(3*N-1 downto 2*N),w8 => d132_in(2*N-1 downto N),w9 => d132_in(N-1 downto 0 ),d_out => d132_out,en_out =>open  ,sof_out=>open   );
CL133: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d133_in(9*N-1 downto 8*N),data2conv2 =>d133_in(8*N-1 downto 7*N),data2conv3 =>d133_in(7*N-1 downto 6*N),data2conv4 =>d133_in(6*N-1 downto 5*N),data2conv5 =>d133_in(5*N-1 downto 4*N),data2conv6 =>d133_in(4*N-1 downto 3*N),data2conv7 =>d133_in(3*N-1 downto 2*N),data2conv8 =>d133_in(2*N-1 downto N),data2conv9 =>d133_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d133_in(9*N-1 downto 8*N),w2 => d133_in(8*N-1 downto 7*N),w3 => d133_in(7*N-1 downto 6*N),w4 => d133_in(6*N-1 downto 5*N),w5 => d133_in(5*N-1 downto 4*N),w6 => d133_in(4*N-1 downto 3*N),w7 => d133_in(3*N-1 downto 2*N),w8 => d133_in(2*N-1 downto N),w9 => d133_in(N-1 downto 0 ),d_out => d133_out,en_out =>open  ,sof_out=>open   );
CL134: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d134_in(9*N-1 downto 8*N),data2conv2 =>d134_in(8*N-1 downto 7*N),data2conv3 =>d134_in(7*N-1 downto 6*N),data2conv4 =>d134_in(6*N-1 downto 5*N),data2conv5 =>d134_in(5*N-1 downto 4*N),data2conv6 =>d134_in(4*N-1 downto 3*N),data2conv7 =>d134_in(3*N-1 downto 2*N),data2conv8 =>d134_in(2*N-1 downto N),data2conv9 =>d134_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d134_in(9*N-1 downto 8*N),w2 => d134_in(8*N-1 downto 7*N),w3 => d134_in(7*N-1 downto 6*N),w4 => d134_in(6*N-1 downto 5*N),w5 => d134_in(5*N-1 downto 4*N),w6 => d134_in(4*N-1 downto 3*N),w7 => d134_in(3*N-1 downto 2*N),w8 => d134_in(2*N-1 downto N),w9 => d134_in(N-1 downto 0 ),d_out => d134_out,en_out =>open  ,sof_out=>open   );
CL135: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d135_in(9*N-1 downto 8*N),data2conv2 =>d135_in(8*N-1 downto 7*N),data2conv3 =>d135_in(7*N-1 downto 6*N),data2conv4 =>d135_in(6*N-1 downto 5*N),data2conv5 =>d135_in(5*N-1 downto 4*N),data2conv6 =>d135_in(4*N-1 downto 3*N),data2conv7 =>d135_in(3*N-1 downto 2*N),data2conv8 =>d135_in(2*N-1 downto N),data2conv9 =>d135_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d135_in(9*N-1 downto 8*N),w2 => d135_in(8*N-1 downto 7*N),w3 => d135_in(7*N-1 downto 6*N),w4 => d135_in(6*N-1 downto 5*N),w5 => d135_in(5*N-1 downto 4*N),w6 => d135_in(4*N-1 downto 3*N),w7 => d135_in(3*N-1 downto 2*N),w8 => d135_in(2*N-1 downto N),w9 => d135_in(N-1 downto 0 ),d_out => d135_out,en_out =>open  ,sof_out=>open   );
CL136: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d136_in(9*N-1 downto 8*N),data2conv2 =>d136_in(8*N-1 downto 7*N),data2conv3 =>d136_in(7*N-1 downto 6*N),data2conv4 =>d136_in(6*N-1 downto 5*N),data2conv5 =>d136_in(5*N-1 downto 4*N),data2conv6 =>d136_in(4*N-1 downto 3*N),data2conv7 =>d136_in(3*N-1 downto 2*N),data2conv8 =>d136_in(2*N-1 downto N),data2conv9 =>d136_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d136_in(9*N-1 downto 8*N),w2 => d136_in(8*N-1 downto 7*N),w3 => d136_in(7*N-1 downto 6*N),w4 => d136_in(6*N-1 downto 5*N),w5 => d136_in(5*N-1 downto 4*N),w6 => d136_in(4*N-1 downto 3*N),w7 => d136_in(3*N-1 downto 2*N),w8 => d136_in(2*N-1 downto N),w9 => d136_in(N-1 downto 0 ),d_out => d136_out,en_out =>open  ,sof_out=>open   );
CL137: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d137_in(9*N-1 downto 8*N),data2conv2 =>d137_in(8*N-1 downto 7*N),data2conv3 =>d137_in(7*N-1 downto 6*N),data2conv4 =>d137_in(6*N-1 downto 5*N),data2conv5 =>d137_in(5*N-1 downto 4*N),data2conv6 =>d137_in(4*N-1 downto 3*N),data2conv7 =>d137_in(3*N-1 downto 2*N),data2conv8 =>d137_in(2*N-1 downto N),data2conv9 =>d137_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d137_in(9*N-1 downto 8*N),w2 => d137_in(8*N-1 downto 7*N),w3 => d137_in(7*N-1 downto 6*N),w4 => d137_in(6*N-1 downto 5*N),w5 => d137_in(5*N-1 downto 4*N),w6 => d137_in(4*N-1 downto 3*N),w7 => d137_in(3*N-1 downto 2*N),w8 => d137_in(2*N-1 downto N),w9 => d137_in(N-1 downto 0 ),d_out => d137_out,en_out =>open  ,sof_out=>open   );
CL138: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d138_in(9*N-1 downto 8*N),data2conv2 =>d138_in(8*N-1 downto 7*N),data2conv3 =>d138_in(7*N-1 downto 6*N),data2conv4 =>d138_in(6*N-1 downto 5*N),data2conv5 =>d138_in(5*N-1 downto 4*N),data2conv6 =>d138_in(4*N-1 downto 3*N),data2conv7 =>d138_in(3*N-1 downto 2*N),data2conv8 =>d138_in(2*N-1 downto N),data2conv9 =>d138_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d138_in(9*N-1 downto 8*N),w2 => d138_in(8*N-1 downto 7*N),w3 => d138_in(7*N-1 downto 6*N),w4 => d138_in(6*N-1 downto 5*N),w5 => d138_in(5*N-1 downto 4*N),w6 => d138_in(4*N-1 downto 3*N),w7 => d138_in(3*N-1 downto 2*N),w8 => d138_in(2*N-1 downto N),w9 => d138_in(N-1 downto 0 ),d_out => d138_out,en_out =>open  ,sof_out=>open   );
CL139: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d139_in(9*N-1 downto 8*N),data2conv2 =>d139_in(8*N-1 downto 7*N),data2conv3 =>d139_in(7*N-1 downto 6*N),data2conv4 =>d139_in(6*N-1 downto 5*N),data2conv5 =>d139_in(5*N-1 downto 4*N),data2conv6 =>d139_in(4*N-1 downto 3*N),data2conv7 =>d139_in(3*N-1 downto 2*N),data2conv8 =>d139_in(2*N-1 downto N),data2conv9 =>d139_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d139_in(9*N-1 downto 8*N),w2 => d139_in(8*N-1 downto 7*N),w3 => d139_in(7*N-1 downto 6*N),w4 => d139_in(6*N-1 downto 5*N),w5 => d139_in(5*N-1 downto 4*N),w6 => d139_in(4*N-1 downto 3*N),w7 => d139_in(3*N-1 downto 2*N),w8 => d139_in(2*N-1 downto N),w9 => d139_in(N-1 downto 0 ),d_out => d139_out,en_out =>open  ,sof_out=>open   );
CL140: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d140_in(9*N-1 downto 8*N),data2conv2 =>d140_in(8*N-1 downto 7*N),data2conv3 =>d140_in(7*N-1 downto 6*N),data2conv4 =>d140_in(6*N-1 downto 5*N),data2conv5 =>d140_in(5*N-1 downto 4*N),data2conv6 =>d140_in(4*N-1 downto 3*N),data2conv7 =>d140_in(3*N-1 downto 2*N),data2conv8 =>d140_in(2*N-1 downto N),data2conv9 =>d140_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d140_in(9*N-1 downto 8*N),w2 => d140_in(8*N-1 downto 7*N),w3 => d140_in(7*N-1 downto 6*N),w4 => d140_in(6*N-1 downto 5*N),w5 => d140_in(5*N-1 downto 4*N),w6 => d140_in(4*N-1 downto 3*N),w7 => d140_in(3*N-1 downto 2*N),w8 => d140_in(2*N-1 downto N),w9 => d140_in(N-1 downto 0 ),d_out => d140_out,en_out =>open  ,sof_out=>open   );
CL141: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d141_in(9*N-1 downto 8*N),data2conv2 =>d141_in(8*N-1 downto 7*N),data2conv3 =>d141_in(7*N-1 downto 6*N),data2conv4 =>d141_in(6*N-1 downto 5*N),data2conv5 =>d141_in(5*N-1 downto 4*N),data2conv6 =>d141_in(4*N-1 downto 3*N),data2conv7 =>d141_in(3*N-1 downto 2*N),data2conv8 =>d141_in(2*N-1 downto N),data2conv9 =>d141_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d141_in(9*N-1 downto 8*N),w2 => d141_in(8*N-1 downto 7*N),w3 => d141_in(7*N-1 downto 6*N),w4 => d141_in(6*N-1 downto 5*N),w5 => d141_in(5*N-1 downto 4*N),w6 => d141_in(4*N-1 downto 3*N),w7 => d141_in(3*N-1 downto 2*N),w8 => d141_in(2*N-1 downto N),w9 => d141_in(N-1 downto 0 ),d_out => d141_out,en_out =>open  ,sof_out=>open   );
CL142: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d142_in(9*N-1 downto 8*N),data2conv2 =>d142_in(8*N-1 downto 7*N),data2conv3 =>d142_in(7*N-1 downto 6*N),data2conv4 =>d142_in(6*N-1 downto 5*N),data2conv5 =>d142_in(5*N-1 downto 4*N),data2conv6 =>d142_in(4*N-1 downto 3*N),data2conv7 =>d142_in(3*N-1 downto 2*N),data2conv8 =>d142_in(2*N-1 downto N),data2conv9 =>d142_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d142_in(9*N-1 downto 8*N),w2 => d142_in(8*N-1 downto 7*N),w3 => d142_in(7*N-1 downto 6*N),w4 => d142_in(6*N-1 downto 5*N),w5 => d142_in(5*N-1 downto 4*N),w6 => d142_in(4*N-1 downto 3*N),w7 => d142_in(3*N-1 downto 2*N),w8 => d142_in(2*N-1 downto N),w9 => d142_in(N-1 downto 0 ),d_out => d142_out,en_out =>open  ,sof_out=>open   );
CL143: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d143_in(9*N-1 downto 8*N),data2conv2 =>d143_in(8*N-1 downto 7*N),data2conv3 =>d143_in(7*N-1 downto 6*N),data2conv4 =>d143_in(6*N-1 downto 5*N),data2conv5 =>d143_in(5*N-1 downto 4*N),data2conv6 =>d143_in(4*N-1 downto 3*N),data2conv7 =>d143_in(3*N-1 downto 2*N),data2conv8 =>d143_in(2*N-1 downto N),data2conv9 =>d143_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d143_in(9*N-1 downto 8*N),w2 => d143_in(8*N-1 downto 7*N),w3 => d143_in(7*N-1 downto 6*N),w4 => d143_in(6*N-1 downto 5*N),w5 => d143_in(5*N-1 downto 4*N),w6 => d143_in(4*N-1 downto 3*N),w7 => d143_in(3*N-1 downto 2*N),w8 => d143_in(2*N-1 downto N),w9 => d143_in(N-1 downto 0 ),d_out => d143_out,en_out =>open  ,sof_out=>open   );
CL144: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d144_in(9*N-1 downto 8*N),data2conv2 =>d144_in(8*N-1 downto 7*N),data2conv3 =>d144_in(7*N-1 downto 6*N),data2conv4 =>d144_in(6*N-1 downto 5*N),data2conv5 =>d144_in(5*N-1 downto 4*N),data2conv6 =>d144_in(4*N-1 downto 3*N),data2conv7 =>d144_in(3*N-1 downto 2*N),data2conv8 =>d144_in(2*N-1 downto N),data2conv9 =>d144_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d144_in(9*N-1 downto 8*N),w2 => d144_in(8*N-1 downto 7*N),w3 => d144_in(7*N-1 downto 6*N),w4 => d144_in(6*N-1 downto 5*N),w5 => d144_in(5*N-1 downto 4*N),w6 => d144_in(4*N-1 downto 3*N),w7 => d144_in(3*N-1 downto 2*N),w8 => d144_in(2*N-1 downto N),w9 => d144_in(N-1 downto 0 ),d_out => d144_out,en_out =>open  ,sof_out=>open   );
CL145: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d145_in(9*N-1 downto 8*N),data2conv2 =>d145_in(8*N-1 downto 7*N),data2conv3 =>d145_in(7*N-1 downto 6*N),data2conv4 =>d145_in(6*N-1 downto 5*N),data2conv5 =>d145_in(5*N-1 downto 4*N),data2conv6 =>d145_in(4*N-1 downto 3*N),data2conv7 =>d145_in(3*N-1 downto 2*N),data2conv8 =>d145_in(2*N-1 downto N),data2conv9 =>d145_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d145_in(9*N-1 downto 8*N),w2 => d145_in(8*N-1 downto 7*N),w3 => d145_in(7*N-1 downto 6*N),w4 => d145_in(6*N-1 downto 5*N),w5 => d145_in(5*N-1 downto 4*N),w6 => d145_in(4*N-1 downto 3*N),w7 => d145_in(3*N-1 downto 2*N),w8 => d145_in(2*N-1 downto N),w9 => d145_in(N-1 downto 0 ),d_out => d145_out,en_out =>open  ,sof_out=>open   );
CL146: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d146_in(9*N-1 downto 8*N),data2conv2 =>d146_in(8*N-1 downto 7*N),data2conv3 =>d146_in(7*N-1 downto 6*N),data2conv4 =>d146_in(6*N-1 downto 5*N),data2conv5 =>d146_in(5*N-1 downto 4*N),data2conv6 =>d146_in(4*N-1 downto 3*N),data2conv7 =>d146_in(3*N-1 downto 2*N),data2conv8 =>d146_in(2*N-1 downto N),data2conv9 =>d146_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d146_in(9*N-1 downto 8*N),w2 => d146_in(8*N-1 downto 7*N),w3 => d146_in(7*N-1 downto 6*N),w4 => d146_in(6*N-1 downto 5*N),w5 => d146_in(5*N-1 downto 4*N),w6 => d146_in(4*N-1 downto 3*N),w7 => d146_in(3*N-1 downto 2*N),w8 => d146_in(2*N-1 downto N),w9 => d146_in(N-1 downto 0 ),d_out => d146_out,en_out =>open  ,sof_out=>open   );
CL147: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d147_in(9*N-1 downto 8*N),data2conv2 =>d147_in(8*N-1 downto 7*N),data2conv3 =>d147_in(7*N-1 downto 6*N),data2conv4 =>d147_in(6*N-1 downto 5*N),data2conv5 =>d147_in(5*N-1 downto 4*N),data2conv6 =>d147_in(4*N-1 downto 3*N),data2conv7 =>d147_in(3*N-1 downto 2*N),data2conv8 =>d147_in(2*N-1 downto N),data2conv9 =>d147_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d147_in(9*N-1 downto 8*N),w2 => d147_in(8*N-1 downto 7*N),w3 => d147_in(7*N-1 downto 6*N),w4 => d147_in(6*N-1 downto 5*N),w5 => d147_in(5*N-1 downto 4*N),w6 => d147_in(4*N-1 downto 3*N),w7 => d147_in(3*N-1 downto 2*N),w8 => d147_in(2*N-1 downto N),w9 => d147_in(N-1 downto 0 ),d_out => d147_out,en_out =>open  ,sof_out=>open   );
CL148: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d148_in(9*N-1 downto 8*N),data2conv2 =>d148_in(8*N-1 downto 7*N),data2conv3 =>d148_in(7*N-1 downto 6*N),data2conv4 =>d148_in(6*N-1 downto 5*N),data2conv5 =>d148_in(5*N-1 downto 4*N),data2conv6 =>d148_in(4*N-1 downto 3*N),data2conv7 =>d148_in(3*N-1 downto 2*N),data2conv8 =>d148_in(2*N-1 downto N),data2conv9 =>d148_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d148_in(9*N-1 downto 8*N),w2 => d148_in(8*N-1 downto 7*N),w3 => d148_in(7*N-1 downto 6*N),w4 => d148_in(6*N-1 downto 5*N),w5 => d148_in(5*N-1 downto 4*N),w6 => d148_in(4*N-1 downto 3*N),w7 => d148_in(3*N-1 downto 2*N),w8 => d148_in(2*N-1 downto N),w9 => d148_in(N-1 downto 0 ),d_out => d148_out,en_out =>open  ,sof_out=>open   );
CL149: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d149_in(9*N-1 downto 8*N),data2conv2 =>d149_in(8*N-1 downto 7*N),data2conv3 =>d149_in(7*N-1 downto 6*N),data2conv4 =>d149_in(6*N-1 downto 5*N),data2conv5 =>d149_in(5*N-1 downto 4*N),data2conv6 =>d149_in(4*N-1 downto 3*N),data2conv7 =>d149_in(3*N-1 downto 2*N),data2conv8 =>d149_in(2*N-1 downto N),data2conv9 =>d149_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d149_in(9*N-1 downto 8*N),w2 => d149_in(8*N-1 downto 7*N),w3 => d149_in(7*N-1 downto 6*N),w4 => d149_in(6*N-1 downto 5*N),w5 => d149_in(5*N-1 downto 4*N),w6 => d149_in(4*N-1 downto 3*N),w7 => d149_in(3*N-1 downto 2*N),w8 => d149_in(2*N-1 downto N),w9 => d149_in(N-1 downto 0 ),d_out => d149_out,en_out =>open  ,sof_out=>open   );
CL150: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d150_in(9*N-1 downto 8*N),data2conv2 =>d150_in(8*N-1 downto 7*N),data2conv3 =>d150_in(7*N-1 downto 6*N),data2conv4 =>d150_in(6*N-1 downto 5*N),data2conv5 =>d150_in(5*N-1 downto 4*N),data2conv6 =>d150_in(4*N-1 downto 3*N),data2conv7 =>d150_in(3*N-1 downto 2*N),data2conv8 =>d150_in(2*N-1 downto N),data2conv9 =>d150_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d150_in(9*N-1 downto 8*N),w2 => d150_in(8*N-1 downto 7*N),w3 => d150_in(7*N-1 downto 6*N),w4 => d150_in(6*N-1 downto 5*N),w5 => d150_in(5*N-1 downto 4*N),w6 => d150_in(4*N-1 downto 3*N),w7 => d150_in(3*N-1 downto 2*N),w8 => d150_in(2*N-1 downto N),w9 => d150_in(N-1 downto 0 ),d_out => d150_out,en_out =>open  ,sof_out=>open   );
CL151: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d151_in(9*N-1 downto 8*N),data2conv2 =>d151_in(8*N-1 downto 7*N),data2conv3 =>d151_in(7*N-1 downto 6*N),data2conv4 =>d151_in(6*N-1 downto 5*N),data2conv5 =>d151_in(5*N-1 downto 4*N),data2conv6 =>d151_in(4*N-1 downto 3*N),data2conv7 =>d151_in(3*N-1 downto 2*N),data2conv8 =>d151_in(2*N-1 downto N),data2conv9 =>d151_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d151_in(9*N-1 downto 8*N),w2 => d151_in(8*N-1 downto 7*N),w3 => d151_in(7*N-1 downto 6*N),w4 => d151_in(6*N-1 downto 5*N),w5 => d151_in(5*N-1 downto 4*N),w6 => d151_in(4*N-1 downto 3*N),w7 => d151_in(3*N-1 downto 2*N),w8 => d151_in(2*N-1 downto N),w9 => d151_in(N-1 downto 0 ),d_out => d151_out,en_out =>open  ,sof_out=>open   );
CL152: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d152_in(9*N-1 downto 8*N),data2conv2 =>d152_in(8*N-1 downto 7*N),data2conv3 =>d152_in(7*N-1 downto 6*N),data2conv4 =>d152_in(6*N-1 downto 5*N),data2conv5 =>d152_in(5*N-1 downto 4*N),data2conv6 =>d152_in(4*N-1 downto 3*N),data2conv7 =>d152_in(3*N-1 downto 2*N),data2conv8 =>d152_in(2*N-1 downto N),data2conv9 =>d152_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d152_in(9*N-1 downto 8*N),w2 => d152_in(8*N-1 downto 7*N),w3 => d152_in(7*N-1 downto 6*N),w4 => d152_in(6*N-1 downto 5*N),w5 => d152_in(5*N-1 downto 4*N),w6 => d152_in(4*N-1 downto 3*N),w7 => d152_in(3*N-1 downto 2*N),w8 => d152_in(2*N-1 downto N),w9 => d152_in(N-1 downto 0 ),d_out => d152_out,en_out =>open  ,sof_out=>open   );
CL153: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d153_in(9*N-1 downto 8*N),data2conv2 =>d153_in(8*N-1 downto 7*N),data2conv3 =>d153_in(7*N-1 downto 6*N),data2conv4 =>d153_in(6*N-1 downto 5*N),data2conv5 =>d153_in(5*N-1 downto 4*N),data2conv6 =>d153_in(4*N-1 downto 3*N),data2conv7 =>d153_in(3*N-1 downto 2*N),data2conv8 =>d153_in(2*N-1 downto N),data2conv9 =>d153_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d153_in(9*N-1 downto 8*N),w2 => d153_in(8*N-1 downto 7*N),w3 => d153_in(7*N-1 downto 6*N),w4 => d153_in(6*N-1 downto 5*N),w5 => d153_in(5*N-1 downto 4*N),w6 => d153_in(4*N-1 downto 3*N),w7 => d153_in(3*N-1 downto 2*N),w8 => d153_in(2*N-1 downto N),w9 => d153_in(N-1 downto 0 ),d_out => d153_out,en_out =>open  ,sof_out=>open   );
CL154: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d154_in(9*N-1 downto 8*N),data2conv2 =>d154_in(8*N-1 downto 7*N),data2conv3 =>d154_in(7*N-1 downto 6*N),data2conv4 =>d154_in(6*N-1 downto 5*N),data2conv5 =>d154_in(5*N-1 downto 4*N),data2conv6 =>d154_in(4*N-1 downto 3*N),data2conv7 =>d154_in(3*N-1 downto 2*N),data2conv8 =>d154_in(2*N-1 downto N),data2conv9 =>d154_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d154_in(9*N-1 downto 8*N),w2 => d154_in(8*N-1 downto 7*N),w3 => d154_in(7*N-1 downto 6*N),w4 => d154_in(6*N-1 downto 5*N),w5 => d154_in(5*N-1 downto 4*N),w6 => d154_in(4*N-1 downto 3*N),w7 => d154_in(3*N-1 downto 2*N),w8 => d154_in(2*N-1 downto N),w9 => d154_in(N-1 downto 0 ),d_out => d154_out,en_out =>open  ,sof_out=>open   );
CL155: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d155_in(9*N-1 downto 8*N),data2conv2 =>d155_in(8*N-1 downto 7*N),data2conv3 =>d155_in(7*N-1 downto 6*N),data2conv4 =>d155_in(6*N-1 downto 5*N),data2conv5 =>d155_in(5*N-1 downto 4*N),data2conv6 =>d155_in(4*N-1 downto 3*N),data2conv7 =>d155_in(3*N-1 downto 2*N),data2conv8 =>d155_in(2*N-1 downto N),data2conv9 =>d155_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d155_in(9*N-1 downto 8*N),w2 => d155_in(8*N-1 downto 7*N),w3 => d155_in(7*N-1 downto 6*N),w4 => d155_in(6*N-1 downto 5*N),w5 => d155_in(5*N-1 downto 4*N),w6 => d155_in(4*N-1 downto 3*N),w7 => d155_in(3*N-1 downto 2*N),w8 => d155_in(2*N-1 downto N),w9 => d155_in(N-1 downto 0 ),d_out => d155_out,en_out =>open  ,sof_out=>open   );
CL156: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d156_in(9*N-1 downto 8*N),data2conv2 =>d156_in(8*N-1 downto 7*N),data2conv3 =>d156_in(7*N-1 downto 6*N),data2conv4 =>d156_in(6*N-1 downto 5*N),data2conv5 =>d156_in(5*N-1 downto 4*N),data2conv6 =>d156_in(4*N-1 downto 3*N),data2conv7 =>d156_in(3*N-1 downto 2*N),data2conv8 =>d156_in(2*N-1 downto N),data2conv9 =>d156_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d156_in(9*N-1 downto 8*N),w2 => d156_in(8*N-1 downto 7*N),w3 => d156_in(7*N-1 downto 6*N),w4 => d156_in(6*N-1 downto 5*N),w5 => d156_in(5*N-1 downto 4*N),w6 => d156_in(4*N-1 downto 3*N),w7 => d156_in(3*N-1 downto 2*N),w8 => d156_in(2*N-1 downto N),w9 => d156_in(N-1 downto 0 ),d_out => d156_out,en_out =>open  ,sof_out=>open   );
CL157: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d157_in(9*N-1 downto 8*N),data2conv2 =>d157_in(8*N-1 downto 7*N),data2conv3 =>d157_in(7*N-1 downto 6*N),data2conv4 =>d157_in(6*N-1 downto 5*N),data2conv5 =>d157_in(5*N-1 downto 4*N),data2conv6 =>d157_in(4*N-1 downto 3*N),data2conv7 =>d157_in(3*N-1 downto 2*N),data2conv8 =>d157_in(2*N-1 downto N),data2conv9 =>d157_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d157_in(9*N-1 downto 8*N),w2 => d157_in(8*N-1 downto 7*N),w3 => d157_in(7*N-1 downto 6*N),w4 => d157_in(6*N-1 downto 5*N),w5 => d157_in(5*N-1 downto 4*N),w6 => d157_in(4*N-1 downto 3*N),w7 => d157_in(3*N-1 downto 2*N),w8 => d157_in(2*N-1 downto N),w9 => d157_in(N-1 downto 0 ),d_out => d157_out,en_out =>open  ,sof_out=>open   );
CL158: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d158_in(9*N-1 downto 8*N),data2conv2 =>d158_in(8*N-1 downto 7*N),data2conv3 =>d158_in(7*N-1 downto 6*N),data2conv4 =>d158_in(6*N-1 downto 5*N),data2conv5 =>d158_in(5*N-1 downto 4*N),data2conv6 =>d158_in(4*N-1 downto 3*N),data2conv7 =>d158_in(3*N-1 downto 2*N),data2conv8 =>d158_in(2*N-1 downto N),data2conv9 =>d158_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d158_in(9*N-1 downto 8*N),w2 => d158_in(8*N-1 downto 7*N),w3 => d158_in(7*N-1 downto 6*N),w4 => d158_in(6*N-1 downto 5*N),w5 => d158_in(5*N-1 downto 4*N),w6 => d158_in(4*N-1 downto 3*N),w7 => d158_in(3*N-1 downto 2*N),w8 => d158_in(2*N-1 downto N),w9 => d158_in(N-1 downto 0 ),d_out => d158_out,en_out =>open  ,sof_out=>open   );
CL159: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d159_in(9*N-1 downto 8*N),data2conv2 =>d159_in(8*N-1 downto 7*N),data2conv3 =>d159_in(7*N-1 downto 6*N),data2conv4 =>d159_in(6*N-1 downto 5*N),data2conv5 =>d159_in(5*N-1 downto 4*N),data2conv6 =>d159_in(4*N-1 downto 3*N),data2conv7 =>d159_in(3*N-1 downto 2*N),data2conv8 =>d159_in(2*N-1 downto N),data2conv9 =>d159_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d159_in(9*N-1 downto 8*N),w2 => d159_in(8*N-1 downto 7*N),w3 => d159_in(7*N-1 downto 6*N),w4 => d159_in(6*N-1 downto 5*N),w5 => d159_in(5*N-1 downto 4*N),w6 => d159_in(4*N-1 downto 3*N),w7 => d159_in(3*N-1 downto 2*N),w8 => d159_in(2*N-1 downto N),w9 => d159_in(N-1 downto 0 ),d_out => d159_out,en_out =>open  ,sof_out=>open   );
CL160: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d160_in(9*N-1 downto 8*N),data2conv2 =>d160_in(8*N-1 downto 7*N),data2conv3 =>d160_in(7*N-1 downto 6*N),data2conv4 =>d160_in(6*N-1 downto 5*N),data2conv5 =>d160_in(5*N-1 downto 4*N),data2conv6 =>d160_in(4*N-1 downto 3*N),data2conv7 =>d160_in(3*N-1 downto 2*N),data2conv8 =>d160_in(2*N-1 downto N),data2conv9 =>d160_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d160_in(9*N-1 downto 8*N),w2 => d160_in(8*N-1 downto 7*N),w3 => d160_in(7*N-1 downto 6*N),w4 => d160_in(6*N-1 downto 5*N),w5 => d160_in(5*N-1 downto 4*N),w6 => d160_in(4*N-1 downto 3*N),w7 => d160_in(3*N-1 downto 2*N),w8 => d160_in(2*N-1 downto N),w9 => d160_in(N-1 downto 0 ),d_out => d160_out,en_out =>open  ,sof_out=>open   );
CL161: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d161_in(9*N-1 downto 8*N),data2conv2 =>d161_in(8*N-1 downto 7*N),data2conv3 =>d161_in(7*N-1 downto 6*N),data2conv4 =>d161_in(6*N-1 downto 5*N),data2conv5 =>d161_in(5*N-1 downto 4*N),data2conv6 =>d161_in(4*N-1 downto 3*N),data2conv7 =>d161_in(3*N-1 downto 2*N),data2conv8 =>d161_in(2*N-1 downto N),data2conv9 =>d161_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d161_in(9*N-1 downto 8*N),w2 => d161_in(8*N-1 downto 7*N),w3 => d161_in(7*N-1 downto 6*N),w4 => d161_in(6*N-1 downto 5*N),w5 => d161_in(5*N-1 downto 4*N),w6 => d161_in(4*N-1 downto 3*N),w7 => d161_in(3*N-1 downto 2*N),w8 => d161_in(2*N-1 downto N),w9 => d161_in(N-1 downto 0 ),d_out => d161_out,en_out =>open  ,sof_out=>open   );
CL162: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d162_in(9*N-1 downto 8*N),data2conv2 =>d162_in(8*N-1 downto 7*N),data2conv3 =>d162_in(7*N-1 downto 6*N),data2conv4 =>d162_in(6*N-1 downto 5*N),data2conv5 =>d162_in(5*N-1 downto 4*N),data2conv6 =>d162_in(4*N-1 downto 3*N),data2conv7 =>d162_in(3*N-1 downto 2*N),data2conv8 =>d162_in(2*N-1 downto N),data2conv9 =>d162_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d162_in(9*N-1 downto 8*N),w2 => d162_in(8*N-1 downto 7*N),w3 => d162_in(7*N-1 downto 6*N),w4 => d162_in(6*N-1 downto 5*N),w5 => d162_in(5*N-1 downto 4*N),w6 => d162_in(4*N-1 downto 3*N),w7 => d162_in(3*N-1 downto 2*N),w8 => d162_in(2*N-1 downto N),w9 => d162_in(N-1 downto 0 ),d_out => d162_out,en_out =>open  ,sof_out=>open   );
CL163: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d163_in(9*N-1 downto 8*N),data2conv2 =>d163_in(8*N-1 downto 7*N),data2conv3 =>d163_in(7*N-1 downto 6*N),data2conv4 =>d163_in(6*N-1 downto 5*N),data2conv5 =>d163_in(5*N-1 downto 4*N),data2conv6 =>d163_in(4*N-1 downto 3*N),data2conv7 =>d163_in(3*N-1 downto 2*N),data2conv8 =>d163_in(2*N-1 downto N),data2conv9 =>d163_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d163_in(9*N-1 downto 8*N),w2 => d163_in(8*N-1 downto 7*N),w3 => d163_in(7*N-1 downto 6*N),w4 => d163_in(6*N-1 downto 5*N),w5 => d163_in(5*N-1 downto 4*N),w6 => d163_in(4*N-1 downto 3*N),w7 => d163_in(3*N-1 downto 2*N),w8 => d163_in(2*N-1 downto N),w9 => d163_in(N-1 downto 0 ),d_out => d163_out,en_out =>open  ,sof_out=>open   );
CL164: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d164_in(9*N-1 downto 8*N),data2conv2 =>d164_in(8*N-1 downto 7*N),data2conv3 =>d164_in(7*N-1 downto 6*N),data2conv4 =>d164_in(6*N-1 downto 5*N),data2conv5 =>d164_in(5*N-1 downto 4*N),data2conv6 =>d164_in(4*N-1 downto 3*N),data2conv7 =>d164_in(3*N-1 downto 2*N),data2conv8 =>d164_in(2*N-1 downto N),data2conv9 =>d164_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d164_in(9*N-1 downto 8*N),w2 => d164_in(8*N-1 downto 7*N),w3 => d164_in(7*N-1 downto 6*N),w4 => d164_in(6*N-1 downto 5*N),w5 => d164_in(5*N-1 downto 4*N),w6 => d164_in(4*N-1 downto 3*N),w7 => d164_in(3*N-1 downto 2*N),w8 => d164_in(2*N-1 downto N),w9 => d164_in(N-1 downto 0 ),d_out => d164_out,en_out =>open  ,sof_out=>open   );
CL165: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d165_in(9*N-1 downto 8*N),data2conv2 =>d165_in(8*N-1 downto 7*N),data2conv3 =>d165_in(7*N-1 downto 6*N),data2conv4 =>d165_in(6*N-1 downto 5*N),data2conv5 =>d165_in(5*N-1 downto 4*N),data2conv6 =>d165_in(4*N-1 downto 3*N),data2conv7 =>d165_in(3*N-1 downto 2*N),data2conv8 =>d165_in(2*N-1 downto N),data2conv9 =>d165_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d165_in(9*N-1 downto 8*N),w2 => d165_in(8*N-1 downto 7*N),w3 => d165_in(7*N-1 downto 6*N),w4 => d165_in(6*N-1 downto 5*N),w5 => d165_in(5*N-1 downto 4*N),w6 => d165_in(4*N-1 downto 3*N),w7 => d165_in(3*N-1 downto 2*N),w8 => d165_in(2*N-1 downto N),w9 => d165_in(N-1 downto 0 ),d_out => d165_out,en_out =>open  ,sof_out=>open   );
CL166: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d166_in(9*N-1 downto 8*N),data2conv2 =>d166_in(8*N-1 downto 7*N),data2conv3 =>d166_in(7*N-1 downto 6*N),data2conv4 =>d166_in(6*N-1 downto 5*N),data2conv5 =>d166_in(5*N-1 downto 4*N),data2conv6 =>d166_in(4*N-1 downto 3*N),data2conv7 =>d166_in(3*N-1 downto 2*N),data2conv8 =>d166_in(2*N-1 downto N),data2conv9 =>d166_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d166_in(9*N-1 downto 8*N),w2 => d166_in(8*N-1 downto 7*N),w3 => d166_in(7*N-1 downto 6*N),w4 => d166_in(6*N-1 downto 5*N),w5 => d166_in(5*N-1 downto 4*N),w6 => d166_in(4*N-1 downto 3*N),w7 => d166_in(3*N-1 downto 2*N),w8 => d166_in(2*N-1 downto N),w9 => d166_in(N-1 downto 0 ),d_out => d166_out,en_out =>open  ,sof_out=>open   );
CL167: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d167_in(9*N-1 downto 8*N),data2conv2 =>d167_in(8*N-1 downto 7*N),data2conv3 =>d167_in(7*N-1 downto 6*N),data2conv4 =>d167_in(6*N-1 downto 5*N),data2conv5 =>d167_in(5*N-1 downto 4*N),data2conv6 =>d167_in(4*N-1 downto 3*N),data2conv7 =>d167_in(3*N-1 downto 2*N),data2conv8 =>d167_in(2*N-1 downto N),data2conv9 =>d167_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d167_in(9*N-1 downto 8*N),w2 => d167_in(8*N-1 downto 7*N),w3 => d167_in(7*N-1 downto 6*N),w4 => d167_in(6*N-1 downto 5*N),w5 => d167_in(5*N-1 downto 4*N),w6 => d167_in(4*N-1 downto 3*N),w7 => d167_in(3*N-1 downto 2*N),w8 => d167_in(2*N-1 downto N),w9 => d167_in(N-1 downto 0 ),d_out => d167_out,en_out =>open  ,sof_out=>open   );
CL168: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d168_in(9*N-1 downto 8*N),data2conv2 =>d168_in(8*N-1 downto 7*N),data2conv3 =>d168_in(7*N-1 downto 6*N),data2conv4 =>d168_in(6*N-1 downto 5*N),data2conv5 =>d168_in(5*N-1 downto 4*N),data2conv6 =>d168_in(4*N-1 downto 3*N),data2conv7 =>d168_in(3*N-1 downto 2*N),data2conv8 =>d168_in(2*N-1 downto N),data2conv9 =>d168_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d168_in(9*N-1 downto 8*N),w2 => d168_in(8*N-1 downto 7*N),w3 => d168_in(7*N-1 downto 6*N),w4 => d168_in(6*N-1 downto 5*N),w5 => d168_in(5*N-1 downto 4*N),w6 => d168_in(4*N-1 downto 3*N),w7 => d168_in(3*N-1 downto 2*N),w8 => d168_in(2*N-1 downto N),w9 => d168_in(N-1 downto 0 ),d_out => d168_out,en_out =>open  ,sof_out=>open   );
CL169: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d169_in(9*N-1 downto 8*N),data2conv2 =>d169_in(8*N-1 downto 7*N),data2conv3 =>d169_in(7*N-1 downto 6*N),data2conv4 =>d169_in(6*N-1 downto 5*N),data2conv5 =>d169_in(5*N-1 downto 4*N),data2conv6 =>d169_in(4*N-1 downto 3*N),data2conv7 =>d169_in(3*N-1 downto 2*N),data2conv8 =>d169_in(2*N-1 downto N),data2conv9 =>d169_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d169_in(9*N-1 downto 8*N),w2 => d169_in(8*N-1 downto 7*N),w3 => d169_in(7*N-1 downto 6*N),w4 => d169_in(6*N-1 downto 5*N),w5 => d169_in(5*N-1 downto 4*N),w6 => d169_in(4*N-1 downto 3*N),w7 => d169_in(3*N-1 downto 2*N),w8 => d169_in(2*N-1 downto N),w9 => d169_in(N-1 downto 0 ),d_out => d169_out,en_out =>open  ,sof_out=>open   );
CL170: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d170_in(9*N-1 downto 8*N),data2conv2 =>d170_in(8*N-1 downto 7*N),data2conv3 =>d170_in(7*N-1 downto 6*N),data2conv4 =>d170_in(6*N-1 downto 5*N),data2conv5 =>d170_in(5*N-1 downto 4*N),data2conv6 =>d170_in(4*N-1 downto 3*N),data2conv7 =>d170_in(3*N-1 downto 2*N),data2conv8 =>d170_in(2*N-1 downto N),data2conv9 =>d170_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d170_in(9*N-1 downto 8*N),w2 => d170_in(8*N-1 downto 7*N),w3 => d170_in(7*N-1 downto 6*N),w4 => d170_in(6*N-1 downto 5*N),w5 => d170_in(5*N-1 downto 4*N),w6 => d170_in(4*N-1 downto 3*N),w7 => d170_in(3*N-1 downto 2*N),w8 => d170_in(2*N-1 downto N),w9 => d170_in(N-1 downto 0 ),d_out => d170_out,en_out =>open  ,sof_out=>open   );
CL171: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d171_in(9*N-1 downto 8*N),data2conv2 =>d171_in(8*N-1 downto 7*N),data2conv3 =>d171_in(7*N-1 downto 6*N),data2conv4 =>d171_in(6*N-1 downto 5*N),data2conv5 =>d171_in(5*N-1 downto 4*N),data2conv6 =>d171_in(4*N-1 downto 3*N),data2conv7 =>d171_in(3*N-1 downto 2*N),data2conv8 =>d171_in(2*N-1 downto N),data2conv9 =>d171_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d171_in(9*N-1 downto 8*N),w2 => d171_in(8*N-1 downto 7*N),w3 => d171_in(7*N-1 downto 6*N),w4 => d171_in(6*N-1 downto 5*N),w5 => d171_in(5*N-1 downto 4*N),w6 => d171_in(4*N-1 downto 3*N),w7 => d171_in(3*N-1 downto 2*N),w8 => d171_in(2*N-1 downto N),w9 => d171_in(N-1 downto 0 ),d_out => d171_out,en_out =>open  ,sof_out=>open   );
CL172: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d172_in(9*N-1 downto 8*N),data2conv2 =>d172_in(8*N-1 downto 7*N),data2conv3 =>d172_in(7*N-1 downto 6*N),data2conv4 =>d172_in(6*N-1 downto 5*N),data2conv5 =>d172_in(5*N-1 downto 4*N),data2conv6 =>d172_in(4*N-1 downto 3*N),data2conv7 =>d172_in(3*N-1 downto 2*N),data2conv8 =>d172_in(2*N-1 downto N),data2conv9 =>d172_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d172_in(9*N-1 downto 8*N),w2 => d172_in(8*N-1 downto 7*N),w3 => d172_in(7*N-1 downto 6*N),w4 => d172_in(6*N-1 downto 5*N),w5 => d172_in(5*N-1 downto 4*N),w6 => d172_in(4*N-1 downto 3*N),w7 => d172_in(3*N-1 downto 2*N),w8 => d172_in(2*N-1 downto N),w9 => d172_in(N-1 downto 0 ),d_out => d172_out,en_out =>open  ,sof_out=>open   );
CL173: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d173_in(9*N-1 downto 8*N),data2conv2 =>d173_in(8*N-1 downto 7*N),data2conv3 =>d173_in(7*N-1 downto 6*N),data2conv4 =>d173_in(6*N-1 downto 5*N),data2conv5 =>d173_in(5*N-1 downto 4*N),data2conv6 =>d173_in(4*N-1 downto 3*N),data2conv7 =>d173_in(3*N-1 downto 2*N),data2conv8 =>d173_in(2*N-1 downto N),data2conv9 =>d173_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d173_in(9*N-1 downto 8*N),w2 => d173_in(8*N-1 downto 7*N),w3 => d173_in(7*N-1 downto 6*N),w4 => d173_in(6*N-1 downto 5*N),w5 => d173_in(5*N-1 downto 4*N),w6 => d173_in(4*N-1 downto 3*N),w7 => d173_in(3*N-1 downto 2*N),w8 => d173_in(2*N-1 downto N),w9 => d173_in(N-1 downto 0 ),d_out => d173_out,en_out =>open  ,sof_out=>open   );
CL174: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d174_in(9*N-1 downto 8*N),data2conv2 =>d174_in(8*N-1 downto 7*N),data2conv3 =>d174_in(7*N-1 downto 6*N),data2conv4 =>d174_in(6*N-1 downto 5*N),data2conv5 =>d174_in(5*N-1 downto 4*N),data2conv6 =>d174_in(4*N-1 downto 3*N),data2conv7 =>d174_in(3*N-1 downto 2*N),data2conv8 =>d174_in(2*N-1 downto N),data2conv9 =>d174_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d174_in(9*N-1 downto 8*N),w2 => d174_in(8*N-1 downto 7*N),w3 => d174_in(7*N-1 downto 6*N),w4 => d174_in(6*N-1 downto 5*N),w5 => d174_in(5*N-1 downto 4*N),w6 => d174_in(4*N-1 downto 3*N),w7 => d174_in(3*N-1 downto 2*N),w8 => d174_in(2*N-1 downto N),w9 => d174_in(N-1 downto 0 ),d_out => d174_out,en_out =>open  ,sof_out=>open   );
CL175: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d175_in(9*N-1 downto 8*N),data2conv2 =>d175_in(8*N-1 downto 7*N),data2conv3 =>d175_in(7*N-1 downto 6*N),data2conv4 =>d175_in(6*N-1 downto 5*N),data2conv5 =>d175_in(5*N-1 downto 4*N),data2conv6 =>d175_in(4*N-1 downto 3*N),data2conv7 =>d175_in(3*N-1 downto 2*N),data2conv8 =>d175_in(2*N-1 downto N),data2conv9 =>d175_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d175_in(9*N-1 downto 8*N),w2 => d175_in(8*N-1 downto 7*N),w3 => d175_in(7*N-1 downto 6*N),w4 => d175_in(6*N-1 downto 5*N),w5 => d175_in(5*N-1 downto 4*N),w6 => d175_in(4*N-1 downto 3*N),w7 => d175_in(3*N-1 downto 2*N),w8 => d175_in(2*N-1 downto N),w9 => d175_in(N-1 downto 0 ),d_out => d175_out,en_out =>open  ,sof_out=>open   );
CL176: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d176_in(9*N-1 downto 8*N),data2conv2 =>d176_in(8*N-1 downto 7*N),data2conv3 =>d176_in(7*N-1 downto 6*N),data2conv4 =>d176_in(6*N-1 downto 5*N),data2conv5 =>d176_in(5*N-1 downto 4*N),data2conv6 =>d176_in(4*N-1 downto 3*N),data2conv7 =>d176_in(3*N-1 downto 2*N),data2conv8 =>d176_in(2*N-1 downto N),data2conv9 =>d176_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d176_in(9*N-1 downto 8*N),w2 => d176_in(8*N-1 downto 7*N),w3 => d176_in(7*N-1 downto 6*N),w4 => d176_in(6*N-1 downto 5*N),w5 => d176_in(5*N-1 downto 4*N),w6 => d176_in(4*N-1 downto 3*N),w7 => d176_in(3*N-1 downto 2*N),w8 => d176_in(2*N-1 downto N),w9 => d176_in(N-1 downto 0 ),d_out => d176_out,en_out =>open  ,sof_out=>open   );
CL177: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d177_in(9*N-1 downto 8*N),data2conv2 =>d177_in(8*N-1 downto 7*N),data2conv3 =>d177_in(7*N-1 downto 6*N),data2conv4 =>d177_in(6*N-1 downto 5*N),data2conv5 =>d177_in(5*N-1 downto 4*N),data2conv6 =>d177_in(4*N-1 downto 3*N),data2conv7 =>d177_in(3*N-1 downto 2*N),data2conv8 =>d177_in(2*N-1 downto N),data2conv9 =>d177_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d177_in(9*N-1 downto 8*N),w2 => d177_in(8*N-1 downto 7*N),w3 => d177_in(7*N-1 downto 6*N),w4 => d177_in(6*N-1 downto 5*N),w5 => d177_in(5*N-1 downto 4*N),w6 => d177_in(4*N-1 downto 3*N),w7 => d177_in(3*N-1 downto 2*N),w8 => d177_in(2*N-1 downto N),w9 => d177_in(N-1 downto 0 ),d_out => d177_out,en_out =>open  ,sof_out=>open   );
CL178: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d178_in(9*N-1 downto 8*N),data2conv2 =>d178_in(8*N-1 downto 7*N),data2conv3 =>d178_in(7*N-1 downto 6*N),data2conv4 =>d178_in(6*N-1 downto 5*N),data2conv5 =>d178_in(5*N-1 downto 4*N),data2conv6 =>d178_in(4*N-1 downto 3*N),data2conv7 =>d178_in(3*N-1 downto 2*N),data2conv8 =>d178_in(2*N-1 downto N),data2conv9 =>d178_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d178_in(9*N-1 downto 8*N),w2 => d178_in(8*N-1 downto 7*N),w3 => d178_in(7*N-1 downto 6*N),w4 => d178_in(6*N-1 downto 5*N),w5 => d178_in(5*N-1 downto 4*N),w6 => d178_in(4*N-1 downto 3*N),w7 => d178_in(3*N-1 downto 2*N),w8 => d178_in(2*N-1 downto N),w9 => d178_in(N-1 downto 0 ),d_out => d178_out,en_out =>open  ,sof_out=>open   );
CL179: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d179_in(9*N-1 downto 8*N),data2conv2 =>d179_in(8*N-1 downto 7*N),data2conv3 =>d179_in(7*N-1 downto 6*N),data2conv4 =>d179_in(6*N-1 downto 5*N),data2conv5 =>d179_in(5*N-1 downto 4*N),data2conv6 =>d179_in(4*N-1 downto 3*N),data2conv7 =>d179_in(3*N-1 downto 2*N),data2conv8 =>d179_in(2*N-1 downto N),data2conv9 =>d179_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d179_in(9*N-1 downto 8*N),w2 => d179_in(8*N-1 downto 7*N),w3 => d179_in(7*N-1 downto 6*N),w4 => d179_in(6*N-1 downto 5*N),w5 => d179_in(5*N-1 downto 4*N),w6 => d179_in(4*N-1 downto 3*N),w7 => d179_in(3*N-1 downto 2*N),w8 => d179_in(2*N-1 downto N),w9 => d179_in(N-1 downto 0 ),d_out => d179_out,en_out =>open  ,sof_out=>open   );
CL180: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d180_in(9*N-1 downto 8*N),data2conv2 =>d180_in(8*N-1 downto 7*N),data2conv3 =>d180_in(7*N-1 downto 6*N),data2conv4 =>d180_in(6*N-1 downto 5*N),data2conv5 =>d180_in(5*N-1 downto 4*N),data2conv6 =>d180_in(4*N-1 downto 3*N),data2conv7 =>d180_in(3*N-1 downto 2*N),data2conv8 =>d180_in(2*N-1 downto N),data2conv9 =>d180_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d180_in(9*N-1 downto 8*N),w2 => d180_in(8*N-1 downto 7*N),w3 => d180_in(7*N-1 downto 6*N),w4 => d180_in(6*N-1 downto 5*N),w5 => d180_in(5*N-1 downto 4*N),w6 => d180_in(4*N-1 downto 3*N),w7 => d180_in(3*N-1 downto 2*N),w8 => d180_in(2*N-1 downto N),w9 => d180_in(N-1 downto 0 ),d_out => d180_out,en_out =>open  ,sof_out=>open   );
CL181: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d181_in(9*N-1 downto 8*N),data2conv2 =>d181_in(8*N-1 downto 7*N),data2conv3 =>d181_in(7*N-1 downto 6*N),data2conv4 =>d181_in(6*N-1 downto 5*N),data2conv5 =>d181_in(5*N-1 downto 4*N),data2conv6 =>d181_in(4*N-1 downto 3*N),data2conv7 =>d181_in(3*N-1 downto 2*N),data2conv8 =>d181_in(2*N-1 downto N),data2conv9 =>d181_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d181_in(9*N-1 downto 8*N),w2 => d181_in(8*N-1 downto 7*N),w3 => d181_in(7*N-1 downto 6*N),w4 => d181_in(6*N-1 downto 5*N),w5 => d181_in(5*N-1 downto 4*N),w6 => d181_in(4*N-1 downto 3*N),w7 => d181_in(3*N-1 downto 2*N),w8 => d181_in(2*N-1 downto N),w9 => d181_in(N-1 downto 0 ),d_out => d181_out,en_out =>open  ,sof_out=>open   );
CL182: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d182_in(9*N-1 downto 8*N),data2conv2 =>d182_in(8*N-1 downto 7*N),data2conv3 =>d182_in(7*N-1 downto 6*N),data2conv4 =>d182_in(6*N-1 downto 5*N),data2conv5 =>d182_in(5*N-1 downto 4*N),data2conv6 =>d182_in(4*N-1 downto 3*N),data2conv7 =>d182_in(3*N-1 downto 2*N),data2conv8 =>d182_in(2*N-1 downto N),data2conv9 =>d182_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d182_in(9*N-1 downto 8*N),w2 => d182_in(8*N-1 downto 7*N),w3 => d182_in(7*N-1 downto 6*N),w4 => d182_in(6*N-1 downto 5*N),w5 => d182_in(5*N-1 downto 4*N),w6 => d182_in(4*N-1 downto 3*N),w7 => d182_in(3*N-1 downto 2*N),w8 => d182_in(2*N-1 downto N),w9 => d182_in(N-1 downto 0 ),d_out => d182_out,en_out =>open  ,sof_out=>open   );
CL183: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d183_in(9*N-1 downto 8*N),data2conv2 =>d183_in(8*N-1 downto 7*N),data2conv3 =>d183_in(7*N-1 downto 6*N),data2conv4 =>d183_in(6*N-1 downto 5*N),data2conv5 =>d183_in(5*N-1 downto 4*N),data2conv6 =>d183_in(4*N-1 downto 3*N),data2conv7 =>d183_in(3*N-1 downto 2*N),data2conv8 =>d183_in(2*N-1 downto N),data2conv9 =>d183_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d183_in(9*N-1 downto 8*N),w2 => d183_in(8*N-1 downto 7*N),w3 => d183_in(7*N-1 downto 6*N),w4 => d183_in(6*N-1 downto 5*N),w5 => d183_in(5*N-1 downto 4*N),w6 => d183_in(4*N-1 downto 3*N),w7 => d183_in(3*N-1 downto 2*N),w8 => d183_in(2*N-1 downto N),w9 => d183_in(N-1 downto 0 ),d_out => d183_out,en_out =>open  ,sof_out=>open   );
CL184: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d184_in(9*N-1 downto 8*N),data2conv2 =>d184_in(8*N-1 downto 7*N),data2conv3 =>d184_in(7*N-1 downto 6*N),data2conv4 =>d184_in(6*N-1 downto 5*N),data2conv5 =>d184_in(5*N-1 downto 4*N),data2conv6 =>d184_in(4*N-1 downto 3*N),data2conv7 =>d184_in(3*N-1 downto 2*N),data2conv8 =>d184_in(2*N-1 downto N),data2conv9 =>d184_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d184_in(9*N-1 downto 8*N),w2 => d184_in(8*N-1 downto 7*N),w3 => d184_in(7*N-1 downto 6*N),w4 => d184_in(6*N-1 downto 5*N),w5 => d184_in(5*N-1 downto 4*N),w6 => d184_in(4*N-1 downto 3*N),w7 => d184_in(3*N-1 downto 2*N),w8 => d184_in(2*N-1 downto N),w9 => d184_in(N-1 downto 0 ),d_out => d184_out,en_out =>open  ,sof_out=>open   );
CL185: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d185_in(9*N-1 downto 8*N),data2conv2 =>d185_in(8*N-1 downto 7*N),data2conv3 =>d185_in(7*N-1 downto 6*N),data2conv4 =>d185_in(6*N-1 downto 5*N),data2conv5 =>d185_in(5*N-1 downto 4*N),data2conv6 =>d185_in(4*N-1 downto 3*N),data2conv7 =>d185_in(3*N-1 downto 2*N),data2conv8 =>d185_in(2*N-1 downto N),data2conv9 =>d185_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d185_in(9*N-1 downto 8*N),w2 => d185_in(8*N-1 downto 7*N),w3 => d185_in(7*N-1 downto 6*N),w4 => d185_in(6*N-1 downto 5*N),w5 => d185_in(5*N-1 downto 4*N),w6 => d185_in(4*N-1 downto 3*N),w7 => d185_in(3*N-1 downto 2*N),w8 => d185_in(2*N-1 downto N),w9 => d185_in(N-1 downto 0 ),d_out => d185_out,en_out =>open  ,sof_out=>open   );
CL186: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d186_in(9*N-1 downto 8*N),data2conv2 =>d186_in(8*N-1 downto 7*N),data2conv3 =>d186_in(7*N-1 downto 6*N),data2conv4 =>d186_in(6*N-1 downto 5*N),data2conv5 =>d186_in(5*N-1 downto 4*N),data2conv6 =>d186_in(4*N-1 downto 3*N),data2conv7 =>d186_in(3*N-1 downto 2*N),data2conv8 =>d186_in(2*N-1 downto N),data2conv9 =>d186_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d186_in(9*N-1 downto 8*N),w2 => d186_in(8*N-1 downto 7*N),w3 => d186_in(7*N-1 downto 6*N),w4 => d186_in(6*N-1 downto 5*N),w5 => d186_in(5*N-1 downto 4*N),w6 => d186_in(4*N-1 downto 3*N),w7 => d186_in(3*N-1 downto 2*N),w8 => d186_in(2*N-1 downto N),w9 => d186_in(N-1 downto 0 ),d_out => d186_out,en_out =>open  ,sof_out=>open   );
CL187: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d187_in(9*N-1 downto 8*N),data2conv2 =>d187_in(8*N-1 downto 7*N),data2conv3 =>d187_in(7*N-1 downto 6*N),data2conv4 =>d187_in(6*N-1 downto 5*N),data2conv5 =>d187_in(5*N-1 downto 4*N),data2conv6 =>d187_in(4*N-1 downto 3*N),data2conv7 =>d187_in(3*N-1 downto 2*N),data2conv8 =>d187_in(2*N-1 downto N),data2conv9 =>d187_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d187_in(9*N-1 downto 8*N),w2 => d187_in(8*N-1 downto 7*N),w3 => d187_in(7*N-1 downto 6*N),w4 => d187_in(6*N-1 downto 5*N),w5 => d187_in(5*N-1 downto 4*N),w6 => d187_in(4*N-1 downto 3*N),w7 => d187_in(3*N-1 downto 2*N),w8 => d187_in(2*N-1 downto N),w9 => d187_in(N-1 downto 0 ),d_out => d187_out,en_out =>open  ,sof_out=>open   );
CL188: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d188_in(9*N-1 downto 8*N),data2conv2 =>d188_in(8*N-1 downto 7*N),data2conv3 =>d188_in(7*N-1 downto 6*N),data2conv4 =>d188_in(6*N-1 downto 5*N),data2conv5 =>d188_in(5*N-1 downto 4*N),data2conv6 =>d188_in(4*N-1 downto 3*N),data2conv7 =>d188_in(3*N-1 downto 2*N),data2conv8 =>d188_in(2*N-1 downto N),data2conv9 =>d188_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d188_in(9*N-1 downto 8*N),w2 => d188_in(8*N-1 downto 7*N),w3 => d188_in(7*N-1 downto 6*N),w4 => d188_in(6*N-1 downto 5*N),w5 => d188_in(5*N-1 downto 4*N),w6 => d188_in(4*N-1 downto 3*N),w7 => d188_in(3*N-1 downto 2*N),w8 => d188_in(2*N-1 downto N),w9 => d188_in(N-1 downto 0 ),d_out => d188_out,en_out =>open  ,sof_out=>open   );
CL189: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d189_in(9*N-1 downto 8*N),data2conv2 =>d189_in(8*N-1 downto 7*N),data2conv3 =>d189_in(7*N-1 downto 6*N),data2conv4 =>d189_in(6*N-1 downto 5*N),data2conv5 =>d189_in(5*N-1 downto 4*N),data2conv6 =>d189_in(4*N-1 downto 3*N),data2conv7 =>d189_in(3*N-1 downto 2*N),data2conv8 =>d189_in(2*N-1 downto N),data2conv9 =>d189_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d189_in(9*N-1 downto 8*N),w2 => d189_in(8*N-1 downto 7*N),w3 => d189_in(7*N-1 downto 6*N),w4 => d189_in(6*N-1 downto 5*N),w5 => d189_in(5*N-1 downto 4*N),w6 => d189_in(4*N-1 downto 3*N),w7 => d189_in(3*N-1 downto 2*N),w8 => d189_in(2*N-1 downto N),w9 => d189_in(N-1 downto 0 ),d_out => d189_out,en_out =>open  ,sof_out=>open   );
CL190: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d190_in(9*N-1 downto 8*N),data2conv2 =>d190_in(8*N-1 downto 7*N),data2conv3 =>d190_in(7*N-1 downto 6*N),data2conv4 =>d190_in(6*N-1 downto 5*N),data2conv5 =>d190_in(5*N-1 downto 4*N),data2conv6 =>d190_in(4*N-1 downto 3*N),data2conv7 =>d190_in(3*N-1 downto 2*N),data2conv8 =>d190_in(2*N-1 downto N),data2conv9 =>d190_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d190_in(9*N-1 downto 8*N),w2 => d190_in(8*N-1 downto 7*N),w3 => d190_in(7*N-1 downto 6*N),w4 => d190_in(6*N-1 downto 5*N),w5 => d190_in(5*N-1 downto 4*N),w6 => d190_in(4*N-1 downto 3*N),w7 => d190_in(3*N-1 downto 2*N),w8 => d190_in(2*N-1 downto N),w9 => d190_in(N-1 downto 0 ),d_out => d190_out,en_out =>open  ,sof_out=>open   );
CL191: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d191_in(9*N-1 downto 8*N),data2conv2 =>d191_in(8*N-1 downto 7*N),data2conv3 =>d191_in(7*N-1 downto 6*N),data2conv4 =>d191_in(6*N-1 downto 5*N),data2conv5 =>d191_in(5*N-1 downto 4*N),data2conv6 =>d191_in(4*N-1 downto 3*N),data2conv7 =>d191_in(3*N-1 downto 2*N),data2conv8 =>d191_in(2*N-1 downto N),data2conv9 =>d191_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d191_in(9*N-1 downto 8*N),w2 => d191_in(8*N-1 downto 7*N),w3 => d191_in(7*N-1 downto 6*N),w4 => d191_in(6*N-1 downto 5*N),w5 => d191_in(5*N-1 downto 4*N),w6 => d191_in(4*N-1 downto 3*N),w7 => d191_in(3*N-1 downto 2*N),w8 => d191_in(2*N-1 downto N),w9 => d191_in(N-1 downto 0 ),d_out => d191_out,en_out =>open  ,sof_out=>open   );
CL192: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d192_in(9*N-1 downto 8*N),data2conv2 =>d192_in(8*N-1 downto 7*N),data2conv3 =>d192_in(7*N-1 downto 6*N),data2conv4 =>d192_in(6*N-1 downto 5*N),data2conv5 =>d192_in(5*N-1 downto 4*N),data2conv6 =>d192_in(4*N-1 downto 3*N),data2conv7 =>d192_in(3*N-1 downto 2*N),data2conv8 =>d192_in(2*N-1 downto N),data2conv9 =>d192_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d192_in(9*N-1 downto 8*N),w2 => d192_in(8*N-1 downto 7*N),w3 => d192_in(7*N-1 downto 6*N),w4 => d192_in(6*N-1 downto 5*N),w5 => d192_in(5*N-1 downto 4*N),w6 => d192_in(4*N-1 downto 3*N),w7 => d192_in(3*N-1 downto 2*N),w8 => d192_in(2*N-1 downto N),w9 => d192_in(N-1 downto 0 ),d_out => d192_out,en_out =>open  ,sof_out=>open   );


CL193: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d193_in(9*N-1 downto 8*N),data2conv2 =>d193_in(8*N-1 downto 7*N),data2conv3 =>d193_in(7*N-1 downto 6*N),data2conv4 =>d193_in(6*N-1 downto 5*N),data2conv5 =>d193_in(5*N-1 downto 4*N),data2conv6 =>d193_in(4*N-1 downto 3*N),data2conv7 =>d193_in(3*N-1 downto 2*N),data2conv8 =>d193_in(2*N-1 downto N),data2conv9 =>d193_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d193_in(9*N-1 downto 8*N),w2 => d193_in(8*N-1 downto 7*N),w3 => d193_in(7*N-1 downto 6*N),w4 => d193_in(6*N-1 downto 5*N),w5 => d193_in(5*N-1 downto 4*N),w6 => d193_in(4*N-1 downto 3*N),w7 => d193_in(3*N-1 downto 2*N),w8 => d193_in(2*N-1 downto N),w9 => d193_in(N-1 downto 0 ),d_out => d193_out,en_out =>open  ,sof_out=>open   );
CL194: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d194_in(9*N-1 downto 8*N),data2conv2 =>d194_in(8*N-1 downto 7*N),data2conv3 =>d194_in(7*N-1 downto 6*N),data2conv4 =>d194_in(6*N-1 downto 5*N),data2conv5 =>d194_in(5*N-1 downto 4*N),data2conv6 =>d194_in(4*N-1 downto 3*N),data2conv7 =>d194_in(3*N-1 downto 2*N),data2conv8 =>d194_in(2*N-1 downto N),data2conv9 =>d194_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d194_in(9*N-1 downto 8*N),w2 => d194_in(8*N-1 downto 7*N),w3 => d194_in(7*N-1 downto 6*N),w4 => d194_in(6*N-1 downto 5*N),w5 => d194_in(5*N-1 downto 4*N),w6 => d194_in(4*N-1 downto 3*N),w7 => d194_in(3*N-1 downto 2*N),w8 => d194_in(2*N-1 downto N),w9 => d194_in(N-1 downto 0 ),d_out => d194_out,en_out =>open  ,sof_out=>open   );
CL195: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d195_in(9*N-1 downto 8*N),data2conv2 =>d195_in(8*N-1 downto 7*N),data2conv3 =>d195_in(7*N-1 downto 6*N),data2conv4 =>d195_in(6*N-1 downto 5*N),data2conv5 =>d195_in(5*N-1 downto 4*N),data2conv6 =>d195_in(4*N-1 downto 3*N),data2conv7 =>d195_in(3*N-1 downto 2*N),data2conv8 =>d195_in(2*N-1 downto N),data2conv9 =>d195_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d195_in(9*N-1 downto 8*N),w2 => d195_in(8*N-1 downto 7*N),w3 => d195_in(7*N-1 downto 6*N),w4 => d195_in(6*N-1 downto 5*N),w5 => d195_in(5*N-1 downto 4*N),w6 => d195_in(4*N-1 downto 3*N),w7 => d195_in(3*N-1 downto 2*N),w8 => d195_in(2*N-1 downto N),w9 => d195_in(N-1 downto 0 ),d_out => d195_out,en_out =>open  ,sof_out=>open   );
CL196: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d196_in(9*N-1 downto 8*N),data2conv2 =>d196_in(8*N-1 downto 7*N),data2conv3 =>d196_in(7*N-1 downto 6*N),data2conv4 =>d196_in(6*N-1 downto 5*N),data2conv5 =>d196_in(5*N-1 downto 4*N),data2conv6 =>d196_in(4*N-1 downto 3*N),data2conv7 =>d196_in(3*N-1 downto 2*N),data2conv8 =>d196_in(2*N-1 downto N),data2conv9 =>d196_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d196_in(9*N-1 downto 8*N),w2 => d196_in(8*N-1 downto 7*N),w3 => d196_in(7*N-1 downto 6*N),w4 => d196_in(6*N-1 downto 5*N),w5 => d196_in(5*N-1 downto 4*N),w6 => d196_in(4*N-1 downto 3*N),w7 => d196_in(3*N-1 downto 2*N),w8 => d196_in(2*N-1 downto N),w9 => d196_in(N-1 downto 0 ),d_out => d196_out,en_out =>open  ,sof_out=>open   );
CL197: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d197_in(9*N-1 downto 8*N),data2conv2 =>d197_in(8*N-1 downto 7*N),data2conv3 =>d197_in(7*N-1 downto 6*N),data2conv4 =>d197_in(6*N-1 downto 5*N),data2conv5 =>d197_in(5*N-1 downto 4*N),data2conv6 =>d197_in(4*N-1 downto 3*N),data2conv7 =>d197_in(3*N-1 downto 2*N),data2conv8 =>d197_in(2*N-1 downto N),data2conv9 =>d197_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d197_in(9*N-1 downto 8*N),w2 => d197_in(8*N-1 downto 7*N),w3 => d197_in(7*N-1 downto 6*N),w4 => d197_in(6*N-1 downto 5*N),w5 => d197_in(5*N-1 downto 4*N),w6 => d197_in(4*N-1 downto 3*N),w7 => d197_in(3*N-1 downto 2*N),w8 => d197_in(2*N-1 downto N),w9 => d197_in(N-1 downto 0 ),d_out => d197_out,en_out =>open  ,sof_out=>open   );
CL198: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d198_in(9*N-1 downto 8*N),data2conv2 =>d198_in(8*N-1 downto 7*N),data2conv3 =>d198_in(7*N-1 downto 6*N),data2conv4 =>d198_in(6*N-1 downto 5*N),data2conv5 =>d198_in(5*N-1 downto 4*N),data2conv6 =>d198_in(4*N-1 downto 3*N),data2conv7 =>d198_in(3*N-1 downto 2*N),data2conv8 =>d198_in(2*N-1 downto N),data2conv9 =>d198_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d198_in(9*N-1 downto 8*N),w2 => d198_in(8*N-1 downto 7*N),w3 => d198_in(7*N-1 downto 6*N),w4 => d198_in(6*N-1 downto 5*N),w5 => d198_in(5*N-1 downto 4*N),w6 => d198_in(4*N-1 downto 3*N),w7 => d198_in(3*N-1 downto 2*N),w8 => d198_in(2*N-1 downto N),w9 => d198_in(N-1 downto 0 ),d_out => d198_out,en_out =>open  ,sof_out=>open   );
CL199: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d199_in(9*N-1 downto 8*N),data2conv2 =>d199_in(8*N-1 downto 7*N),data2conv3 =>d199_in(7*N-1 downto 6*N),data2conv4 =>d199_in(6*N-1 downto 5*N),data2conv5 =>d199_in(5*N-1 downto 4*N),data2conv6 =>d199_in(4*N-1 downto 3*N),data2conv7 =>d199_in(3*N-1 downto 2*N),data2conv8 =>d199_in(2*N-1 downto N),data2conv9 =>d199_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d199_in(9*N-1 downto 8*N),w2 => d199_in(8*N-1 downto 7*N),w3 => d199_in(7*N-1 downto 6*N),w4 => d199_in(6*N-1 downto 5*N),w5 => d199_in(5*N-1 downto 4*N),w6 => d199_in(4*N-1 downto 3*N),w7 => d199_in(3*N-1 downto 2*N),w8 => d199_in(2*N-1 downto N),w9 => d199_in(N-1 downto 0 ),d_out => d199_out,en_out =>open  ,sof_out=>open   );
CL200: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d200_in(9*N-1 downto 8*N),data2conv2 =>d200_in(8*N-1 downto 7*N),data2conv3 =>d200_in(7*N-1 downto 6*N),data2conv4 =>d200_in(6*N-1 downto 5*N),data2conv5 =>d200_in(5*N-1 downto 4*N),data2conv6 =>d200_in(4*N-1 downto 3*N),data2conv7 =>d200_in(3*N-1 downto 2*N),data2conv8 =>d200_in(2*N-1 downto N),data2conv9 =>d200_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d200_in(9*N-1 downto 8*N),w2 => d200_in(8*N-1 downto 7*N),w3 => d200_in(7*N-1 downto 6*N),w4 => d200_in(6*N-1 downto 5*N),w5 => d200_in(5*N-1 downto 4*N),w6 => d200_in(4*N-1 downto 3*N),w7 => d200_in(3*N-1 downto 2*N),w8 => d200_in(2*N-1 downto N),w9 => d200_in(N-1 downto 0 ),d_out => d200_out,en_out =>open  ,sof_out=>open   );
CL201: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d201_in(9*N-1 downto 8*N),data2conv2 =>d201_in(8*N-1 downto 7*N),data2conv3 =>d201_in(7*N-1 downto 6*N),data2conv4 =>d201_in(6*N-1 downto 5*N),data2conv5 =>d201_in(5*N-1 downto 4*N),data2conv6 =>d201_in(4*N-1 downto 3*N),data2conv7 =>d201_in(3*N-1 downto 2*N),data2conv8 =>d201_in(2*N-1 downto N),data2conv9 =>d201_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d201_in(9*N-1 downto 8*N),w2 => d201_in(8*N-1 downto 7*N),w3 => d201_in(7*N-1 downto 6*N),w4 => d201_in(6*N-1 downto 5*N),w5 => d201_in(5*N-1 downto 4*N),w6 => d201_in(4*N-1 downto 3*N),w7 => d201_in(3*N-1 downto 2*N),w8 => d201_in(2*N-1 downto N),w9 => d201_in(N-1 downto 0 ),d_out => d201_out,en_out =>open  ,sof_out=>open   );
CL202: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d202_in(9*N-1 downto 8*N),data2conv2 =>d202_in(8*N-1 downto 7*N),data2conv3 =>d202_in(7*N-1 downto 6*N),data2conv4 =>d202_in(6*N-1 downto 5*N),data2conv5 =>d202_in(5*N-1 downto 4*N),data2conv6 =>d202_in(4*N-1 downto 3*N),data2conv7 =>d202_in(3*N-1 downto 2*N),data2conv8 =>d202_in(2*N-1 downto N),data2conv9 =>d202_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d202_in(9*N-1 downto 8*N),w2 => d202_in(8*N-1 downto 7*N),w3 => d202_in(7*N-1 downto 6*N),w4 => d202_in(6*N-1 downto 5*N),w5 => d202_in(5*N-1 downto 4*N),w6 => d202_in(4*N-1 downto 3*N),w7 => d202_in(3*N-1 downto 2*N),w8 => d202_in(2*N-1 downto N),w9 => d202_in(N-1 downto 0 ),d_out => d202_out,en_out =>open  ,sof_out=>open   );
CL203: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d203_in(9*N-1 downto 8*N),data2conv2 =>d203_in(8*N-1 downto 7*N),data2conv3 =>d203_in(7*N-1 downto 6*N),data2conv4 =>d203_in(6*N-1 downto 5*N),data2conv5 =>d203_in(5*N-1 downto 4*N),data2conv6 =>d203_in(4*N-1 downto 3*N),data2conv7 =>d203_in(3*N-1 downto 2*N),data2conv8 =>d203_in(2*N-1 downto N),data2conv9 =>d203_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d203_in(9*N-1 downto 8*N),w2 => d203_in(8*N-1 downto 7*N),w3 => d203_in(7*N-1 downto 6*N),w4 => d203_in(6*N-1 downto 5*N),w5 => d203_in(5*N-1 downto 4*N),w6 => d203_in(4*N-1 downto 3*N),w7 => d203_in(3*N-1 downto 2*N),w8 => d203_in(2*N-1 downto N),w9 => d203_in(N-1 downto 0 ),d_out => d203_out,en_out =>open  ,sof_out=>open   );
CL204: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d204_in(9*N-1 downto 8*N),data2conv2 =>d204_in(8*N-1 downto 7*N),data2conv3 =>d204_in(7*N-1 downto 6*N),data2conv4 =>d204_in(6*N-1 downto 5*N),data2conv5 =>d204_in(5*N-1 downto 4*N),data2conv6 =>d204_in(4*N-1 downto 3*N),data2conv7 =>d204_in(3*N-1 downto 2*N),data2conv8 =>d204_in(2*N-1 downto N),data2conv9 =>d204_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d204_in(9*N-1 downto 8*N),w2 => d204_in(8*N-1 downto 7*N),w3 => d204_in(7*N-1 downto 6*N),w4 => d204_in(6*N-1 downto 5*N),w5 => d204_in(5*N-1 downto 4*N),w6 => d204_in(4*N-1 downto 3*N),w7 => d204_in(3*N-1 downto 2*N),w8 => d204_in(2*N-1 downto N),w9 => d204_in(N-1 downto 0 ),d_out => d204_out,en_out =>open  ,sof_out=>open   );
CL205: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d205_in(9*N-1 downto 8*N),data2conv2 =>d205_in(8*N-1 downto 7*N),data2conv3 =>d205_in(7*N-1 downto 6*N),data2conv4 =>d205_in(6*N-1 downto 5*N),data2conv5 =>d205_in(5*N-1 downto 4*N),data2conv6 =>d205_in(4*N-1 downto 3*N),data2conv7 =>d205_in(3*N-1 downto 2*N),data2conv8 =>d205_in(2*N-1 downto N),data2conv9 =>d205_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d205_in(9*N-1 downto 8*N),w2 => d205_in(8*N-1 downto 7*N),w3 => d205_in(7*N-1 downto 6*N),w4 => d205_in(6*N-1 downto 5*N),w5 => d205_in(5*N-1 downto 4*N),w6 => d205_in(4*N-1 downto 3*N),w7 => d205_in(3*N-1 downto 2*N),w8 => d205_in(2*N-1 downto N),w9 => d205_in(N-1 downto 0 ),d_out => d205_out,en_out =>open  ,sof_out=>open   );
CL206: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d206_in(9*N-1 downto 8*N),data2conv2 =>d206_in(8*N-1 downto 7*N),data2conv3 =>d206_in(7*N-1 downto 6*N),data2conv4 =>d206_in(6*N-1 downto 5*N),data2conv5 =>d206_in(5*N-1 downto 4*N),data2conv6 =>d206_in(4*N-1 downto 3*N),data2conv7 =>d206_in(3*N-1 downto 2*N),data2conv8 =>d206_in(2*N-1 downto N),data2conv9 =>d206_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d206_in(9*N-1 downto 8*N),w2 => d206_in(8*N-1 downto 7*N),w3 => d206_in(7*N-1 downto 6*N),w4 => d206_in(6*N-1 downto 5*N),w5 => d206_in(5*N-1 downto 4*N),w6 => d206_in(4*N-1 downto 3*N),w7 => d206_in(3*N-1 downto 2*N),w8 => d206_in(2*N-1 downto N),w9 => d206_in(N-1 downto 0 ),d_out => d206_out,en_out =>open  ,sof_out=>open   );
CL207: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d207_in(9*N-1 downto 8*N),data2conv2 =>d207_in(8*N-1 downto 7*N),data2conv3 =>d207_in(7*N-1 downto 6*N),data2conv4 =>d207_in(6*N-1 downto 5*N),data2conv5 =>d207_in(5*N-1 downto 4*N),data2conv6 =>d207_in(4*N-1 downto 3*N),data2conv7 =>d207_in(3*N-1 downto 2*N),data2conv8 =>d207_in(2*N-1 downto N),data2conv9 =>d207_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d207_in(9*N-1 downto 8*N),w2 => d207_in(8*N-1 downto 7*N),w3 => d207_in(7*N-1 downto 6*N),w4 => d207_in(6*N-1 downto 5*N),w5 => d207_in(5*N-1 downto 4*N),w6 => d207_in(4*N-1 downto 3*N),w7 => d207_in(3*N-1 downto 2*N),w8 => d207_in(2*N-1 downto N),w9 => d207_in(N-1 downto 0 ),d_out => d207_out,en_out =>open  ,sof_out=>open   );
CL208: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d208_in(9*N-1 downto 8*N),data2conv2 =>d208_in(8*N-1 downto 7*N),data2conv3 =>d208_in(7*N-1 downto 6*N),data2conv4 =>d208_in(6*N-1 downto 5*N),data2conv5 =>d208_in(5*N-1 downto 4*N),data2conv6 =>d208_in(4*N-1 downto 3*N),data2conv7 =>d208_in(3*N-1 downto 2*N),data2conv8 =>d208_in(2*N-1 downto N),data2conv9 =>d208_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d208_in(9*N-1 downto 8*N),w2 => d208_in(8*N-1 downto 7*N),w3 => d208_in(7*N-1 downto 6*N),w4 => d208_in(6*N-1 downto 5*N),w5 => d208_in(5*N-1 downto 4*N),w6 => d208_in(4*N-1 downto 3*N),w7 => d208_in(3*N-1 downto 2*N),w8 => d208_in(2*N-1 downto N),w9 => d208_in(N-1 downto 0 ),d_out => d208_out,en_out =>open  ,sof_out=>open   );
CL209: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d209_in(9*N-1 downto 8*N),data2conv2 =>d209_in(8*N-1 downto 7*N),data2conv3 =>d209_in(7*N-1 downto 6*N),data2conv4 =>d209_in(6*N-1 downto 5*N),data2conv5 =>d209_in(5*N-1 downto 4*N),data2conv6 =>d209_in(4*N-1 downto 3*N),data2conv7 =>d209_in(3*N-1 downto 2*N),data2conv8 =>d209_in(2*N-1 downto N),data2conv9 =>d209_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d209_in(9*N-1 downto 8*N),w2 => d209_in(8*N-1 downto 7*N),w3 => d209_in(7*N-1 downto 6*N),w4 => d209_in(6*N-1 downto 5*N),w5 => d209_in(5*N-1 downto 4*N),w6 => d209_in(4*N-1 downto 3*N),w7 => d209_in(3*N-1 downto 2*N),w8 => d209_in(2*N-1 downto N),w9 => d209_in(N-1 downto 0 ),d_out => d209_out,en_out =>open  ,sof_out=>open   );
CL210: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d210_in(9*N-1 downto 8*N),data2conv2 =>d210_in(8*N-1 downto 7*N),data2conv3 =>d210_in(7*N-1 downto 6*N),data2conv4 =>d210_in(6*N-1 downto 5*N),data2conv5 =>d210_in(5*N-1 downto 4*N),data2conv6 =>d210_in(4*N-1 downto 3*N),data2conv7 =>d210_in(3*N-1 downto 2*N),data2conv8 =>d210_in(2*N-1 downto N),data2conv9 =>d210_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d210_in(9*N-1 downto 8*N),w2 => d210_in(8*N-1 downto 7*N),w3 => d210_in(7*N-1 downto 6*N),w4 => d210_in(6*N-1 downto 5*N),w5 => d210_in(5*N-1 downto 4*N),w6 => d210_in(4*N-1 downto 3*N),w7 => d210_in(3*N-1 downto 2*N),w8 => d210_in(2*N-1 downto N),w9 => d210_in(N-1 downto 0 ),d_out => d210_out,en_out =>open  ,sof_out=>open   );
CL211: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d211_in(9*N-1 downto 8*N),data2conv2 =>d211_in(8*N-1 downto 7*N),data2conv3 =>d211_in(7*N-1 downto 6*N),data2conv4 =>d211_in(6*N-1 downto 5*N),data2conv5 =>d211_in(5*N-1 downto 4*N),data2conv6 =>d211_in(4*N-1 downto 3*N),data2conv7 =>d211_in(3*N-1 downto 2*N),data2conv8 =>d211_in(2*N-1 downto N),data2conv9 =>d211_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d211_in(9*N-1 downto 8*N),w2 => d211_in(8*N-1 downto 7*N),w3 => d211_in(7*N-1 downto 6*N),w4 => d211_in(6*N-1 downto 5*N),w5 => d211_in(5*N-1 downto 4*N),w6 => d211_in(4*N-1 downto 3*N),w7 => d211_in(3*N-1 downto 2*N),w8 => d211_in(2*N-1 downto N),w9 => d211_in(N-1 downto 0 ),d_out => d211_out,en_out =>open  ,sof_out=>open   );
CL212: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d212_in(9*N-1 downto 8*N),data2conv2 =>d212_in(8*N-1 downto 7*N),data2conv3 =>d212_in(7*N-1 downto 6*N),data2conv4 =>d212_in(6*N-1 downto 5*N),data2conv5 =>d212_in(5*N-1 downto 4*N),data2conv6 =>d212_in(4*N-1 downto 3*N),data2conv7 =>d212_in(3*N-1 downto 2*N),data2conv8 =>d212_in(2*N-1 downto N),data2conv9 =>d212_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d212_in(9*N-1 downto 8*N),w2 => d212_in(8*N-1 downto 7*N),w3 => d212_in(7*N-1 downto 6*N),w4 => d212_in(6*N-1 downto 5*N),w5 => d212_in(5*N-1 downto 4*N),w6 => d212_in(4*N-1 downto 3*N),w7 => d212_in(3*N-1 downto 2*N),w8 => d212_in(2*N-1 downto N),w9 => d212_in(N-1 downto 0 ),d_out => d212_out,en_out =>open  ,sof_out=>open   );
CL213: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d213_in(9*N-1 downto 8*N),data2conv2 =>d213_in(8*N-1 downto 7*N),data2conv3 =>d213_in(7*N-1 downto 6*N),data2conv4 =>d213_in(6*N-1 downto 5*N),data2conv5 =>d213_in(5*N-1 downto 4*N),data2conv6 =>d213_in(4*N-1 downto 3*N),data2conv7 =>d213_in(3*N-1 downto 2*N),data2conv8 =>d213_in(2*N-1 downto N),data2conv9 =>d213_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d213_in(9*N-1 downto 8*N),w2 => d213_in(8*N-1 downto 7*N),w3 => d213_in(7*N-1 downto 6*N),w4 => d213_in(6*N-1 downto 5*N),w5 => d213_in(5*N-1 downto 4*N),w6 => d213_in(4*N-1 downto 3*N),w7 => d213_in(3*N-1 downto 2*N),w8 => d213_in(2*N-1 downto N),w9 => d213_in(N-1 downto 0 ),d_out => d213_out,en_out =>open  ,sof_out=>open   );
CL214: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d214_in(9*N-1 downto 8*N),data2conv2 =>d214_in(8*N-1 downto 7*N),data2conv3 =>d214_in(7*N-1 downto 6*N),data2conv4 =>d214_in(6*N-1 downto 5*N),data2conv5 =>d214_in(5*N-1 downto 4*N),data2conv6 =>d214_in(4*N-1 downto 3*N),data2conv7 =>d214_in(3*N-1 downto 2*N),data2conv8 =>d214_in(2*N-1 downto N),data2conv9 =>d214_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d214_in(9*N-1 downto 8*N),w2 => d214_in(8*N-1 downto 7*N),w3 => d214_in(7*N-1 downto 6*N),w4 => d214_in(6*N-1 downto 5*N),w5 => d214_in(5*N-1 downto 4*N),w6 => d214_in(4*N-1 downto 3*N),w7 => d214_in(3*N-1 downto 2*N),w8 => d214_in(2*N-1 downto N),w9 => d214_in(N-1 downto 0 ),d_out => d214_out,en_out =>open  ,sof_out=>open   );
CL215: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d215_in(9*N-1 downto 8*N),data2conv2 =>d215_in(8*N-1 downto 7*N),data2conv3 =>d215_in(7*N-1 downto 6*N),data2conv4 =>d215_in(6*N-1 downto 5*N),data2conv5 =>d215_in(5*N-1 downto 4*N),data2conv6 =>d215_in(4*N-1 downto 3*N),data2conv7 =>d215_in(3*N-1 downto 2*N),data2conv8 =>d215_in(2*N-1 downto N),data2conv9 =>d215_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d215_in(9*N-1 downto 8*N),w2 => d215_in(8*N-1 downto 7*N),w3 => d215_in(7*N-1 downto 6*N),w4 => d215_in(6*N-1 downto 5*N),w5 => d215_in(5*N-1 downto 4*N),w6 => d215_in(4*N-1 downto 3*N),w7 => d215_in(3*N-1 downto 2*N),w8 => d215_in(2*N-1 downto N),w9 => d215_in(N-1 downto 0 ),d_out => d215_out,en_out =>open  ,sof_out=>open   );
CL216: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d216_in(9*N-1 downto 8*N),data2conv2 =>d216_in(8*N-1 downto 7*N),data2conv3 =>d216_in(7*N-1 downto 6*N),data2conv4 =>d216_in(6*N-1 downto 5*N),data2conv5 =>d216_in(5*N-1 downto 4*N),data2conv6 =>d216_in(4*N-1 downto 3*N),data2conv7 =>d216_in(3*N-1 downto 2*N),data2conv8 =>d216_in(2*N-1 downto N),data2conv9 =>d216_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d216_in(9*N-1 downto 8*N),w2 => d216_in(8*N-1 downto 7*N),w3 => d216_in(7*N-1 downto 6*N),w4 => d216_in(6*N-1 downto 5*N),w5 => d216_in(5*N-1 downto 4*N),w6 => d216_in(4*N-1 downto 3*N),w7 => d216_in(3*N-1 downto 2*N),w8 => d216_in(2*N-1 downto N),w9 => d216_in(N-1 downto 0 ),d_out => d216_out,en_out =>open  ,sof_out=>open   );
CL217: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d217_in(9*N-1 downto 8*N),data2conv2 =>d217_in(8*N-1 downto 7*N),data2conv3 =>d217_in(7*N-1 downto 6*N),data2conv4 =>d217_in(6*N-1 downto 5*N),data2conv5 =>d217_in(5*N-1 downto 4*N),data2conv6 =>d217_in(4*N-1 downto 3*N),data2conv7 =>d217_in(3*N-1 downto 2*N),data2conv8 =>d217_in(2*N-1 downto N),data2conv9 =>d217_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d217_in(9*N-1 downto 8*N),w2 => d217_in(8*N-1 downto 7*N),w3 => d217_in(7*N-1 downto 6*N),w4 => d217_in(6*N-1 downto 5*N),w5 => d217_in(5*N-1 downto 4*N),w6 => d217_in(4*N-1 downto 3*N),w7 => d217_in(3*N-1 downto 2*N),w8 => d217_in(2*N-1 downto N),w9 => d217_in(N-1 downto 0 ),d_out => d217_out,en_out =>open  ,sof_out=>open   );
CL218: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d218_in(9*N-1 downto 8*N),data2conv2 =>d218_in(8*N-1 downto 7*N),data2conv3 =>d218_in(7*N-1 downto 6*N),data2conv4 =>d218_in(6*N-1 downto 5*N),data2conv5 =>d218_in(5*N-1 downto 4*N),data2conv6 =>d218_in(4*N-1 downto 3*N),data2conv7 =>d218_in(3*N-1 downto 2*N),data2conv8 =>d218_in(2*N-1 downto N),data2conv9 =>d218_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d218_in(9*N-1 downto 8*N),w2 => d218_in(8*N-1 downto 7*N),w3 => d218_in(7*N-1 downto 6*N),w4 => d218_in(6*N-1 downto 5*N),w5 => d218_in(5*N-1 downto 4*N),w6 => d218_in(4*N-1 downto 3*N),w7 => d218_in(3*N-1 downto 2*N),w8 => d218_in(2*N-1 downto N),w9 => d218_in(N-1 downto 0 ),d_out => d218_out,en_out =>open  ,sof_out=>open   );
CL219: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d219_in(9*N-1 downto 8*N),data2conv2 =>d219_in(8*N-1 downto 7*N),data2conv3 =>d219_in(7*N-1 downto 6*N),data2conv4 =>d219_in(6*N-1 downto 5*N),data2conv5 =>d219_in(5*N-1 downto 4*N),data2conv6 =>d219_in(4*N-1 downto 3*N),data2conv7 =>d219_in(3*N-1 downto 2*N),data2conv8 =>d219_in(2*N-1 downto N),data2conv9 =>d219_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d219_in(9*N-1 downto 8*N),w2 => d219_in(8*N-1 downto 7*N),w3 => d219_in(7*N-1 downto 6*N),w4 => d219_in(6*N-1 downto 5*N),w5 => d219_in(5*N-1 downto 4*N),w6 => d219_in(4*N-1 downto 3*N),w7 => d219_in(3*N-1 downto 2*N),w8 => d219_in(2*N-1 downto N),w9 => d219_in(N-1 downto 0 ),d_out => d219_out,en_out =>open  ,sof_out=>open   );
CL220: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d220_in(9*N-1 downto 8*N),data2conv2 =>d220_in(8*N-1 downto 7*N),data2conv3 =>d220_in(7*N-1 downto 6*N),data2conv4 =>d220_in(6*N-1 downto 5*N),data2conv5 =>d220_in(5*N-1 downto 4*N),data2conv6 =>d220_in(4*N-1 downto 3*N),data2conv7 =>d220_in(3*N-1 downto 2*N),data2conv8 =>d220_in(2*N-1 downto N),data2conv9 =>d220_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d220_in(9*N-1 downto 8*N),w2 => d220_in(8*N-1 downto 7*N),w3 => d220_in(7*N-1 downto 6*N),w4 => d220_in(6*N-1 downto 5*N),w5 => d220_in(5*N-1 downto 4*N),w6 => d220_in(4*N-1 downto 3*N),w7 => d220_in(3*N-1 downto 2*N),w8 => d220_in(2*N-1 downto N),w9 => d220_in(N-1 downto 0 ),d_out => d220_out,en_out =>open  ,sof_out=>open   );
CL221: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d221_in(9*N-1 downto 8*N),data2conv2 =>d221_in(8*N-1 downto 7*N),data2conv3 =>d221_in(7*N-1 downto 6*N),data2conv4 =>d221_in(6*N-1 downto 5*N),data2conv5 =>d221_in(5*N-1 downto 4*N),data2conv6 =>d221_in(4*N-1 downto 3*N),data2conv7 =>d221_in(3*N-1 downto 2*N),data2conv8 =>d221_in(2*N-1 downto N),data2conv9 =>d221_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d221_in(9*N-1 downto 8*N),w2 => d221_in(8*N-1 downto 7*N),w3 => d221_in(7*N-1 downto 6*N),w4 => d221_in(6*N-1 downto 5*N),w5 => d221_in(5*N-1 downto 4*N),w6 => d221_in(4*N-1 downto 3*N),w7 => d221_in(3*N-1 downto 2*N),w8 => d221_in(2*N-1 downto N),w9 => d221_in(N-1 downto 0 ),d_out => d221_out,en_out =>open  ,sof_out=>open   );
CL222: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d222_in(9*N-1 downto 8*N),data2conv2 =>d222_in(8*N-1 downto 7*N),data2conv3 =>d222_in(7*N-1 downto 6*N),data2conv4 =>d222_in(6*N-1 downto 5*N),data2conv5 =>d222_in(5*N-1 downto 4*N),data2conv6 =>d222_in(4*N-1 downto 3*N),data2conv7 =>d222_in(3*N-1 downto 2*N),data2conv8 =>d222_in(2*N-1 downto N),data2conv9 =>d222_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d222_in(9*N-1 downto 8*N),w2 => d222_in(8*N-1 downto 7*N),w3 => d222_in(7*N-1 downto 6*N),w4 => d222_in(6*N-1 downto 5*N),w5 => d222_in(5*N-1 downto 4*N),w6 => d222_in(4*N-1 downto 3*N),w7 => d222_in(3*N-1 downto 2*N),w8 => d222_in(2*N-1 downto N),w9 => d222_in(N-1 downto 0 ),d_out => d222_out,en_out =>open  ,sof_out=>open   );
CL223: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d223_in(9*N-1 downto 8*N),data2conv2 =>d223_in(8*N-1 downto 7*N),data2conv3 =>d223_in(7*N-1 downto 6*N),data2conv4 =>d223_in(6*N-1 downto 5*N),data2conv5 =>d223_in(5*N-1 downto 4*N),data2conv6 =>d223_in(4*N-1 downto 3*N),data2conv7 =>d223_in(3*N-1 downto 2*N),data2conv8 =>d223_in(2*N-1 downto N),data2conv9 =>d223_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d223_in(9*N-1 downto 8*N),w2 => d223_in(8*N-1 downto 7*N),w3 => d223_in(7*N-1 downto 6*N),w4 => d223_in(6*N-1 downto 5*N),w5 => d223_in(5*N-1 downto 4*N),w6 => d223_in(4*N-1 downto 3*N),w7 => d223_in(3*N-1 downto 2*N),w8 => d223_in(2*N-1 downto N),w9 => d223_in(N-1 downto 0 ),d_out => d223_out,en_out =>open  ,sof_out=>open   );
CL224: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d224_in(9*N-1 downto 8*N),data2conv2 =>d224_in(8*N-1 downto 7*N),data2conv3 =>d224_in(7*N-1 downto 6*N),data2conv4 =>d224_in(6*N-1 downto 5*N),data2conv5 =>d224_in(5*N-1 downto 4*N),data2conv6 =>d224_in(4*N-1 downto 3*N),data2conv7 =>d224_in(3*N-1 downto 2*N),data2conv8 =>d224_in(2*N-1 downto N),data2conv9 =>d224_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d224_in(9*N-1 downto 8*N),w2 => d224_in(8*N-1 downto 7*N),w3 => d224_in(7*N-1 downto 6*N),w4 => d224_in(6*N-1 downto 5*N),w5 => d224_in(5*N-1 downto 4*N),w6 => d224_in(4*N-1 downto 3*N),w7 => d224_in(3*N-1 downto 2*N),w8 => d224_in(2*N-1 downto N),w9 => d224_in(N-1 downto 0 ),d_out => d224_out,en_out =>open  ,sof_out=>open   );
CL225: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d225_in(9*N-1 downto 8*N),data2conv2 =>d225_in(8*N-1 downto 7*N),data2conv3 =>d225_in(7*N-1 downto 6*N),data2conv4 =>d225_in(6*N-1 downto 5*N),data2conv5 =>d225_in(5*N-1 downto 4*N),data2conv6 =>d225_in(4*N-1 downto 3*N),data2conv7 =>d225_in(3*N-1 downto 2*N),data2conv8 =>d225_in(2*N-1 downto N),data2conv9 =>d225_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d225_in(9*N-1 downto 8*N),w2 => d225_in(8*N-1 downto 7*N),w3 => d225_in(7*N-1 downto 6*N),w4 => d225_in(6*N-1 downto 5*N),w5 => d225_in(5*N-1 downto 4*N),w6 => d225_in(4*N-1 downto 3*N),w7 => d225_in(3*N-1 downto 2*N),w8 => d225_in(2*N-1 downto N),w9 => d225_in(N-1 downto 0 ),d_out => d225_out,en_out =>open  ,sof_out=>open   );
CL226: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d226_in(9*N-1 downto 8*N),data2conv2 =>d226_in(8*N-1 downto 7*N),data2conv3 =>d226_in(7*N-1 downto 6*N),data2conv4 =>d226_in(6*N-1 downto 5*N),data2conv5 =>d226_in(5*N-1 downto 4*N),data2conv6 =>d226_in(4*N-1 downto 3*N),data2conv7 =>d226_in(3*N-1 downto 2*N),data2conv8 =>d226_in(2*N-1 downto N),data2conv9 =>d226_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d226_in(9*N-1 downto 8*N),w2 => d226_in(8*N-1 downto 7*N),w3 => d226_in(7*N-1 downto 6*N),w4 => d226_in(6*N-1 downto 5*N),w5 => d226_in(5*N-1 downto 4*N),w6 => d226_in(4*N-1 downto 3*N),w7 => d226_in(3*N-1 downto 2*N),w8 => d226_in(2*N-1 downto N),w9 => d226_in(N-1 downto 0 ),d_out => d226_out,en_out =>open  ,sof_out=>open   );
CL227: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d227_in(9*N-1 downto 8*N),data2conv2 =>d227_in(8*N-1 downto 7*N),data2conv3 =>d227_in(7*N-1 downto 6*N),data2conv4 =>d227_in(6*N-1 downto 5*N),data2conv5 =>d227_in(5*N-1 downto 4*N),data2conv6 =>d227_in(4*N-1 downto 3*N),data2conv7 =>d227_in(3*N-1 downto 2*N),data2conv8 =>d227_in(2*N-1 downto N),data2conv9 =>d227_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d227_in(9*N-1 downto 8*N),w2 => d227_in(8*N-1 downto 7*N),w3 => d227_in(7*N-1 downto 6*N),w4 => d227_in(6*N-1 downto 5*N),w5 => d227_in(5*N-1 downto 4*N),w6 => d227_in(4*N-1 downto 3*N),w7 => d227_in(3*N-1 downto 2*N),w8 => d227_in(2*N-1 downto N),w9 => d227_in(N-1 downto 0 ),d_out => d227_out,en_out =>open  ,sof_out=>open   );
CL228: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d228_in(9*N-1 downto 8*N),data2conv2 =>d228_in(8*N-1 downto 7*N),data2conv3 =>d228_in(7*N-1 downto 6*N),data2conv4 =>d228_in(6*N-1 downto 5*N),data2conv5 =>d228_in(5*N-1 downto 4*N),data2conv6 =>d228_in(4*N-1 downto 3*N),data2conv7 =>d228_in(3*N-1 downto 2*N),data2conv8 =>d228_in(2*N-1 downto N),data2conv9 =>d228_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d228_in(9*N-1 downto 8*N),w2 => d228_in(8*N-1 downto 7*N),w3 => d228_in(7*N-1 downto 6*N),w4 => d228_in(6*N-1 downto 5*N),w5 => d228_in(5*N-1 downto 4*N),w6 => d228_in(4*N-1 downto 3*N),w7 => d228_in(3*N-1 downto 2*N),w8 => d228_in(2*N-1 downto N),w9 => d228_in(N-1 downto 0 ),d_out => d228_out,en_out =>open  ,sof_out=>open   );
CL229: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d229_in(9*N-1 downto 8*N),data2conv2 =>d229_in(8*N-1 downto 7*N),data2conv3 =>d229_in(7*N-1 downto 6*N),data2conv4 =>d229_in(6*N-1 downto 5*N),data2conv5 =>d229_in(5*N-1 downto 4*N),data2conv6 =>d229_in(4*N-1 downto 3*N),data2conv7 =>d229_in(3*N-1 downto 2*N),data2conv8 =>d229_in(2*N-1 downto N),data2conv9 =>d229_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d229_in(9*N-1 downto 8*N),w2 => d229_in(8*N-1 downto 7*N),w3 => d229_in(7*N-1 downto 6*N),w4 => d229_in(6*N-1 downto 5*N),w5 => d229_in(5*N-1 downto 4*N),w6 => d229_in(4*N-1 downto 3*N),w7 => d229_in(3*N-1 downto 2*N),w8 => d229_in(2*N-1 downto N),w9 => d229_in(N-1 downto 0 ),d_out => d229_out,en_out =>open  ,sof_out=>open   );
CL230: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d230_in(9*N-1 downto 8*N),data2conv2 =>d230_in(8*N-1 downto 7*N),data2conv3 =>d230_in(7*N-1 downto 6*N),data2conv4 =>d230_in(6*N-1 downto 5*N),data2conv5 =>d230_in(5*N-1 downto 4*N),data2conv6 =>d230_in(4*N-1 downto 3*N),data2conv7 =>d230_in(3*N-1 downto 2*N),data2conv8 =>d230_in(2*N-1 downto N),data2conv9 =>d230_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d230_in(9*N-1 downto 8*N),w2 => d230_in(8*N-1 downto 7*N),w3 => d230_in(7*N-1 downto 6*N),w4 => d230_in(6*N-1 downto 5*N),w5 => d230_in(5*N-1 downto 4*N),w6 => d230_in(4*N-1 downto 3*N),w7 => d230_in(3*N-1 downto 2*N),w8 => d230_in(2*N-1 downto N),w9 => d230_in(N-1 downto 0 ),d_out => d230_out,en_out =>open  ,sof_out=>open   );
CL231: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d231_in(9*N-1 downto 8*N),data2conv2 =>d231_in(8*N-1 downto 7*N),data2conv3 =>d231_in(7*N-1 downto 6*N),data2conv4 =>d231_in(6*N-1 downto 5*N),data2conv5 =>d231_in(5*N-1 downto 4*N),data2conv6 =>d231_in(4*N-1 downto 3*N),data2conv7 =>d231_in(3*N-1 downto 2*N),data2conv8 =>d231_in(2*N-1 downto N),data2conv9 =>d231_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d231_in(9*N-1 downto 8*N),w2 => d231_in(8*N-1 downto 7*N),w3 => d231_in(7*N-1 downto 6*N),w4 => d231_in(6*N-1 downto 5*N),w5 => d231_in(5*N-1 downto 4*N),w6 => d231_in(4*N-1 downto 3*N),w7 => d231_in(3*N-1 downto 2*N),w8 => d231_in(2*N-1 downto N),w9 => d231_in(N-1 downto 0 ),d_out => d231_out,en_out =>open  ,sof_out=>open   );
CL232: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d232_in(9*N-1 downto 8*N),data2conv2 =>d232_in(8*N-1 downto 7*N),data2conv3 =>d232_in(7*N-1 downto 6*N),data2conv4 =>d232_in(6*N-1 downto 5*N),data2conv5 =>d232_in(5*N-1 downto 4*N),data2conv6 =>d232_in(4*N-1 downto 3*N),data2conv7 =>d232_in(3*N-1 downto 2*N),data2conv8 =>d232_in(2*N-1 downto N),data2conv9 =>d232_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d232_in(9*N-1 downto 8*N),w2 => d232_in(8*N-1 downto 7*N),w3 => d232_in(7*N-1 downto 6*N),w4 => d232_in(6*N-1 downto 5*N),w5 => d232_in(5*N-1 downto 4*N),w6 => d232_in(4*N-1 downto 3*N),w7 => d232_in(3*N-1 downto 2*N),w8 => d232_in(2*N-1 downto N),w9 => d232_in(N-1 downto 0 ),d_out => d232_out,en_out =>open  ,sof_out=>open   );
CL233: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d233_in(9*N-1 downto 8*N),data2conv2 =>d233_in(8*N-1 downto 7*N),data2conv3 =>d233_in(7*N-1 downto 6*N),data2conv4 =>d233_in(6*N-1 downto 5*N),data2conv5 =>d233_in(5*N-1 downto 4*N),data2conv6 =>d233_in(4*N-1 downto 3*N),data2conv7 =>d233_in(3*N-1 downto 2*N),data2conv8 =>d233_in(2*N-1 downto N),data2conv9 =>d233_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d233_in(9*N-1 downto 8*N),w2 => d233_in(8*N-1 downto 7*N),w3 => d233_in(7*N-1 downto 6*N),w4 => d233_in(6*N-1 downto 5*N),w5 => d233_in(5*N-1 downto 4*N),w6 => d233_in(4*N-1 downto 3*N),w7 => d233_in(3*N-1 downto 2*N),w8 => d233_in(2*N-1 downto N),w9 => d233_in(N-1 downto 0 ),d_out => d233_out,en_out =>open  ,sof_out=>open   );
CL234: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d234_in(9*N-1 downto 8*N),data2conv2 =>d234_in(8*N-1 downto 7*N),data2conv3 =>d234_in(7*N-1 downto 6*N),data2conv4 =>d234_in(6*N-1 downto 5*N),data2conv5 =>d234_in(5*N-1 downto 4*N),data2conv6 =>d234_in(4*N-1 downto 3*N),data2conv7 =>d234_in(3*N-1 downto 2*N),data2conv8 =>d234_in(2*N-1 downto N),data2conv9 =>d234_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d234_in(9*N-1 downto 8*N),w2 => d234_in(8*N-1 downto 7*N),w3 => d234_in(7*N-1 downto 6*N),w4 => d234_in(6*N-1 downto 5*N),w5 => d234_in(5*N-1 downto 4*N),w6 => d234_in(4*N-1 downto 3*N),w7 => d234_in(3*N-1 downto 2*N),w8 => d234_in(2*N-1 downto N),w9 => d234_in(N-1 downto 0 ),d_out => d234_out,en_out =>open  ,sof_out=>open   );
CL235: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d235_in(9*N-1 downto 8*N),data2conv2 =>d235_in(8*N-1 downto 7*N),data2conv3 =>d235_in(7*N-1 downto 6*N),data2conv4 =>d235_in(6*N-1 downto 5*N),data2conv5 =>d235_in(5*N-1 downto 4*N),data2conv6 =>d235_in(4*N-1 downto 3*N),data2conv7 =>d235_in(3*N-1 downto 2*N),data2conv8 =>d235_in(2*N-1 downto N),data2conv9 =>d235_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d235_in(9*N-1 downto 8*N),w2 => d235_in(8*N-1 downto 7*N),w3 => d235_in(7*N-1 downto 6*N),w4 => d235_in(6*N-1 downto 5*N),w5 => d235_in(5*N-1 downto 4*N),w6 => d235_in(4*N-1 downto 3*N),w7 => d235_in(3*N-1 downto 2*N),w8 => d235_in(2*N-1 downto N),w9 => d235_in(N-1 downto 0 ),d_out => d235_out,en_out =>open  ,sof_out=>open   );
CL236: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d236_in(9*N-1 downto 8*N),data2conv2 =>d236_in(8*N-1 downto 7*N),data2conv3 =>d236_in(7*N-1 downto 6*N),data2conv4 =>d236_in(6*N-1 downto 5*N),data2conv5 =>d236_in(5*N-1 downto 4*N),data2conv6 =>d236_in(4*N-1 downto 3*N),data2conv7 =>d236_in(3*N-1 downto 2*N),data2conv8 =>d236_in(2*N-1 downto N),data2conv9 =>d236_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d236_in(9*N-1 downto 8*N),w2 => d236_in(8*N-1 downto 7*N),w3 => d236_in(7*N-1 downto 6*N),w4 => d236_in(6*N-1 downto 5*N),w5 => d236_in(5*N-1 downto 4*N),w6 => d236_in(4*N-1 downto 3*N),w7 => d236_in(3*N-1 downto 2*N),w8 => d236_in(2*N-1 downto N),w9 => d236_in(N-1 downto 0 ),d_out => d236_out,en_out =>open  ,sof_out=>open   );
CL237: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d237_in(9*N-1 downto 8*N),data2conv2 =>d237_in(8*N-1 downto 7*N),data2conv3 =>d237_in(7*N-1 downto 6*N),data2conv4 =>d237_in(6*N-1 downto 5*N),data2conv5 =>d237_in(5*N-1 downto 4*N),data2conv6 =>d237_in(4*N-1 downto 3*N),data2conv7 =>d237_in(3*N-1 downto 2*N),data2conv8 =>d237_in(2*N-1 downto N),data2conv9 =>d237_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d237_in(9*N-1 downto 8*N),w2 => d237_in(8*N-1 downto 7*N),w3 => d237_in(7*N-1 downto 6*N),w4 => d237_in(6*N-1 downto 5*N),w5 => d237_in(5*N-1 downto 4*N),w6 => d237_in(4*N-1 downto 3*N),w7 => d237_in(3*N-1 downto 2*N),w8 => d237_in(2*N-1 downto N),w9 => d237_in(N-1 downto 0 ),d_out => d237_out,en_out =>open  ,sof_out=>open   );
CL238: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d238_in(9*N-1 downto 8*N),data2conv2 =>d238_in(8*N-1 downto 7*N),data2conv3 =>d238_in(7*N-1 downto 6*N),data2conv4 =>d238_in(6*N-1 downto 5*N),data2conv5 =>d238_in(5*N-1 downto 4*N),data2conv6 =>d238_in(4*N-1 downto 3*N),data2conv7 =>d238_in(3*N-1 downto 2*N),data2conv8 =>d238_in(2*N-1 downto N),data2conv9 =>d238_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d238_in(9*N-1 downto 8*N),w2 => d238_in(8*N-1 downto 7*N),w3 => d238_in(7*N-1 downto 6*N),w4 => d238_in(6*N-1 downto 5*N),w5 => d238_in(5*N-1 downto 4*N),w6 => d238_in(4*N-1 downto 3*N),w7 => d238_in(3*N-1 downto 2*N),w8 => d238_in(2*N-1 downto N),w9 => d238_in(N-1 downto 0 ),d_out => d238_out,en_out =>open  ,sof_out=>open   );
CL239: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d239_in(9*N-1 downto 8*N),data2conv2 =>d239_in(8*N-1 downto 7*N),data2conv3 =>d239_in(7*N-1 downto 6*N),data2conv4 =>d239_in(6*N-1 downto 5*N),data2conv5 =>d239_in(5*N-1 downto 4*N),data2conv6 =>d239_in(4*N-1 downto 3*N),data2conv7 =>d239_in(3*N-1 downto 2*N),data2conv8 =>d239_in(2*N-1 downto N),data2conv9 =>d239_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d239_in(9*N-1 downto 8*N),w2 => d239_in(8*N-1 downto 7*N),w3 => d239_in(7*N-1 downto 6*N),w4 => d239_in(6*N-1 downto 5*N),w5 => d239_in(5*N-1 downto 4*N),w6 => d239_in(4*N-1 downto 3*N),w7 => d239_in(3*N-1 downto 2*N),w8 => d239_in(2*N-1 downto N),w9 => d239_in(N-1 downto 0 ),d_out => d239_out,en_out =>open  ,sof_out=>open   );
CL240: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d240_in(9*N-1 downto 8*N),data2conv2 =>d240_in(8*N-1 downto 7*N),data2conv3 =>d240_in(7*N-1 downto 6*N),data2conv4 =>d240_in(6*N-1 downto 5*N),data2conv5 =>d240_in(5*N-1 downto 4*N),data2conv6 =>d240_in(4*N-1 downto 3*N),data2conv7 =>d240_in(3*N-1 downto 2*N),data2conv8 =>d240_in(2*N-1 downto N),data2conv9 =>d240_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d240_in(9*N-1 downto 8*N),w2 => d240_in(8*N-1 downto 7*N),w3 => d240_in(7*N-1 downto 6*N),w4 => d240_in(6*N-1 downto 5*N),w5 => d240_in(5*N-1 downto 4*N),w6 => d240_in(4*N-1 downto 3*N),w7 => d240_in(3*N-1 downto 2*N),w8 => d240_in(2*N-1 downto N),w9 => d240_in(N-1 downto 0 ),d_out => d240_out,en_out =>open  ,sof_out=>open   );
CL241: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d241_in(9*N-1 downto 8*N),data2conv2 =>d241_in(8*N-1 downto 7*N),data2conv3 =>d241_in(7*N-1 downto 6*N),data2conv4 =>d241_in(6*N-1 downto 5*N),data2conv5 =>d241_in(5*N-1 downto 4*N),data2conv6 =>d241_in(4*N-1 downto 3*N),data2conv7 =>d241_in(3*N-1 downto 2*N),data2conv8 =>d241_in(2*N-1 downto N),data2conv9 =>d241_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d241_in(9*N-1 downto 8*N),w2 => d241_in(8*N-1 downto 7*N),w3 => d241_in(7*N-1 downto 6*N),w4 => d241_in(6*N-1 downto 5*N),w5 => d241_in(5*N-1 downto 4*N),w6 => d241_in(4*N-1 downto 3*N),w7 => d241_in(3*N-1 downto 2*N),w8 => d241_in(2*N-1 downto N),w9 => d241_in(N-1 downto 0 ),d_out => d241_out,en_out =>open  ,sof_out=>open   );
CL242: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d242_in(9*N-1 downto 8*N),data2conv2 =>d242_in(8*N-1 downto 7*N),data2conv3 =>d242_in(7*N-1 downto 6*N),data2conv4 =>d242_in(6*N-1 downto 5*N),data2conv5 =>d242_in(5*N-1 downto 4*N),data2conv6 =>d242_in(4*N-1 downto 3*N),data2conv7 =>d242_in(3*N-1 downto 2*N),data2conv8 =>d242_in(2*N-1 downto N),data2conv9 =>d242_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d242_in(9*N-1 downto 8*N),w2 => d242_in(8*N-1 downto 7*N),w3 => d242_in(7*N-1 downto 6*N),w4 => d242_in(6*N-1 downto 5*N),w5 => d242_in(5*N-1 downto 4*N),w6 => d242_in(4*N-1 downto 3*N),w7 => d242_in(3*N-1 downto 2*N),w8 => d242_in(2*N-1 downto N),w9 => d242_in(N-1 downto 0 ),d_out => d242_out,en_out =>open  ,sof_out=>open   );
CL243: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d243_in(9*N-1 downto 8*N),data2conv2 =>d243_in(8*N-1 downto 7*N),data2conv3 =>d243_in(7*N-1 downto 6*N),data2conv4 =>d243_in(6*N-1 downto 5*N),data2conv5 =>d243_in(5*N-1 downto 4*N),data2conv6 =>d243_in(4*N-1 downto 3*N),data2conv7 =>d243_in(3*N-1 downto 2*N),data2conv8 =>d243_in(2*N-1 downto N),data2conv9 =>d243_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d243_in(9*N-1 downto 8*N),w2 => d243_in(8*N-1 downto 7*N),w3 => d243_in(7*N-1 downto 6*N),w4 => d243_in(6*N-1 downto 5*N),w5 => d243_in(5*N-1 downto 4*N),w6 => d243_in(4*N-1 downto 3*N),w7 => d243_in(3*N-1 downto 2*N),w8 => d243_in(2*N-1 downto N),w9 => d243_in(N-1 downto 0 ),d_out => d243_out,en_out =>open  ,sof_out=>open   );
CL244: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d244_in(9*N-1 downto 8*N),data2conv2 =>d244_in(8*N-1 downto 7*N),data2conv3 =>d244_in(7*N-1 downto 6*N),data2conv4 =>d244_in(6*N-1 downto 5*N),data2conv5 =>d244_in(5*N-1 downto 4*N),data2conv6 =>d244_in(4*N-1 downto 3*N),data2conv7 =>d244_in(3*N-1 downto 2*N),data2conv8 =>d244_in(2*N-1 downto N),data2conv9 =>d244_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d244_in(9*N-1 downto 8*N),w2 => d244_in(8*N-1 downto 7*N),w3 => d244_in(7*N-1 downto 6*N),w4 => d244_in(6*N-1 downto 5*N),w5 => d244_in(5*N-1 downto 4*N),w6 => d244_in(4*N-1 downto 3*N),w7 => d244_in(3*N-1 downto 2*N),w8 => d244_in(2*N-1 downto N),w9 => d244_in(N-1 downto 0 ),d_out => d244_out,en_out =>open  ,sof_out=>open   );
CL245: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d245_in(9*N-1 downto 8*N),data2conv2 =>d245_in(8*N-1 downto 7*N),data2conv3 =>d245_in(7*N-1 downto 6*N),data2conv4 =>d245_in(6*N-1 downto 5*N),data2conv5 =>d245_in(5*N-1 downto 4*N),data2conv6 =>d245_in(4*N-1 downto 3*N),data2conv7 =>d245_in(3*N-1 downto 2*N),data2conv8 =>d245_in(2*N-1 downto N),data2conv9 =>d245_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d245_in(9*N-1 downto 8*N),w2 => d245_in(8*N-1 downto 7*N),w3 => d245_in(7*N-1 downto 6*N),w4 => d245_in(6*N-1 downto 5*N),w5 => d245_in(5*N-1 downto 4*N),w6 => d245_in(4*N-1 downto 3*N),w7 => d245_in(3*N-1 downto 2*N),w8 => d245_in(2*N-1 downto N),w9 => d245_in(N-1 downto 0 ),d_out => d245_out,en_out =>open  ,sof_out=>open   );
CL246: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d246_in(9*N-1 downto 8*N),data2conv2 =>d246_in(8*N-1 downto 7*N),data2conv3 =>d246_in(7*N-1 downto 6*N),data2conv4 =>d246_in(6*N-1 downto 5*N),data2conv5 =>d246_in(5*N-1 downto 4*N),data2conv6 =>d246_in(4*N-1 downto 3*N),data2conv7 =>d246_in(3*N-1 downto 2*N),data2conv8 =>d246_in(2*N-1 downto N),data2conv9 =>d246_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d246_in(9*N-1 downto 8*N),w2 => d246_in(8*N-1 downto 7*N),w3 => d246_in(7*N-1 downto 6*N),w4 => d246_in(6*N-1 downto 5*N),w5 => d246_in(5*N-1 downto 4*N),w6 => d246_in(4*N-1 downto 3*N),w7 => d246_in(3*N-1 downto 2*N),w8 => d246_in(2*N-1 downto N),w9 => d246_in(N-1 downto 0 ),d_out => d246_out,en_out =>open  ,sof_out=>open   );
CL247: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d247_in(9*N-1 downto 8*N),data2conv2 =>d247_in(8*N-1 downto 7*N),data2conv3 =>d247_in(7*N-1 downto 6*N),data2conv4 =>d247_in(6*N-1 downto 5*N),data2conv5 =>d247_in(5*N-1 downto 4*N),data2conv6 =>d247_in(4*N-1 downto 3*N),data2conv7 =>d247_in(3*N-1 downto 2*N),data2conv8 =>d247_in(2*N-1 downto N),data2conv9 =>d247_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d247_in(9*N-1 downto 8*N),w2 => d247_in(8*N-1 downto 7*N),w3 => d247_in(7*N-1 downto 6*N),w4 => d247_in(6*N-1 downto 5*N),w5 => d247_in(5*N-1 downto 4*N),w6 => d247_in(4*N-1 downto 3*N),w7 => d247_in(3*N-1 downto 2*N),w8 => d247_in(2*N-1 downto N),w9 => d247_in(N-1 downto 0 ),d_out => d247_out,en_out =>open  ,sof_out=>open   );
CL248: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d248_in(9*N-1 downto 8*N),data2conv2 =>d248_in(8*N-1 downto 7*N),data2conv3 =>d248_in(7*N-1 downto 6*N),data2conv4 =>d248_in(6*N-1 downto 5*N),data2conv5 =>d248_in(5*N-1 downto 4*N),data2conv6 =>d248_in(4*N-1 downto 3*N),data2conv7 =>d248_in(3*N-1 downto 2*N),data2conv8 =>d248_in(2*N-1 downto N),data2conv9 =>d248_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d248_in(9*N-1 downto 8*N),w2 => d248_in(8*N-1 downto 7*N),w3 => d248_in(7*N-1 downto 6*N),w4 => d248_in(6*N-1 downto 5*N),w5 => d248_in(5*N-1 downto 4*N),w6 => d248_in(4*N-1 downto 3*N),w7 => d248_in(3*N-1 downto 2*N),w8 => d248_in(2*N-1 downto N),w9 => d248_in(N-1 downto 0 ),d_out => d248_out,en_out =>open  ,sof_out=>open   );
CL249: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d249_in(9*N-1 downto 8*N),data2conv2 =>d249_in(8*N-1 downto 7*N),data2conv3 =>d249_in(7*N-1 downto 6*N),data2conv4 =>d249_in(6*N-1 downto 5*N),data2conv5 =>d249_in(5*N-1 downto 4*N),data2conv6 =>d249_in(4*N-1 downto 3*N),data2conv7 =>d249_in(3*N-1 downto 2*N),data2conv8 =>d249_in(2*N-1 downto N),data2conv9 =>d249_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d249_in(9*N-1 downto 8*N),w2 => d249_in(8*N-1 downto 7*N),w3 => d249_in(7*N-1 downto 6*N),w4 => d249_in(6*N-1 downto 5*N),w5 => d249_in(5*N-1 downto 4*N),w6 => d249_in(4*N-1 downto 3*N),w7 => d249_in(3*N-1 downto 2*N),w8 => d249_in(2*N-1 downto N),w9 => d249_in(N-1 downto 0 ),d_out => d249_out,en_out =>open  ,sof_out=>open   );
CL250: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d250_in(9*N-1 downto 8*N),data2conv2 =>d250_in(8*N-1 downto 7*N),data2conv3 =>d250_in(7*N-1 downto 6*N),data2conv4 =>d250_in(6*N-1 downto 5*N),data2conv5 =>d250_in(5*N-1 downto 4*N),data2conv6 =>d250_in(4*N-1 downto 3*N),data2conv7 =>d250_in(3*N-1 downto 2*N),data2conv8 =>d250_in(2*N-1 downto N),data2conv9 =>d250_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d250_in(9*N-1 downto 8*N),w2 => d250_in(8*N-1 downto 7*N),w3 => d250_in(7*N-1 downto 6*N),w4 => d250_in(6*N-1 downto 5*N),w5 => d250_in(5*N-1 downto 4*N),w6 => d250_in(4*N-1 downto 3*N),w7 => d250_in(3*N-1 downto 2*N),w8 => d250_in(2*N-1 downto N),w9 => d250_in(N-1 downto 0 ),d_out => d250_out,en_out =>open  ,sof_out=>open   );
CL251: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d251_in(9*N-1 downto 8*N),data2conv2 =>d251_in(8*N-1 downto 7*N),data2conv3 =>d251_in(7*N-1 downto 6*N),data2conv4 =>d251_in(6*N-1 downto 5*N),data2conv5 =>d251_in(5*N-1 downto 4*N),data2conv6 =>d251_in(4*N-1 downto 3*N),data2conv7 =>d251_in(3*N-1 downto 2*N),data2conv8 =>d251_in(2*N-1 downto N),data2conv9 =>d251_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d251_in(9*N-1 downto 8*N),w2 => d251_in(8*N-1 downto 7*N),w3 => d251_in(7*N-1 downto 6*N),w4 => d251_in(6*N-1 downto 5*N),w5 => d251_in(5*N-1 downto 4*N),w6 => d251_in(4*N-1 downto 3*N),w7 => d251_in(3*N-1 downto 2*N),w8 => d251_in(2*N-1 downto N),w9 => d251_in(N-1 downto 0 ),d_out => d251_out,en_out =>open  ,sof_out=>open   );
CL252: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d252_in(9*N-1 downto 8*N),data2conv2 =>d252_in(8*N-1 downto 7*N),data2conv3 =>d252_in(7*N-1 downto 6*N),data2conv4 =>d252_in(6*N-1 downto 5*N),data2conv5 =>d252_in(5*N-1 downto 4*N),data2conv6 =>d252_in(4*N-1 downto 3*N),data2conv7 =>d252_in(3*N-1 downto 2*N),data2conv8 =>d252_in(2*N-1 downto N),data2conv9 =>d252_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d252_in(9*N-1 downto 8*N),w2 => d252_in(8*N-1 downto 7*N),w3 => d252_in(7*N-1 downto 6*N),w4 => d252_in(6*N-1 downto 5*N),w5 => d252_in(5*N-1 downto 4*N),w6 => d252_in(4*N-1 downto 3*N),w7 => d252_in(3*N-1 downto 2*N),w8 => d252_in(2*N-1 downto N),w9 => d252_in(N-1 downto 0 ),d_out => d252_out,en_out =>open  ,sof_out=>open   );
CL253: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d253_in(9*N-1 downto 8*N),data2conv2 =>d253_in(8*N-1 downto 7*N),data2conv3 =>d253_in(7*N-1 downto 6*N),data2conv4 =>d253_in(6*N-1 downto 5*N),data2conv5 =>d253_in(5*N-1 downto 4*N),data2conv6 =>d253_in(4*N-1 downto 3*N),data2conv7 =>d253_in(3*N-1 downto 2*N),data2conv8 =>d253_in(2*N-1 downto N),data2conv9 =>d253_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d253_in(9*N-1 downto 8*N),w2 => d253_in(8*N-1 downto 7*N),w3 => d253_in(7*N-1 downto 6*N),w4 => d253_in(6*N-1 downto 5*N),w5 => d253_in(5*N-1 downto 4*N),w6 => d253_in(4*N-1 downto 3*N),w7 => d253_in(3*N-1 downto 2*N),w8 => d253_in(2*N-1 downto N),w9 => d253_in(N-1 downto 0 ),d_out => d253_out,en_out =>open  ,sof_out=>open   );
CL254: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d254_in(9*N-1 downto 8*N),data2conv2 =>d254_in(8*N-1 downto 7*N),data2conv3 =>d254_in(7*N-1 downto 6*N),data2conv4 =>d254_in(6*N-1 downto 5*N),data2conv5 =>d254_in(5*N-1 downto 4*N),data2conv6 =>d254_in(4*N-1 downto 3*N),data2conv7 =>d254_in(3*N-1 downto 2*N),data2conv8 =>d254_in(2*N-1 downto N),data2conv9 =>d254_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d254_in(9*N-1 downto 8*N),w2 => d254_in(8*N-1 downto 7*N),w3 => d254_in(7*N-1 downto 6*N),w4 => d254_in(6*N-1 downto 5*N),w5 => d254_in(5*N-1 downto 4*N),w6 => d254_in(4*N-1 downto 3*N),w7 => d254_in(3*N-1 downto 2*N),w8 => d254_in(2*N-1 downto N),w9 => d254_in(N-1 downto 0 ),d_out => d254_out,en_out =>open  ,sof_out=>open   );
CL255: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d255_in(9*N-1 downto 8*N),data2conv2 =>d255_in(8*N-1 downto 7*N),data2conv3 =>d255_in(7*N-1 downto 6*N),data2conv4 =>d255_in(6*N-1 downto 5*N),data2conv5 =>d255_in(5*N-1 downto 4*N),data2conv6 =>d255_in(4*N-1 downto 3*N),data2conv7 =>d255_in(3*N-1 downto 2*N),data2conv8 =>d255_in(2*N-1 downto N),data2conv9 =>d255_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d255_in(9*N-1 downto 8*N),w2 => d255_in(8*N-1 downto 7*N),w3 => d255_in(7*N-1 downto 6*N),w4 => d255_in(6*N-1 downto 5*N),w5 => d255_in(5*N-1 downto 4*N),w6 => d255_in(4*N-1 downto 3*N),w7 => d255_in(3*N-1 downto 2*N),w8 => d255_in(2*N-1 downto N),w9 => d255_in(N-1 downto 0 ),d_out => d255_out,en_out =>open  ,sof_out=>open   );
CL256: ConvLayer1 generic map (mult_sum=>mult_sum,N=>N,M=>M,W=>W,SR=>SR) port map(clk=>clk,rst=>rst,data2conv1 =>d256_in(9*N-1 downto 8*N),data2conv2 =>d256_in(8*N-1 downto 7*N),data2conv3 =>d256_in(7*N-1 downto 6*N),data2conv4 =>d256_in(6*N-1 downto 5*N),data2conv5 =>d256_in(5*N-1 downto 4*N),data2conv6 =>d256_in(4*N-1 downto 3*N),data2conv7 =>d256_in(3*N-1 downto 2*N),data2conv8 =>d256_in(2*N-1 downto N),data2conv9 =>d256_in(N-1 downto 0 ),en_in =>en_in,sof_in =>sof_in,w1 => d256_in(9*N-1 downto 8*N),w2 => d256_in(8*N-1 downto 7*N),w3 => d256_in(7*N-1 downto 6*N),w4 => d256_in(6*N-1 downto 5*N),w5 => d256_in(5*N-1 downto 4*N),w6 => d256_in(4*N-1 downto 3*N),w7 => d256_in(3*N-1 downto 2*N),w8 => d256_in(2*N-1 downto N),w9 => d256_in(N-1 downto 0 ),d_out => d256_out,en_out =>open  ,sof_out=>open   );

  p_sums: process (clk)
  begin
    if rising_edge(clk) then
       sum1  <= (d01_out(d01_out'left) & d01_out(d01_out'left) & d01_out) +  (d02_out(d02_out'left) & d02_out(d02_out'left) & d02_out) + (d03_out(d03_out'left) & d03_out(d03_out'left) & d03_out) +  (d03_out(d03_out'left) & d03_out(d03_out'left) & d03_out);  
       sum2  <= (d05_out(d05_out'left) & d05_out(d05_out'left) & d05_out) +  (d06_out(d06_out'left) & d06_out(d06_out'left) & d06_out) + (d07_out(d07_out'left) & d07_out(d07_out'left) & d07_out) +  (d07_out(d07_out'left) & d07_out(d07_out'left) & d07_out);  
       sum3  <= (d09_out(d09_out'left) & d09_out(d09_out'left) & d09_out) +  (d10_out(d10_out'left) & d10_out(d10_out'left) & d10_out) + (d11_out(d11_out'left) & d11_out(d11_out'left) & d11_out) +  (d11_out(d11_out'left) & d11_out(d11_out'left) & d11_out);  
       sum4  <= (d13_out(d13_out'left) & d13_out(d13_out'left) & d13_out) +  (d14_out(d14_out'left) & d14_out(d14_out'left) & d14_out) + (d15_out(d15_out'left) & d15_out(d15_out'left) & d15_out) +  (d15_out(d15_out'left) & d15_out(d15_out'left) & d15_out);  
       sum5  <= (d17_out(d17_out'left) & d17_out(d17_out'left) & d17_out) +  (d18_out(d18_out'left) & d18_out(d18_out'left) & d18_out) + (d19_out(d19_out'left) & d19_out(d19_out'left) & d19_out) +  (d19_out(d19_out'left) & d19_out(d19_out'left) & d19_out);  
       sum6  <= (d21_out(d21_out'left) & d21_out(d21_out'left) & d21_out) +  (d22_out(d22_out'left) & d22_out(d22_out'left) & d22_out) + (d23_out(d23_out'left) & d23_out(d23_out'left) & d23_out) +  (d23_out(d23_out'left) & d23_out(d23_out'left) & d23_out);  
       sum7  <= (d25_out(d25_out'left) & d25_out(d25_out'left) & d25_out) +  (d26_out(d26_out'left) & d26_out(d26_out'left) & d26_out) + (d27_out(d27_out'left) & d27_out(d27_out'left) & d27_out) +  (d27_out(d27_out'left) & d27_out(d27_out'left) & d27_out);  
       sum8  <= (d29_out(d29_out'left) & d29_out(d29_out'left) & d29_out) +  (d30_out(d30_out'left) & d30_out(d30_out'left) & d30_out) + (d31_out(d31_out'left) & d31_out(d31_out'left) & d31_out) +  (d31_out(d31_out'left) & d31_out(d31_out'left) & d31_out);  
       sum9  <= (d33_out(d33_out'left) & d33_out(d33_out'left) & d33_out) +  (d34_out(d34_out'left) & d34_out(d34_out'left) & d34_out) + (d35_out(d35_out'left) & d35_out(d35_out'left) & d35_out) +  (d35_out(d35_out'left) & d35_out(d35_out'left) & d35_out);  
       sum10 <= (d37_out(d37_out'left) & d37_out(d37_out'left) & d37_out) +  (d38_out(d38_out'left) & d38_out(d38_out'left) & d38_out) + (d39_out(d39_out'left) & d39_out(d39_out'left) & d39_out) +  (d39_out(d39_out'left) & d39_out(d39_out'left) & d39_out);  
       sum11 <= (d41_out(d41_out'left) & d41_out(d41_out'left) & d41_out) +  (d42_out(d42_out'left) & d42_out(d42_out'left) & d42_out) + (d43_out(d43_out'left) & d43_out(d43_out'left) & d43_out) +  (d43_out(d43_out'left) & d43_out(d43_out'left) & d43_out);  
       sum12 <= (d45_out(d45_out'left) & d45_out(d45_out'left) & d45_out) +  (d46_out(d46_out'left) & d46_out(d46_out'left) & d46_out) + (d47_out(d47_out'left) & d47_out(d47_out'left) & d47_out) +  (d47_out(d47_out'left) & d47_out(d47_out'left) & d47_out);  
       sum13 <= (d49_out(d49_out'left) & d49_out(d49_out'left) & d49_out) +  (d50_out(d50_out'left) & d50_out(d50_out'left) & d50_out) + (d51_out(d51_out'left) & d51_out(d51_out'left) & d51_out) +  (d51_out(d51_out'left) & d51_out(d51_out'left) & d51_out);  
       sum14 <= (d53_out(d53_out'left) & d53_out(d53_out'left) & d53_out) +  (d54_out(d54_out'left) & d54_out(d54_out'left) & d54_out) + (d55_out(d55_out'left) & d55_out(d55_out'left) & d55_out) +  (d55_out(d55_out'left) & d55_out(d55_out'left) & d55_out);  
       sum15 <= (d57_out(d57_out'left) & d57_out(d57_out'left) & d57_out) +  (d58_out(d58_out'left) & d58_out(d58_out'left) & d58_out) + (d59_out(d59_out'left) & d59_out(d59_out'left) & d59_out) +  (d59_out(d59_out'left) & d59_out(d59_out'left) & d59_out);  
       sum16 <= (d61_out(d61_out'left) & d61_out(d61_out'left) & d61_out) +  (d62_out(d62_out'left) & d62_out(d62_out'left) & d62_out) + (d63_out(d63_out'left) & d63_out(d63_out'left) & d63_out) +  (d63_out(d63_out'left) & d63_out(d63_out'left) & d63_out);  
       sum22 <= (d65_out (d65_out 'left) & d65_out (d65_out 'left) & d65_out ) + (d66_out (d66_out 'left) & d66_out (d66_out 'left) & d66_out ) + (d67_out (d67_out 'left) & d67_out (d67_out 'left) & d67_out ) + (d68_out (d68_out 'left) & d68_out (d68_out 'left) & d68_out );
       sum23 <= (d69_out (d69_out 'left) & d69_out (d69_out 'left) & d69_out ) + (d70_out (d70_out 'left) & d70_out (d70_out 'left) & d70_out ) + (d71_out (d71_out 'left) & d71_out (d71_out 'left) & d71_out ) + (d72_out (d72_out 'left) & d72_out (d72_out 'left) & d72_out );
       sum24 <= (d73_out (d73_out 'left) & d73_out (d73_out 'left) & d73_out ) + (d74_out (d74_out 'left) & d74_out (d74_out 'left) & d74_out ) + (d75_out (d75_out 'left) & d75_out (d75_out 'left) & d75_out ) + (d76_out (d76_out 'left) & d76_out (d76_out 'left) & d76_out );
       sum25 <= (d77_out (d77_out 'left) & d77_out (d77_out 'left) & d77_out ) + (d78_out (d78_out 'left) & d78_out (d78_out 'left) & d78_out ) + (d79_out (d79_out 'left) & d79_out (d79_out 'left) & d79_out ) + (d80_out (d80_out 'left) & d80_out (d80_out 'left) & d80_out );
       sum26 <= (d81_out (d81_out 'left) & d81_out (d81_out 'left) & d81_out ) + (d82_out (d82_out 'left) & d82_out (d82_out 'left) & d82_out ) + (d83_out (d83_out 'left) & d83_out (d83_out 'left) & d83_out ) + (d84_out (d84_out 'left) & d84_out (d84_out 'left) & d84_out );
       sum27 <= (d85_out (d85_out 'left) & d85_out (d85_out 'left) & d85_out ) + (d86_out (d86_out 'left) & d86_out (d86_out 'left) & d86_out ) + (d87_out (d87_out 'left) & d87_out (d87_out 'left) & d87_out ) + (d88_out (d88_out 'left) & d88_out (d88_out 'left) & d88_out );
       sum28 <= (d89_out (d89_out 'left) & d89_out (d89_out 'left) & d89_out ) + (d90_out (d90_out 'left) & d90_out (d90_out 'left) & d90_out ) + (d91_out (d91_out 'left) & d91_out (d91_out 'left) & d91_out ) + (d92_out (d92_out 'left) & d92_out (d92_out 'left) & d92_out );
       sum29 <= (d93_out (d93_out 'left) & d93_out (d93_out 'left) & d93_out ) + (d94_out (d94_out 'left) & d94_out (d94_out 'left) & d94_out ) + (d95_out (d95_out 'left) & d95_out (d95_out 'left) & d95_out ) + (d96_out (d96_out 'left) & d96_out (d96_out 'left) & d96_out );
       sum30 <= (d97_out (d97_out 'left) & d97_out (d97_out 'left) & d97_out ) + (d98_out (d98_out 'left) & d98_out (d98_out 'left) & d98_out ) + (d99_out (d99_out 'left) & d99_out (d99_out 'left) & d99_out ) + (d100_out(d100_out'left) & d100_out(d100_out'left) & d100_out);
       sum31 <= (d101_out(d101_out'left) & d101_out(d101_out'left) & d101_out) + (d102_out(d102_out'left) & d102_out(d102_out'left) & d102_out) + (d103_out(d103_out'left) & d103_out(d103_out'left) & d103_out) + (d104_out(d104_out'left) & d104_out(d104_out'left) & d104_out);
       sum32 <= (d105_out(d105_out'left) & d105_out(d105_out'left) & d105_out) + (d106_out(d106_out'left) & d106_out(d106_out'left) & d106_out) + (d107_out(d107_out'left) & d107_out(d107_out'left) & d107_out) + (d108_out(d108_out'left) & d108_out(d108_out'left) & d108_out);
       sum33 <= (d109_out(d109_out'left) & d109_out(d109_out'left) & d109_out) + (d110_out(d110_out'left) & d110_out(d110_out'left) & d110_out) + (d111_out(d111_out'left) & d111_out(d111_out'left) & d111_out) + (d112_out(d112_out'left) & d112_out(d112_out'left) & d112_out);
       sum34 <= (d113_out(d113_out'left) & d113_out(d113_out'left) & d113_out) + (d114_out(d114_out'left) & d114_out(d114_out'left) & d114_out) + (d115_out(d115_out'left) & d115_out(d115_out'left) & d115_out) + (d116_out(d116_out'left) & d116_out(d116_out'left) & d116_out);
       sum35 <= (d117_out(d117_out'left) & d117_out(d117_out'left) & d117_out) + (d118_out(d118_out'left) & d118_out(d118_out'left) & d118_out) + (d119_out(d119_out'left) & d119_out(d119_out'left) & d119_out) + (d120_out(d120_out'left) & d120_out(d120_out'left) & d120_out);
       sum36 <= (d121_out(d121_out'left) & d121_out(d121_out'left) & d121_out) + (d122_out(d122_out'left) & d122_out(d122_out'left) & d122_out) + (d123_out(d123_out'left) & d123_out(d123_out'left) & d123_out) + (d124_out(d124_out'left) & d124_out(d124_out'left) & d124_out);
       sum37 <= (d125_out(d125_out'left) & d125_out(d125_out'left) & d125_out) + (d126_out(d126_out'left) & d126_out(d126_out'left) & d126_out) + (d127_out(d127_out'left) & d127_out(d127_out'left) & d127_out) + (d128_out(d128_out'left) & d128_out(d128_out'left) & d128_out);

       sum44 <= (d129_out(d129_out'left) & d129_out(d129_out'left) & d129_out) + (d130_out(d130_out'left) & d130_out(d130_out'left) & d130_out) + (d131_out(d131_out'left) & d131_out(d131_out'left) & d131_out) + (d132_out(d132_out'left) & d132_out(d132_out'left) & d132_out);
       sum45 <= (d133_out(d133_out'left) & d133_out(d133_out'left) & d133_out) + (d134_out(d134_out'left) & d134_out(d134_out'left) & d134_out) + (d135_out(d135_out'left) & d135_out(d135_out'left) & d135_out) + (d136_out(d136_out'left) & d136_out(d136_out'left) & d136_out);
       sum46 <= (d137_out(d137_out'left) & d137_out(d137_out'left) & d137_out) + (d138_out(d138_out'left) & d138_out(d138_out'left) & d138_out) + (d139_out(d139_out'left) & d139_out(d139_out'left) & d139_out) + (d140_out(d140_out'left) & d140_out(d140_out'left) & d140_out);
       sum47 <= (d141_out(d141_out'left) & d141_out(d141_out'left) & d141_out) + (d142_out(d142_out'left) & d142_out(d142_out'left) & d142_out) + (d143_out(d143_out'left) & d143_out(d143_out'left) & d143_out) + (d144_out(d144_out'left) & d144_out(d144_out'left) & d144_out);
       sum48 <= (d145_out(d145_out'left) & d145_out(d145_out'left) & d145_out) + (d146_out(d146_out'left) & d146_out(d146_out'left) & d146_out) + (d147_out(d147_out'left) & d147_out(d147_out'left) & d147_out) + (d148_out(d148_out'left) & d148_out(d148_out'left) & d148_out);
       sum49 <= (d149_out(d149_out'left) & d149_out(d149_out'left) & d149_out) + (d150_out(d150_out'left) & d150_out(d150_out'left) & d150_out) + (d151_out(d151_out'left) & d151_out(d151_out'left) & d151_out) + (d152_out(d152_out'left) & d152_out(d152_out'left) & d152_out);
       sum50 <= (d153_out(d153_out'left) & d153_out(d153_out'left) & d153_out) + (d154_out(d154_out'left) & d154_out(d154_out'left) & d154_out) + (d155_out(d155_out'left) & d155_out(d155_out'left) & d155_out) + (d156_out(d156_out'left) & d156_out(d156_out'left) & d156_out);
       sum51 <= (d157_out(d157_out'left) & d157_out(d157_out'left) & d157_out) + (d158_out(d158_out'left) & d158_out(d158_out'left) & d158_out) + (d159_out(d159_out'left) & d159_out(d159_out'left) & d159_out) + (d160_out(d160_out'left) & d160_out(d160_out'left) & d160_out);
       sum52 <= (d161_out(d161_out'left) & d161_out(d161_out'left) & d161_out) + (d162_out(d162_out'left) & d162_out(d162_out'left) & d162_out) + (d163_out(d163_out'left) & d163_out(d163_out'left) & d163_out) + (d164_out(d164_out'left) & d164_out(d164_out'left) & d164_out);
       sum53 <= (d165_out(d165_out'left) & d165_out(d165_out'left) & d165_out) + (d166_out(d166_out'left) & d166_out(d166_out'left) & d166_out) + (d167_out(d167_out'left) & d167_out(d167_out'left) & d167_out) + (d168_out(d168_out'left) & d168_out(d168_out'left) & d168_out);
       sum54 <= (d169_out(d169_out'left) & d169_out(d169_out'left) & d169_out) + (d170_out(d170_out'left) & d170_out(d170_out'left) & d170_out) + (d171_out(d171_out'left) & d171_out(d171_out'left) & d171_out) + (d172_out(d172_out'left) & d172_out(d172_out'left) & d172_out);
       sum55 <= (d173_out(d173_out'left) & d173_out(d173_out'left) & d173_out) + (d174_out(d174_out'left) & d174_out(d174_out'left) & d174_out) + (d175_out(d175_out'left) & d175_out(d175_out'left) & d175_out) + (d176_out(d176_out'left) & d176_out(d176_out'left) & d176_out);
       sum56 <= (d177_out(d177_out'left) & d177_out(d177_out'left) & d177_out) + (d178_out(d178_out'left) & d178_out(d178_out'left) & d178_out) + (d179_out(d179_out'left) & d179_out(d179_out'left) & d179_out) + (d180_out(d180_out'left) & d180_out(d180_out'left) & d180_out);
       sum57 <= (d181_out(d181_out'left) & d181_out(d181_out'left) & d181_out) + (d182_out(d182_out'left) & d182_out(d182_out'left) & d182_out) + (d183_out(d183_out'left) & d183_out(d183_out'left) & d183_out) + (d184_out(d184_out'left) & d184_out(d184_out'left) & d184_out);
       sum58 <= (d185_out(d185_out'left) & d185_out(d185_out'left) & d185_out) + (d186_out(d186_out'left) & d186_out(d186_out'left) & d186_out) + (d187_out(d187_out'left) & d187_out(d187_out'left) & d187_out) + (d188_out(d188_out'left) & d188_out(d188_out'left) & d188_out);
       sum59 <= (d189_out(d189_out'left) & d189_out(d189_out'left) & d189_out) + (d190_out(d190_out'left) & d190_out(d190_out'left) & d190_out) + (d191_out(d191_out'left) & d191_out(d191_out'left) & d191_out) + (d192_out(d192_out'left) & d192_out(d192_out'left) & d192_out);
       sum60 <= (d193_out(d193_out'left) & d193_out(d193_out'left) & d193_out) + (d194_out(d194_out'left) & d194_out(d194_out'left) & d194_out) + (d195_out(d195_out'left) & d195_out(d195_out'left) & d195_out) + (d196_out(d196_out'left) & d196_out(d196_out'left) & d196_out);
       sum61 <= (d197_out(d197_out'left) & d197_out(d197_out'left) & d197_out) + (d198_out(d198_out'left) & d198_out(d198_out'left) & d198_out) + (d199_out(d199_out'left) & d199_out(d199_out'left) & d199_out) + (d200_out(d200_out'left) & d200_out(d200_out'left) & d200_out);
       sum62 <= (d201_out(d201_out'left) & d201_out(d201_out'left) & d201_out) + (d202_out(d202_out'left) & d202_out(d202_out'left) & d202_out) + (d203_out(d203_out'left) & d203_out(d203_out'left) & d203_out) + (d204_out(d204_out'left) & d204_out(d204_out'left) & d204_out);
       sum63 <= (d205_out(d205_out'left) & d205_out(d205_out'left) & d205_out) + (d206_out(d206_out'left) & d206_out(d206_out'left) & d206_out) + (d207_out(d207_out'left) & d207_out(d207_out'left) & d207_out) + (d208_out(d208_out'left) & d208_out(d208_out'left) & d208_out);
       sum64 <= (d209_out(d209_out'left) & d209_out(d209_out'left) & d209_out) + (d210_out(d210_out'left) & d210_out(d210_out'left) & d210_out) + (d211_out(d211_out'left) & d211_out(d211_out'left) & d211_out) + (d212_out(d212_out'left) & d212_out(d212_out'left) & d212_out);
       sum65 <= (d213_out(d213_out'left) & d213_out(d213_out'left) & d213_out) + (d214_out(d214_out'left) & d214_out(d214_out'left) & d214_out) + (d215_out(d215_out'left) & d215_out(d215_out'left) & d215_out) + (d216_out(d216_out'left) & d216_out(d216_out'left) & d216_out);
       sum66 <= (d217_out(d217_out'left) & d217_out(d217_out'left) & d217_out) + (d218_out(d218_out'left) & d218_out(d218_out'left) & d218_out) + (d219_out(d219_out'left) & d219_out(d219_out'left) & d219_out) + (d220_out(d220_out'left) & d220_out(d220_out'left) & d220_out);
       sum67 <= (d221_out(d221_out'left) & d221_out(d221_out'left) & d221_out) + (d222_out(d222_out'left) & d222_out(d222_out'left) & d222_out) + (d223_out(d223_out'left) & d223_out(d223_out'left) & d223_out) + (d224_out(d224_out'left) & d224_out(d224_out'left) & d224_out);
       sum68 <= (d225_out(d225_out'left) & d225_out(d225_out'left) & d225_out) + (d226_out(d226_out'left) & d226_out(d226_out'left) & d226_out) + (d227_out(d227_out'left) & d227_out(d227_out'left) & d227_out) + (d228_out(d228_out'left) & d228_out(d228_out'left) & d228_out);
       sum69 <= (d229_out(d229_out'left) & d229_out(d229_out'left) & d229_out) + (d230_out(d230_out'left) & d230_out(d230_out'left) & d230_out) + (d231_out(d231_out'left) & d231_out(d231_out'left) & d231_out) + (d232_out(d232_out'left) & d232_out(d232_out'left) & d232_out);
       sum70 <= (d233_out(d233_out'left) & d233_out(d233_out'left) & d233_out) + (d234_out(d234_out'left) & d234_out(d234_out'left) & d234_out) + (d235_out(d235_out'left) & d235_out(d235_out'left) & d235_out) + (d236_out(d236_out'left) & d236_out(d236_out'left) & d236_out);
       sum71 <= (d237_out(d237_out'left) & d237_out(d237_out'left) & d237_out) + (d238_out(d238_out'left) & d238_out(d238_out'left) & d238_out) + (d239_out(d239_out'left) & d239_out(d239_out'left) & d239_out) + (d240_out(d240_out'left) & d240_out(d240_out'left) & d240_out);
       sum72 <= (d241_out(d241_out'left) & d241_out(d241_out'left) & d241_out) + (d242_out(d242_out'left) & d242_out(d242_out'left) & d242_out) + (d243_out(d243_out'left) & d243_out(d243_out'left) & d243_out) + (d244_out(d244_out'left) & d244_out(d244_out'left) & d244_out);
       sum73 <= (d245_out(d245_out'left) & d245_out(d245_out'left) & d245_out) + (d246_out(d246_out'left) & d246_out(d246_out'left) & d246_out) + (d247_out(d247_out'left) & d247_out(d247_out'left) & d247_out) + (d248_out(d248_out'left) & d248_out(d248_out'left) & d248_out);
       sum74 <= (d249_out(d249_out'left) & d249_out(d249_out'left) & d249_out) + (d250_out(d250_out'left) & d250_out(d250_out'left) & d250_out) + (d251_out(d251_out'left) & d251_out(d251_out'left) & d251_out) + (d252_out(d252_out'left) & d252_out(d252_out'left) & d252_out);
       sum75 <= (d253_out(d253_out'left) & d253_out(d253_out'left) & d253_out) + (d254_out(d254_out'left) & d254_out(d254_out'left) & d254_out) + (d255_out(d255_out'left) & d255_out(d255_out'left) & d255_out) + (d256_out(d256_out'left) & d256_out(d256_out'left) & d256_out);

       sum17 <= (sum1(sum1  'left) & sum1(sum1  'left) & sum1 ) + (sum2(sum2  'left) & sum2(sum2  'left) & sum2 ) + (sum3(sum3  'left) & sum3(sum3  'left) & sum3 ) + (sum4(sum4  'left) & sum4(sum4  'left) & sum4 );  
       sum18 <= (sum5(sum5  'left) & sum5(sum5  'left) & sum5 ) + (sum6(sum6  'left) & sum6(sum6  'left) & sum6 ) + (sum7(sum7  'left) & sum7(sum7  'left) & sum7 ) + (sum8(sum8  'left) & sum8(sum8  'left) & sum8 );  
       sum19 <= (sum9(sum9  'left) & sum9(sum9  'left) & sum9 ) + (sum10(sum10'left) & sum10(sum10'left) & sum10) + (sum11(sum11'left) & sum11(sum11'left) & sum11) + (sum12(sum12'left) & sum12(sum12'left) & sum12);
       sum20 <= (sum13(sum13'left) & sum13(sum13'left) & sum13) + (sum14(sum14'left) & sum14(sum14'left) & sum14) + (sum15(sum15'left) & sum15(sum15'left) & sum15) + (sum16(sum16'left) & sum16(sum16'left) & sum16);
       sum38 <= (sum22(sum22'left) & sum22(sum22'left) & sum22) + (sum23(sum23'left) & sum23(sum23'left) & sum23) + (sum24(sum24'left) & sum24(sum24'left) & sum24) + (sum25(sum25'left) & sum25(sum25'left) & sum25);
       sum39 <= (sum26(sum26'left) & sum26(sum26'left) & sum26) + (sum27(sum27'left) & sum27(sum27'left) & sum27) + (sum28(sum28'left) & sum28(sum28'left) & sum28) + (sum29(sum29'left) & sum29(sum29'left) & sum29);
       sum40 <= (sum30(sum30'left) & sum30(sum30'left) & sum30) + (sum31(sum31'left) & sum31(sum31'left) & sum31) + (sum32(sum32'left) & sum32(sum32'left) & sum32) + (sum33(sum33'left) & sum33(sum33'left) & sum33);
       sum41 <= (sum34(sum34'left) & sum34(sum34'left) & sum34) + (sum35(sum35'left) & sum35(sum35'left) & sum35) + (sum36(sum36'left) & sum36(sum36'left) & sum36) + (sum37(sum37'left) & sum37(sum37'left) & sum37);

       sum76 <= (sum44(sum44'left) & sum44(sum44'left) & sum44) + (sum45(sum45'left) & sum45(sum45'left) & sum45) + (sum46(sum46'left) & sum46(sum46'left) & sum46) + (sum47(sum47'left) & sum47(sum47'left) & sum47);
       sum77 <= (sum48(sum48'left) & sum48(sum48'left) & sum48) + (sum49(sum49'left) & sum49(sum49'left) & sum49) + (sum50(sum50'left) & sum50(sum50'left) & sum50) + (sum51(sum51'left) & sum51(sum51'left) & sum51);
       sum78 <= (sum52(sum52'left) & sum52(sum52'left) & sum52) + (sum53(sum53'left) & sum53(sum53'left) & sum53) + (sum54(sum54'left) & sum54(sum54'left) & sum54) + (sum55(sum55'left) & sum55(sum55'left) & sum55);
       sum79 <= (sum56(sum56'left) & sum56(sum56'left) & sum56) + (sum57(sum57'left) & sum57(sum57'left) & sum57) + (sum58(sum58'left) & sum58(sum58'left) & sum58) + (sum59(sum59'left) & sum59(sum59'left) & sum59);
       sum80 <= (sum60(sum60'left) & sum60(sum60'left) & sum60) + (sum61(sum61'left) & sum61(sum61'left) & sum61) + (sum62(sum62'left) & sum62(sum62'left) & sum62) + (sum63(sum63'left) & sum63(sum63'left) & sum63);
       sum81 <= (sum64(sum64'left) & sum64(sum64'left) & sum64) + (sum65(sum65'left) & sum65(sum65'left) & sum65) + (sum66(sum66'left) & sum66(sum66'left) & sum66) + (sum67(sum67'left) & sum67(sum67'left) & sum67);
       sum82 <= (sum68(sum68'left) & sum68(sum68'left) & sum68) + (sum69(sum69'left) & sum69(sum69'left) & sum69) + (sum70(sum70'left) & sum70(sum70'left) & sum70) + (sum71(sum71'left) & sum71(sum71'left) & sum71);
       sum83 <= (sum72(sum72'left) & sum72(sum72'left) & sum72) + (sum73(sum73'left) & sum73(sum73'left) & sum73) + (sum74(sum74'left) & sum74(sum74'left) & sum74) + (sum75(sum75'left) & sum75(sum75'left) & sum75);


       sum21 <= (sum17(sum17'left) & sum17(sum17'left) & sum17) + (sum18(sum18'left) & sum18(sum18'left) & sum18) + (sum19(sum19'left) & sum19(sum19'left) & sum19) + (sum20(sum20'left) & sum20(sum20'left) & sum20); 
       sum42 <= (sum38(sum38'left) & sum38(sum38'left) & sum38) + (sum39(sum39'left) & sum39(sum39'left) & sum39) + (sum40(sum40'left) & sum40(sum40'left) & sum40) + (sum41(sum41'left) & sum41(sum41'left) & sum41);

       sum84 <= (sum76(sum76'left) & sum76(sum76'left) & sum76) + (sum77(sum77'left) & sum77(sum77'left) & sum77) + (sum78(sum78'left) & sum78(sum78'left) & sum78) + (sum79(sum79'left) & sum79(sum79'left) & sum79); 
       sum85 <= (sum80(sum80'left) & sum80(sum80'left) & sum80) + (sum81(sum81'left) & sum81(sum81'left) & sum81) + (sum82(sum82'left) & sum82(sum82'left) & sum82) + (sum83(sum83'left) & sum83(sum83'left) & sum83);

       sum43 <= (sum21(sum21'left) & sum21(sum21'left) & sum21) + (sum42(sum42'left) & sum42(sum42'left) & sum42) + (sum84(sum84'left) & sum84(sum84'left) & sum84) + (sum85(sum85'left) & sum85(sum85'left) & sum85);
    end if;
  end process p_sums;

d_out <= sum43(sum43'left downto sum43'left -W +1);

end a;