package entropy_encoder_pack is 
type Dout_type  is array ( 0 to 32 ) of std_logic_vector(7-1 downto 0);
end package entropy_encoder_pack;
